--------------------------------------------------------------------------------
-- Company: UNIVERSITY OF MARYLAND
--
-- File: USB_EXEC.vhd
-- File history:  REV A
--     
-- Description: 
--      THIS MODULE LOOKS AT THE USB INTERFACE SIGNALS TO DETERMINE WHEN THE MODULE HAS BEEN ACTIVATED IN THE SYNC 245 MODE.
--      THE SYNC 245 MODE IS EVIDENT ONCE THE 60 MHZ CLOCK IS PRESENT.
--      BASICALLY, A COUNTER RUNNING FROM THE 60 MHZ DOMAIN DIRECT FROM THE USB MODULE IS ENABLED BY THE 40 MHZ DOMAIN TO DETERMINE THE STATUS OF THE 60MHZ DOMAIN CLOCK.
--      THE USB INTERFACE IS ENABLED IN 2 STEPS ONCE AN ACTIVE CLOCK IS DETECTED.  
--      (1) THE CCC_60M USED TO GENERATED AN ON-BOARD SYNCHRONOUS 60 MHZ CLOCK IS ENABLED.
--      (2) ONCE THE CCC_60M LOCK IS ASSERTED, THEN A SYNCHRONOUS RELEASE OF THE RESET SIGNAL DEDICATED ONLY FOR THE USB_INTERFACE.VHD IS PERFORMED.
--
-- Targeted device: <Family::ProASIC3E> <Die::A3PE1500> <Package::208 PQFP>
-- Author: <Name>
--
--------------------------------------------------------------------------------

library IEEE;

use IEEE.std_logic_1164.all;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_MISC.ALL;

library proasic3e;
use proasic3e.all;

entity USB_EXEC is
port (
            RESETB              :   IN      STD_LOGIC;                      -- ACTIVE LOW RESET
            CLK_40MHZ_GEN       :   IN      STD_LOGIC;                      -- CLOCK SYNCHRONOUS TO THE 160MHZ CCC CLOCK FROM THE SERIALIZER

            CLK60MHZ            :   IN      STD_LOGIC;                      -- CLOCK FROM THE USM MODULE DERIVED FROM A 12MHZ CRYSTAL ON-BOARD THE USB MODULE PLL
                                                                            -- THIS CLOCK IS NOT ACTIVE AT POWER ON.  REQUIRES USB HOST ACTION TO ENABLE THE OUTPUT.
            USB_RESET_B         :   OUT     STD_LOGIC                       -- ACTIVE LOW RESET DEDICATED FOR THE USB VHDL STATE MACHINE--SYCHRONOUS RELEASE RELATIVE TO THE 60 MHZ CLOCK

    );

end USB_EXEC;

architecture RTL_LOGIC of USB_EXEC is

--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
-- DEFINE INTERNAL SIGNALS
--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++

-- CLK60MHZ CLOCK DOMAIN SIGNALS
    SIGNAL  N_T_CNT60M, T_CNT60M                :   STD_LOGIC_VECTOR(7 DOWNTO 0);       -- TEST COUNTER USED TO VERIFY USB CLOCK IS RUNNING

    SIGNAL  CNT_EN_60M0S                        :   STD_LOGIC;                          -- ENABLE DERIVED FROM THE 40 MHZ CLOCK DOMAIN, BUT BEING RESYNC'D TO THE 60 MHZ CLOCK DOMAIN
    SIGNAL  CNT_EN_60M1S                        :   STD_LOGIC;                          --  "
    SIGNAL  CNT_EN_60M2S                        :   STD_LOGIC;                          --  "  --> USE THIS RESYNC'D VERSION OF THE FLAG

    SIGNAL  N_TERMCNT_FG60M, TERMCNT_FG60M      :   STD_LOGIC;                          -- TERMINAL COUNT FLAG GENERATED BY THE 60MHZ TEST COUNTER

    SIGNAL  USB_EN_60M_S                        :   STD_LOGIC;                          -- USB ENABLE FROM THE 40 MHZ CLOCK DOMAIN, BUT BEING RESYNC'D TO THE 60 MHZ CLOCK DOMAIN
    SIGNAL  USB_EN_60M_1S                       :   STD_LOGIC;                          --  "
    SIGNAL  USB_EN_60M_2S                       :   STD_LOGIC;                          --  "  --> USE THIS RESYNC'D VERSION OF THE FLAG

-- CLK_40MHZ_GEN DOMAIN SIGNALS
    SIGNAL  N_CNT_EN_40M, CNT_EN_40M            :   STD_LOGIC;                          -- COUNTER ENABLE GENERATED BY THE 40 MHZ CLOCK DOMAIN FOR THE 60 MHZ CLOCK DOMAIN COUNTER

    SIGNAL  TERMCNT_FG40M0S                     :   STD_LOGIC;                          -- TERM-COINT FLAG FROM THE 60 MHZ CLOCK DOMAIN, BUT BEING RESYNC'D TO THE 40 MHZ CLOCK DOMAIN
    SIGNAL  TERMCNT_FG40M1S                     :   STD_LOGIC;                          --  "
    SIGNAL  TERMCNT_FG40M2S                     :   STD_LOGIC;                          --  "  --> USE THIS RESYNC'D VERSION OF THE FLAG

    SIGNAL  N_USB_EN_40M, USB_EN_40M            :   STD_LOGIC;                          -- ACTIVE HIGH ENABLE FOR THE USB_INTERFACE.VHD MODULE GENERATED BY THE 40 MHZ CLOCK DOMAIN

-- DEFINE THE STATES FOR THE 40 MHZ CLOCK DOMAIN STATE MACHINE THAT CONTROLS WHEN THE USB_INTERFACE.VHD IS ENABLED
    TYPE TEST_SM_STATES IS   ( INIT, CHK_1ST_TEST, CLR_FOR_2ND_TEST, CHK_2ND_TEST, SIT_SS );
    SIGNAL N_TEST_SM, TEST_SM                   :   TEST_SM_STATES;

begin

--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
-- DEFINE INTERNAL REGISTERS
--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
-- 60 MHZ CLOCK DOMAIN
    REG60M:PROCESS(CLK60MHZ, RESETB)
        BEGIN
            IF (RESETB = '0')   THEN 
                T_CNT60M        <=  (OTHERS => '0');

                CNT_EN_60M0S    <=  '0';
                CNT_EN_60M1S    <=  '0';
                CNT_EN_60M2S    <=  '0';

                TERMCNT_FG60M   <=  '0';

                USB_EN_60M_S    <=  '0';
                USB_EN_60M_1S   <=  '0';
                USB_EN_60M_2S   <=  '0';

            ELSIF (CLK60MHZ'EVENT AND CLK60MHZ='1')   THEN
                T_CNT60M        <=  N_T_CNT60M;                     -- 60 MHZ TEST COUNTER

                CNT_EN_60M0S    <=  CNT_EN_40M;                     -- CLOCK DOMAIN CROSSING RESYNC ASSIGNMENTS
                CNT_EN_60M1S    <=  CNT_EN_60M0S;                   --  "
                CNT_EN_60M2S    <=  CNT_EN_60M1S;                   --  "  --> USE THIS RESYNC'D VERSION OF THE SIGNAL

                TERMCNT_FG60M   <=  N_TERMCNT_FG60M;

                USB_EN_60M_S    <=  USB_EN_40M;
                USB_EN_60M_1S   <=  USB_EN_60M_S;
                USB_EN_60M_2S   <=  USB_EN_60M_1S;

            END IF;

        END PROCESS REG60M;

-- 40 MHZ CLOCK DOMAIN
    REG40M:PROCESS(CLK_40MHZ_GEN, RESETB)
        BEGIN
            IF (RESETB = '0')   THEN 
                CNT_EN_40M      <=  '0';

                TEST_SM         <=  INIT;

                TERMCNT_FG40M0S <=  '0';
                TERMCNT_FG40M1S <=  '0';
                TERMCNT_FG40M2S <=  '0';

                USB_EN_40M      <=  '0';                            -- ACTIVE HIGH--SO KEEP DISABLED AS DEFAULT
                
            ELSIF (CLK_40MHZ_GEN'EVENT AND CLK_40MHZ_GEN='1')   THEN
                CNT_EN_40M      <=  N_CNT_EN_40M;

                TEST_SM         <=  N_TEST_SM;

                TERMCNT_FG40M0S <=  TERMCNT_FG60M;                  -- CLOCK DOMAIN CROSSING RESYNC ASSIGNMENTS
                TERMCNT_FG40M1S <=  TERMCNT_FG40M0S;                --  "
                TERMCNT_FG40M2S <=  TERMCNT_FG40M1S;                --  "  --> USE THIS RESYNC'D VERSION OF THE SIGNAL

                USB_EN_40M      <=  N_USB_EN_40M;

            END IF;

        END PROCESS REG40M;

--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
-- DEFINE TEST COUNT OPERATION THAT USES THE 60 MHZ CLOCK DOMAIN
--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++

    TEST_60M:PROCESS(T_CNT60M, CNT_EN_60M2S)
        BEGIN

        -- OPERATE THE 60 MHZ COUNTER WHEN ENABLED
            IF CNT_EN_60M2S = '1'    THEN                   -- USE THE ENEABLE SIGNAL RE-SYNC'D TO THIS DOMAIN

                IF T_CNT60M = ("11111111") THEN             -- PERMANANTLY SET THE TERMCNT_FG60M FLAG WHEN a 255 COUNT IS ACHIEVED
                    N_T_CNT60M          <=  T_CNT60M;
                    N_TERMCNT_FG60M     <=  '1';
                ELSE
                    N_T_CNT60M          <=  T_CNT60M + '1';
                    N_TERMCNT_FG60M     <=  '0';
                END IF;

            ELSE                                            -- CLEAR THE COUNT AND TERMCNT_FG60M FLAG WHENEVER THE COUNTER IS DISABLED
                N_T_CNT60M      <=  ("00000000");
                N_TERMCNT_FG60M <=  '0';

            END IF;

        END PROCESS TEST_60M;

--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
-- DEFINE THE STATE MACHINE THAT CONTROLS THE USB_INTERFACE.VHD PROCESS MASTER ENABLE.  THIS PROCESS USES THE 40 MHZ CLOCK DOMAIN.
--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
    USB_EN_SM:PROCESS(TEST_SM, TERMCNT_FG40M2S)
        BEGIN

            CASE TEST_SM IS

                WHEN INIT       =>                              -- INITIAL POR STATE FOR THE STATE MACHINE
                    N_TEST_SM       <=  CHK_1ST_TEST;
                    N_CNT_EN_40M    <=  '0';
                    N_USB_EN_40M    <=  '0';                    -- ACTIVE HIGH--KEEP THE USB_INTERFACE.VHD MODULE DISABLED

                WHEN CHK_1ST_TEST =>                            -- WAIT HERE UNTIL THE ENABLED 60 MHZ TEST COUNTER REACHES A TERMINAL COUNT
                    N_CNT_EN_40M    <=  '1';                    -- ENABLE THE 60 MHZ TEST COUNTER
                    N_USB_EN_40M    <=  '0';                    -- ACTIVE HIGH--KEEP THE USB_INTERFACE.VHD MODULE DISABLED

                    IF TERMCNT_FG40M2S = '1' THEN
                        N_TEST_SM       <=  CLR_FOR_2ND_TEST;   -- REPEAT TEST A SECOND TIME
                        N_CNT_EN_40M    <=  '0';                -- DISABLE THE 60 MHZ TEST COUNTER (OVER-WRITES ABOVE ASSIGNMENT)
                    ELSE
                        N_TEST_SM       <=  CHK_1ST_TEST;
                    END IF;

                WHEN CLR_FOR_2ND_TEST =>                        -- REPEAT THE TEST
                    N_CNT_EN_40M    <=  '0';                    -- DISABLE THE 60 MHZ TEST COUNTER
                    N_USB_EN_40M    <=  '0';                    -- ACTIVE HIGH--KEEP THE USB_INTERFACE.VHD MODULE DISABLED

                    IF TERMCNT_FG40M2S = '0' THEN               -- WAIT FOR THE 60 MHZ COUNTER TO RESET BACK TO 0
                        N_TEST_SM       <=  CHK_2ND_TEST;       -- REPEAT TEST A SECOND TIME
                    ELSE
                        N_TEST_SM       <=  CLR_FOR_2ND_TEST;
                    END IF;

                WHEN CHK_2ND_TEST =>                            -- 2ND TEST--WAIT HERE UNTIL THE ENABLED 60 MHZ TEST COUNTER REACHES A TERMINAL COUNT
                    N_CNT_EN_40M    <=  '1';                    -- RE-ENABLE THE 60 MHZ TEST COUNTER
                    N_USB_EN_40M    <=  '0';                    -- ACTIVE HIGH--KEEP THE USB_INTERFACE.VHD MODULE DISABLED

                    IF TERMCNT_FG40M2S = '1' THEN
                        N_TEST_SM       <=  SIT_SS;
                    ELSE
                        N_TEST_SM       <=  CHK_2ND_TEST;
                    END IF;

                WHEN SIT_SS     =>                              -- 2 TESTS COMPLETE-SIT HERE AT STEADY STATE INDEFINITLY (UNTIL ANOTHER POR)
                    N_TEST_SM       <=  SIT_SS;
                    N_CNT_EN_40M    <=  '0';                    -- DISABLE THE 60 MHZ TEST COUNTER TO SAVE THE POWER
                    N_USB_EN_40M    <=  '1';                    -- ACTIVE HIGH--KEEP THE USB_INTERFACE.VHD MODULE DISABLED

                WHEN OTHERS     =>
                    N_TEST_SM       <=  INIT;
                    N_CNT_EN_40M    <=  '0';                    -- DISABLE THE 60 MHZ TEST COUNTER
                    N_USB_EN_40M    <=  '0';                    -- ACTIVE HIGH--ENABLE THE USB_INTERFACE.VHD MODULE !!!!!!!

            END CASE;

    END PROCESS USB_EN_SM;

--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
-- CONNECT INTERNAL SIGNALS TO EXTERNAL PORTS
USB_RESET_B     <=  USB_EN_60M_2S;

end RTL_LOGIC;
