-- Version: v11.9 SP2 11.9.2.1

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SLAVE_DES320S_1_17 is

    port( ELK_RX_SER_WORD_1      : out   std_logic_vector(7 downto 0);
          BIT_OS_SEL_2_0         : in    std_logic;
          BIT_OS_SEL_1           : in    std_logic_vector(2 downto 0);
          BIT_OS_SEL_0_0         : in    std_logic;
          BIT_OS_SEL_0_d0        : in    std_logic;
          CLK_40M_GL             : in    std_logic;
          CCC_160M_FXD           : in    std_logic;
          ELK_IN_R               : in    std_logic;
          ELK_IN_F               : in    std_logic;
          MASTER_DCB_POR_B_i_0_i : in    std_logic;
          CCC_160M_ADJ           : in    std_logic
        );

end SLAVE_DES320S_1_17;

architecture DEF_ARCH of SLAVE_DES320S_1_17 is 

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal N_17, \ARB_BYTE[0]_net_1\, \ARB_BYTE[4]_net_1\, N_18, 
        \ARB_BYTE[1]_net_1\, \ARB_BYTE[5]_net_1\, N_19, 
        \ARB_BYTE[2]_net_1\, \ARB_BYTE[6]_net_1\, N_20, 
        \ARB_BYTE[3]_net_1\, \ARB_BYTE[7]_net_1\, N_21, 
        \ARB_BYTE[8]_net_1\, N_22, \ARB_BYTE[9]_net_1\, N_23, 
        \ARB_BYTE[10]_net_1\, N_24, \ARB_BYTE[11]_net_1\, N_31, 
        \ARB_BYTE[12]_net_1\, N_32, \ARB_BYTE[13]_net_1\, N_33, 
        N_34, N_35, N_36, N_37, N_38, N_39, N_40, N_56, 
        \ARB_BYTE[14]_net_1\, N_64, \N_RECD_SER_WORD[0]\, 
        \N_RECD_SER_WORD[1]\, \N_RECD_SER_WORD[2]\, 
        \N_RECD_SER_WORD[3]\, \N_RECD_SER_WORD[4]\, 
        \N_RECD_SER_WORD[5]\, \N_RECD_SER_WORD[6]\, 
        \N_RECD_SER_WORD[7]\, \ADJ_SER_IN_F_0DEL\, 
        \ADJ_SER_IN_R_0DEL\, \ADJ_SER_IN_F_1DEL\, 
        \ADJ_SER_IN_R_1DEL\, \Q[0]_net_1\, \ADJ_Q[0]_net_1\, 
        \Q[1]_net_1\, \ADJ_Q[1]_net_1\, \Q[2]_net_1\, 
        \ADJ_Q[2]_net_1\, \Q[3]_net_1\, \ADJ_Q[3]_net_1\, 
        \Q[4]_net_1\, \ADJ_Q[4]_net_1\, \Q[5]_net_1\, 
        \ADJ_Q[5]_net_1\, \Q[6]_net_1\, \ADJ_Q[6]_net_1\, 
        \Q[7]_net_1\, \ADJ_Q[7]_net_1\, \Q[8]_net_1\, 
        \ADJ_Q[8]_net_1\, \Q[9]_net_1\, \ADJ_Q[9]_net_1\, 
        \Q[10]_net_1\, \ADJ_Q[10]_net_1\, \Q[11]_net_1\, 
        \ADJ_Q[11]_net_1\, \Q[12]_net_1\, \ADJ_Q[12]_net_1\, 
        \Q[13]_net_1\, \ADJ_Q[13]_net_1\, \Q[14]_net_1\, 
        \ADJ_Q[14]_net_1\, \ARB_WRD_40M_FIXED[0]_net_1\, 
        \ARB_WRD_40M_FIXED[1]_net_1\, 
        \ARB_WRD_40M_FIXED[2]_net_1\, 
        \ARB_WRD_40M_FIXED[3]_net_1\, 
        \ARB_WRD_40M_FIXED[4]_net_1\, 
        \ARB_WRD_40M_FIXED[5]_net_1\, 
        \ARB_WRD_40M_FIXED[6]_net_1\, 
        \ARB_WRD_40M_FIXED[7]_net_1\, 
        \ARB_WRD_40M_FIXED[8]_net_1\, 
        \ARB_WRD_40M_FIXED[9]_net_1\, 
        \ARB_WRD_40M_FIXED[10]_net_1\, 
        \ARB_WRD_40M_FIXED[11]_net_1\, 
        \ARB_WRD_40M_FIXED[12]_net_1\, 
        \ARB_WRD_40M_FIXED[13]_net_1\, 
        \ARB_WRD_40M_FIXED[14]_net_1\, \GND\, \VCC\ : std_logic;

begin 


    \RECD_SER_WORD_RNO[5]\ : MX2
      port map(A => N_38, B => N_39, S => BIT_OS_SEL_2_0, Y => 
        \N_RECD_SER_WORD[5]\);
    
    \ARB_WRD_40M_FIXED[9]\ : DFN1C0
      port map(D => \Q[9]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[9]_net_1\);
    
    \ADJ_Q[4]\ : DFN1C0
      port map(D => \ADJ_Q[2]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[4]_net_1\);
    
    \ARB_BYTE[6]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[6]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[6]_net_1\);
    
    ADJ_SER_IN_F_1DEL : DFN1C0
      port map(D => \ADJ_SER_IN_F_0DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_F_1DEL\);
    
    \ARB_BYTE[0]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[0]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[0]_net_1\);
    
    \Q[11]\ : DFN1C0
      port map(D => \ADJ_Q[11]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[11]_net_1\);
    
    \ADJ_Q[8]\ : DFN1C0
      port map(D => \ADJ_Q[6]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[8]_net_1\);
    
    \ARB_BYTE_RNI30OT1[13]\ : MX2
      port map(A => N_24, B => N_32, S => BIT_OS_SEL_0_0, Y => 
        N_40);
    
    \ARB_BYTE_RNIDOP9[4]\ : MX2
      port map(A => \ARB_BYTE[4]_net_1\, B => \ARB_BYTE[8]_net_1\, 
        S => BIT_OS_SEL_0_d0, Y => N_21);
    
    \ADJ_Q[6]\ : DFN1C0
      port map(D => \ADJ_Q[4]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[6]_net_1\);
    
    \ADJ_Q[12]\ : DFN1C0
      port map(D => \ADJ_Q[10]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[12]_net_1\);
    
    \RECD_SER_WORD_RNO_1[0]\ : MX2
      port map(A => \ARB_BYTE[0]_net_1\, B => \ARB_BYTE[4]_net_1\, 
        S => BIT_OS_SEL_0_d0, Y => N_17);
    
    \Q[1]\ : DFN1C0
      port map(D => \ADJ_Q[1]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[1]_net_1\);
    
    \ARB_BYTE_RNI7IP9[1]\ : MX2
      port map(A => \ARB_BYTE[1]_net_1\, B => \ARB_BYTE[5]_net_1\, 
        S => BIT_OS_SEL_0_d0, Y => N_18);
    
    \ARB_BYTE[4]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[4]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[4]_net_1\);
    
    \ADJ_Q[2]\ : DFN1C0
      port map(D => \ADJ_Q[0]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[2]_net_1\);
    
    \RECD_SER_WORD_RNO_1[7]\ : MX2
      port map(A => \ARB_BYTE[10]_net_1\, B => 
        \ARB_BYTE[14]_net_1\, S => BIT_OS_SEL_1(2), Y => N_56);
    
    \RECD_SER_WORD[4]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[4]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_1(4));
    
    \Q[5]\ : DFN1C0
      port map(D => \ADJ_Q[5]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[5]_net_1\);
    
    \ADJ_Q[11]\ : DFN1C0
      port map(D => \ADJ_Q[9]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[11]_net_1\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \ADJ_Q[3]\ : DFN1C0
      port map(D => \ADJ_Q[1]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[3]_net_1\);
    
    \Q[10]\ : DFN1C0
      port map(D => \ADJ_Q[10]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[10]_net_1\);
    
    \ARB_WRD_40M_FIXED[6]\ : DFN1C0
      port map(D => \Q[6]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[6]_net_1\);
    
    \ARB_WRD_40M_FIXED[1]\ : DFN1C0
      port map(D => \Q[1]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[1]_net_1\);
    
    \RECD_SER_WORD[3]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[3]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_1(3));
    
    \RECD_SER_WORD[0]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[0]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_1(0));
    
    \RECD_SER_WORD_RNO[3]\ : MX2
      port map(A => N_36, B => N_37, S => BIT_OS_SEL_2_0, Y => 
        \N_RECD_SER_WORD[3]\);
    
    \Q[0]\ : DFN1C0
      port map(D => \ADJ_Q[0]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[0]_net_1\);
    
    \ARB_BYTE_RNITAP11[1]\ : MX2
      port map(A => N_18, B => N_20, S => BIT_OS_SEL_0_0, Y => 
        N_34);
    
    \RECD_SER_WORD_RNO_0[7]\ : MX2
      port map(A => N_31, B => N_56, S => BIT_OS_SEL_1(1), Y => 
        N_64);
    
    \Q[7]\ : DFN1C0
      port map(D => \ADJ_Q[7]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[7]_net_1\);
    
    \ARB_BYTE[14]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[14]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[14]_net_1\);
    
    \ARB_WRD_40M_FIXED[2]\ : DFN1C0
      port map(D => \Q[2]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[2]_net_1\);
    
    \ARB_WRD_40M_FIXED[14]\ : DFN1C0
      port map(D => \Q[14]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[14]_net_1\);
    
    \RECD_SER_WORD_RNO[2]\ : MX2
      port map(A => N_35, B => N_36, S => BIT_OS_SEL_1(0), Y => 
        \N_RECD_SER_WORD[2]\);
    
    \ARB_BYTE_RNIOQON[6]\ : MX2
      port map(A => \ARB_BYTE[6]_net_1\, B => 
        \ARB_BYTE[10]_net_1\, S => BIT_OS_SEL_0_d0, Y => N_23);
    
    \ARB_BYTE[2]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[2]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[2]_net_1\);
    
    \ADJ_Q[7]\ : DFN1C0
      port map(D => \ADJ_Q[5]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[7]_net_1\);
    
    \ARB_BYTE[8]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[8]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[8]_net_1\);
    
    \RECD_SER_WORD[5]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[5]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_1(5));
    
    \ARB_BYTE_RNISUON[12]\ : MX2
      port map(A => \ARB_BYTE[8]_net_1\, B => 
        \ARB_BYTE[12]_net_1\, S => BIT_OS_SEL_0_d0, Y => N_31);
    
    \ARB_BYTE[12]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[12]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[12]_net_1\);
    
    \RECD_SER_WORD[1]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[1]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_1(1));
    
    \ARB_BYTE_RNIBMP9[3]\ : MX2
      port map(A => \ARB_BYTE[3]_net_1\, B => \ARB_BYTE[7]_net_1\, 
        S => BIT_OS_SEL_0_d0, Y => N_20);
    
    \Q[3]\ : DFN1C0
      port map(D => \ADJ_Q[3]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[3]_net_1\);
    
    ADJ_SER_IN_F_0DEL : DFN1C0
      port map(D => ELK_IN_F, CLK => CCC_160M_ADJ, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_F_0DEL\);
    
    \RECD_SER_WORD_RNO[7]\ : MX2
      port map(A => N_40, B => N_64, S => BIT_OS_SEL_2_0, Y => 
        \N_RECD_SER_WORD[7]\);
    
    \RECD_SER_WORD_RNO[1]\ : MX2
      port map(A => N_34, B => N_35, S => BIT_OS_SEL_1(0), Y => 
        \N_RECD_SER_WORD[1]\);
    
    \ARB_WRD_40M_FIXED[4]\ : DFN1C0
      port map(D => \Q[4]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[4]_net_1\);
    
    \RECD_SER_WORD_RNO[0]\ : MX2
      port map(A => N_33, B => N_34, S => BIT_OS_SEL_1(0), Y => 
        \N_RECD_SER_WORD[0]\);
    
    \Q[6]\ : DFN1C0
      port map(D => \ADJ_Q[6]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[6]_net_1\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \ARB_WRD_40M_FIXED[8]\ : DFN1C0
      port map(D => \Q[8]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[8]_net_1\);
    
    \ARB_BYTE[11]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[11]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[11]_net_1\);
    
    \Q[9]\ : DFN1C0
      port map(D => \ADJ_Q[9]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[9]_net_1\);
    
    \Q[14]\ : DFN1C0
      port map(D => \ADJ_Q[14]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[14]_net_1\);
    
    ADJ_SER_IN_R_0DEL : DFN1C0
      port map(D => ELK_IN_R, CLK => CCC_160M_ADJ, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_R_0DEL\);
    
    \Q[13]\ : DFN1C0
      port map(D => \ADJ_Q[13]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[13]_net_1\);
    
    \ARB_BYTE_RNI1FP11[2]\ : MX2
      port map(A => N_19, B => N_21, S => BIT_OS_SEL_0_0, Y => 
        N_35);
    
    \ARB_BYTE[9]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[9]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[9]_net_1\);
    
    ADJ_SER_IN_R_1DEL : DFN1C0
      port map(D => \ADJ_SER_IN_R_0DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_R_1DEL\);
    
    \ARB_BYTE[10]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[10]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[10]_net_1\);
    
    \ADJ_Q[9]\ : DFN1C0
      port map(D => \ADJ_Q[7]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[9]_net_1\);
    
    \RECD_SER_WORD[7]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[7]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_1(7));
    
    \ARB_WRD_40M_FIXED[5]\ : DFN1C0
      port map(D => \Q[5]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[5]_net_1\);
    
    \ARB_WRD_40M_FIXED[12]\ : DFN1C0
      port map(D => \Q[12]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[12]_net_1\);
    
    \ARB_WRD_40M_FIXED[11]\ : DFN1C0
      port map(D => \Q[11]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[11]_net_1\);
    
    \ARB_WRD_40M_FIXED[0]\ : DFN1C0
      port map(D => \Q[0]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[0]_net_1\);
    
    \ADJ_Q[10]\ : DFN1C0
      port map(D => \ADJ_Q[8]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[10]_net_1\);
    
    \Q[2]\ : DFN1C0
      port map(D => \ADJ_Q[2]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[2]_net_1\);
    
    \ARB_BYTE_RNIGLOF1[4]\ : MX2
      port map(A => N_21, B => N_23, S => BIT_OS_SEL_0_0, Y => 
        N_37);
    
    \ADJ_Q[1]\ : DFN1C0
      port map(D => \ADJ_SER_IN_F_1DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[1]_net_1\);
    
    \RECD_SER_WORD[6]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[6]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_1(6));
    
    \RECD_SER_WORD[2]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[2]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_1(2));
    
    \ARB_BYTE_RNIVRNT1[6]\ : MX2
      port map(A => N_23, B => N_31, S => BIT_OS_SEL_0_0, Y => 
        N_39);
    
    \ARB_BYTE_RNIU0PN[13]\ : MX2
      port map(A => \ARB_BYTE[9]_net_1\, B => 
        \ARB_BYTE[13]_net_1\, S => BIT_OS_SEL_0_d0, Y => N_32);
    
    \ADJ_Q[13]\ : DFN1C0
      port map(D => \ADJ_Q[11]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[13]_net_1\);
    
    \Q[8]\ : DFN1C0
      port map(D => \ADJ_Q[8]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[8]_net_1\);
    
    \ARB_BYTE[5]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[5]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[5]_net_1\);
    
    \ADJ_Q[14]\ : DFN1C0
      port map(D => \ADJ_Q[12]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[14]_net_1\);
    
    \RECD_SER_WORD_RNO[4]\ : MX2
      port map(A => N_37, B => N_38, S => BIT_OS_SEL_2_0, Y => 
        \N_RECD_SER_WORD[4]\);
    
    \Q[12]\ : DFN1C0
      port map(D => \ADJ_Q[12]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[12]_net_1\);
    
    \ARB_BYTE[13]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[13]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[13]_net_1\);
    
    \ARB_WRD_40M_FIXED[3]\ : DFN1C0
      port map(D => \Q[3]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[3]_net_1\);
    
    \ARB_BYTE[7]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[7]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[7]_net_1\);
    
    \RECD_SER_WORD_RNO_0[0]\ : MX2
      port map(A => N_17, B => N_19, S => BIT_OS_SEL_0_0, Y => 
        N_33);
    
    \Q[4]\ : DFN1C0
      port map(D => \ADJ_Q[4]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[4]_net_1\);
    
    \ARB_WRD_40M_FIXED[7]\ : DFN1C0
      port map(D => \Q[7]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[7]_net_1\);
    
    \RECD_SER_WORD_RNO[6]\ : MX2
      port map(A => N_39, B => N_40, S => BIT_OS_SEL_2_0, Y => 
        \N_RECD_SER_WORD[6]\);
    
    \ARB_BYTE[3]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[3]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[3]_net_1\);
    
    \ADJ_Q[5]\ : DFN1C0
      port map(D => \ADJ_Q[3]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[5]_net_1\);
    
    \ARB_BYTE_RNI5JP11[3]\ : MX2
      port map(A => N_20, B => N_22, S => BIT_OS_SEL_0_0, Y => 
        N_36);
    
    \ARB_BYTE[1]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[1]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[1]_net_1\);
    
    \ARB_BYTE_RNI9KP9[2]\ : MX2
      port map(A => \ARB_BYTE[2]_net_1\, B => \ARB_BYTE[6]_net_1\, 
        S => BIT_OS_SEL_0_d0, Y => N_19);
    
    \ARB_WRD_40M_FIXED[13]\ : DFN1C0
      port map(D => \Q[13]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[13]_net_1\);
    
    \ARB_BYTE_RNIFQP9[5]\ : MX2
      port map(A => \ARB_BYTE[5]_net_1\, B => \ARB_BYTE[9]_net_1\, 
        S => BIT_OS_SEL_0_d0, Y => N_22);
    
    \ADJ_Q[0]\ : DFN1C0
      port map(D => \ADJ_SER_IN_R_1DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[0]_net_1\);
    
    \ARB_BYTE_RNIKPOF1[5]\ : MX2
      port map(A => N_22, B => N_24, S => BIT_OS_SEL_0_0, Y => 
        N_38);
    
    \ARB_WRD_40M_FIXED[10]\ : DFN1C0
      port map(D => \Q[10]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[10]_net_1\);
    
    \ARB_BYTE_RNIQSON[11]\ : MX2
      port map(A => \ARB_BYTE[7]_net_1\, B => 
        \ARB_BYTE[11]_net_1\, S => BIT_OS_SEL_0_d0, Y => N_24);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SER320M_3_34_1 is

    port( ELK_TX_DAT                 : in    std_logic_vector(7 downto 0);
          MASTER_SALT_POR_B_i_0_i_4  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_16 : in    std_logic;
          ELK_OUT_R_i_0              : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_1  : in    std_logic;
          ELK_OUT_F_i_0              : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_7  : in    std_logic;
          CLK_40M_GL                 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_14 : in    std_logic;
          CCC_160M_FXD               : in    std_logic
        );

end SER320M_3_34_1;

architecture DEF_ARCH of SER320M_3_34_1 is 

  component DFI1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          QN  : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component DFN1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

    signal SER_OUT_RI_i, \SER_CMD_WORD_R[3]_net_1\, SER_OUT_FI_i, 
        \SER_CMD_WORD_F[3]_net_1\, \N_SER_CMD_WORD_R[0]\, 
        \START_RISE\, \N_SER_CMD_WORD_F[0]\, 
        \N_SER_CMD_WORD_R[3]\, \SER_CMD_WORD_R[2]_net_1\, 
        \N_SER_CMD_WORD_R[2]\, \SER_CMD_WORD_R[1]_net_1\, 
        \N_SER_CMD_WORD_R[1]\, \SER_CMD_WORD_R[0]_net_1\, 
        \N_SER_CMD_WORD_F[3]\, \SER_CMD_WORD_F[2]_net_1\, 
        \N_SER_CMD_WORD_F[2]\, \SER_CMD_WORD_F[1]_net_1\, 
        \N_SER_CMD_WORD_F[1]\, \SER_CMD_WORD_F[0]_net_1\, 
        N_START_RISE, \CLK40M_GEN_DEL0\, \GND\, \VCC\
         : std_logic;

begin 


    SER_OUT_FI : DFI1C0
      port map(D => \SER_CMD_WORD_F[3]_net_1\, CLK => 
        CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_14, QN => 
        SER_OUT_FI_i);
    
    \SER_CMD_WORD_F[3]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[3]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_7, Q => 
        \SER_CMD_WORD_F[3]_net_1\);
    
    \SER_CMD_WORD_R[1]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[1]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_4, Q => 
        \SER_CMD_WORD_R[1]_net_1\);
    
    \SER_CMD_WORD_R[2]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[2]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_4, Q => 
        \SER_CMD_WORD_R[2]_net_1\);
    
    \SER_CMD_WORD_R_RNO[3]\ : MX2
      port map(A => \SER_CMD_WORD_R[2]_net_1\, B => ELK_TX_DAT(7), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_R[3]\);
    
    \SER_CMD_WORD_R_RNO[0]\ : NOR2B
      port map(A => \START_RISE\, B => ELK_TX_DAT(1), Y => 
        \N_SER_CMD_WORD_R[0]\);
    
    \SER_CMD_WORD_F[0]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[0]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_7, Q => 
        \SER_CMD_WORD_F[0]_net_1\);
    
    \SER_CMD_WORD_R_RNO[1]\ : MX2
      port map(A => \SER_CMD_WORD_R[0]_net_1\, B => ELK_TX_DAT(3), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_R[1]\);
    
    \SER_CMD_WORD_F_RNO[2]\ : MX2
      port map(A => \SER_CMD_WORD_F[1]_net_1\, B => ELK_TX_DAT(4), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_F[2]\);
    
    \SER_CMD_WORD_F_RNO[3]\ : MX2
      port map(A => \SER_CMD_WORD_F[2]_net_1\, B => ELK_TX_DAT(6), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_F[3]\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    CLK40M_GEN_DEL0 : DFN1C0
      port map(D => CLK_40M_GL, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_7, Q => \CLK40M_GEN_DEL0\);
    
    SER_OUT_RI : DFI1C0
      port map(D => \SER_CMD_WORD_R[3]_net_1\, CLK => 
        CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_14, QN => 
        SER_OUT_RI_i);
    
    \SER_CMD_WORD_F[2]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[2]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_7, Q => 
        \SER_CMD_WORD_F[2]_net_1\);
    
    \SER_CMD_WORD_F_RNO[1]\ : MX2
      port map(A => \SER_CMD_WORD_F[0]_net_1\, B => ELK_TX_DAT(2), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_F[1]\);
    
    \SER_CMD_WORD_R[0]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[0]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_4, Q => 
        \SER_CMD_WORD_R[0]_net_1\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    START_RISE : DFN1C0
      port map(D => N_START_RISE, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_4, Q => \START_RISE\);
    
    \SER_CMD_WORD_R[3]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[3]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_4, Q => 
        \SER_CMD_WORD_R[3]_net_1\);
    
    \SER_CMD_WORD_F_RNO[0]\ : NOR2B
      port map(A => \START_RISE\, B => ELK_TX_DAT(0), Y => 
        \N_SER_CMD_WORD_F[0]\);
    
    SER_OUT_RDEL : DFN1P0
      port map(D => SER_OUT_RI_i, CLK => CCC_160M_FXD, PRE => 
        MASTER_SALT_POR_B_i_0_i_16, Q => ELK_OUT_R_i_0);
    
    \SER_CMD_WORD_F[1]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[1]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_7, Q => 
        \SER_CMD_WORD_F[1]_net_1\);
    
    START_RISE_RNO : NOR2B
      port map(A => \CLK40M_GEN_DEL0\, B => CLK_40M_GL, Y => 
        N_START_RISE);
    
    \SER_CMD_WORD_R_RNO[2]\ : MX2
      port map(A => \SER_CMD_WORD_R[1]_net_1\, B => ELK_TX_DAT(5), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_R[2]\);
    
    SER_OUT_FDEL : DFN1P0
      port map(D => SER_OUT_FI_i, CLK => CCC_160M_FXD, PRE => 
        MASTER_SALT_POR_B_i_0_i_1, Q => ELK_OUT_F_i_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity DDR_BIDIR_LVDS_DUAL_CLK_1 is

    port( DCB_SALT_SEL_c_i : in    std_logic;
          ELK1_DAT_P       : inout std_logic := 'Z';
          ELK1_DAT_N       : inout std_logic := 'Z';
          ELK_OUT_R_i_0    : in    std_logic;
          ELK_OUT_F_i_0    : in    std_logic;
          CCC_160M_FXD     : in    std_logic;
          CCC_160M_ADJ     : in    std_logic;
          ELK_IN_DDR_F_i   : out   std_logic;
          ELK_IN_DDR_R_i   : out   std_logic
        );

end DDR_BIDIR_LVDS_DUAL_CLK_1;

architecture DEF_ARCH of DDR_BIDIR_LVDS_DUAL_CLK_1 is 

  component DDR_REG
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          QR  : out   std_logic;
          QF  : out   std_logic
        );
  end component;

  component DDR_OUT
    port( DR  : in    std_logic := 'U';
          DF  : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component BIBUF_LVDS
    port( PADP : inout   std_logic;
          PADN : inout   std_logic;
          D    : in    std_logic := 'U';
          E    : in    std_logic := 'U';
          Y    : out   std_logic
        );
  end component;

  component INV
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal ELK_IN_DDR_R, ELK_IN_DDR_F, 
        DDR_BIDIR_LVDS_DUAL_CLK_1_GND, BIBUF_LVDS_0_Y, 
        DDR_OUT_0_Q, \VCC\ : std_logic;

begin 


    DDR_REG_0 : DDR_REG
      port map(D => BIBUF_LVDS_0_Y, CLK => CCC_160M_ADJ, CLR => 
        DDR_BIDIR_LVDS_DUAL_CLK_1_GND, QR => ELK_IN_DDR_R, QF => 
        ELK_IN_DDR_F);
    
    DDR_OUT_0 : DDR_OUT
      port map(DR => ELK_OUT_R_i_0, DF => ELK_OUT_F_i_0, CLK => 
        CCC_160M_FXD, CLR => DDR_BIDIR_LVDS_DUAL_CLK_1_GND, Q => 
        DDR_OUT_0_Q);
    
    BIBUF_LVDS_0 : BIBUF_LVDS
      port map(PADP => ELK1_DAT_P, PADN => ELK1_DAT_N, D => 
        DDR_OUT_0_Q, E => DCB_SALT_SEL_c_i, Y => BIBUF_LVDS_0_Y);
    
    DDR_REG_0_RNI7PO8_0 : INV
      port map(A => ELK_IN_DDR_R, Y => ELK_IN_DDR_R_i);
    
    DDR_REG_0_RNI7PO8 : INV
      port map(A => ELK_IN_DDR_F, Y => ELK_IN_DDR_F_i);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    GND_i : GND
      port map(Y => DDR_BIDIR_LVDS_DUAL_CLK_1_GND);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SYNC_DAT_SEL_1 is

    port( ELK_TX_DAT                 : out   std_logic_vector(7 downto 0);
          PATT_ELK_DAT_1             : in    std_logic_vector(7 downto 0);
          OP_MODE_c_5_0              : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_11 : in    std_logic;
          CLK_40M_GL                 : in    std_logic
        );

end SYNC_DAT_SEL_1;

architecture DEF_ARCH of SYNC_DAT_SEL_1 is 

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \N_SERDAT[0]\, \N_SERDAT[1]\, \N_SERDAT[2]\, 
        \N_SERDAT[3]\, \N_SERDAT[4]\, \N_SERDAT[5]\, 
        \N_SERDAT[6]\, \N_SERDAT[7]\, \GND\, \VCC\ : std_logic;

begin 


    \SERDAT_RNO[4]\ : NOR2A
      port map(A => PATT_ELK_DAT_1(4), B => OP_MODE_c_5_0, Y => 
        \N_SERDAT[4]\);
    
    \SERDAT_RNO[0]\ : NOR2A
      port map(A => PATT_ELK_DAT_1(0), B => OP_MODE_c_5_0, Y => 
        \N_SERDAT[0]\);
    
    \SERDAT[6]\ : DFN1C0
      port map(D => \N_SERDAT[6]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_11, Q => ELK_TX_DAT(6));
    
    \SERDAT[4]\ : DFN1C0
      port map(D => \N_SERDAT[4]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_11, Q => ELK_TX_DAT(4));
    
    \SERDAT_RNO[7]\ : OR2
      port map(A => PATT_ELK_DAT_1(7), B => OP_MODE_c_5_0, Y => 
        \N_SERDAT[7]\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \SERDAT_RNO[3]\ : OR2
      port map(A => PATT_ELK_DAT_1(3), B => OP_MODE_c_5_0, Y => 
        \N_SERDAT[3]\);
    
    \SERDAT_RNO[2]\ : OR2
      port map(A => PATT_ELK_DAT_1(2), B => OP_MODE_c_5_0, Y => 
        \N_SERDAT[2]\);
    
    \SERDAT[5]\ : DFN1C0
      port map(D => \N_SERDAT[5]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_11, Q => ELK_TX_DAT(5));
    
    \SERDAT[7]\ : DFN1C0
      port map(D => \N_SERDAT[7]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_11, Q => ELK_TX_DAT(7));
    
    GND_i : GND
      port map(Y => \GND\);
    
    \SERDAT_RNO[5]\ : NOR2A
      port map(A => PATT_ELK_DAT_1(5), B => OP_MODE_c_5_0, Y => 
        \N_SERDAT[5]\);
    
    \SERDAT[0]\ : DFN1C0
      port map(D => \N_SERDAT[0]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_11, Q => ELK_TX_DAT(0));
    
    \SERDAT_RNO[6]\ : NOR2A
      port map(A => PATT_ELK_DAT_1(6), B => OP_MODE_c_5_0, Y => 
        \N_SERDAT[6]\);
    
    \SERDAT[1]\ : DFN1C0
      port map(D => \N_SERDAT[1]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_11, Q => ELK_TX_DAT(1));
    
    \SERDAT_RNO[1]\ : OR2
      port map(A => PATT_ELK_DAT_1(1), B => OP_MODE_c_5_0, Y => 
        \N_SERDAT[1]\);
    
    \SERDAT[3]\ : DFN1C0
      port map(D => \N_SERDAT[3]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_11, Q => ELK_TX_DAT(3));
    
    \SERDAT[2]\ : DFN1C0
      port map(D => \N_SERDAT[2]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_11, Q => ELK_TX_DAT(2));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity ELINK_SLAVE_INV_2 is

    port( BIT_OS_SEL_0_d0            : in    std_logic;
          BIT_OS_SEL_0_0             : in    std_logic;
          BIT_OS_SEL_1               : in    std_logic_vector(2 downto 0);
          BIT_OS_SEL_2_0             : in    std_logic;
          ELK_RX_SER_WORD_1          : out   std_logic_vector(7 downto 0);
          OP_MODE_c_5_0              : in    std_logic;
          PATT_ELK_DAT_1             : in    std_logic_vector(7 downto 0);
          MASTER_DCB_POR_B_i_0_i     : in    std_logic;
          ELK1_DAT_N                 : inout std_logic := 'Z';
          ELK1_DAT_P                 : inout std_logic := 'Z';
          DCB_SALT_SEL_c_i           : in    std_logic;
          CCC_160M_FXD               : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_14 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_7  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_1  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_16 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_4  : in    std_logic;
          CLK_40M_GL                 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_11 : in    std_logic;
          DEV_RST_B_c_0              : in    std_logic;
          CCC_160M_ADJ               : in    std_logic
        );

end ELINK_SLAVE_INV_2;

architecture DEF_ARCH of ELINK_SLAVE_INV_2 is 

  component SLAVE_DES320S_1_17
    port( ELK_RX_SER_WORD_1      : out   std_logic_vector(7 downto 0);
          BIT_OS_SEL_2_0         : in    std_logic := 'U';
          BIT_OS_SEL_1           : in    std_logic_vector(2 downto 0) := (others => 'U');
          BIT_OS_SEL_0_0         : in    std_logic := 'U';
          BIT_OS_SEL_0_d0        : in    std_logic := 'U';
          CLK_40M_GL             : in    std_logic := 'U';
          CCC_160M_FXD           : in    std_logic := 'U';
          ELK_IN_R               : in    std_logic := 'U';
          ELK_IN_F               : in    std_logic := 'U';
          MASTER_DCB_POR_B_i_0_i : in    std_logic := 'U';
          CCC_160M_ADJ           : in    std_logic := 'U'
        );
  end component;

  component SER320M_3_34_1
    port( ELK_TX_DAT                 : in    std_logic_vector(7 downto 0) := (others => 'U');
          MASTER_SALT_POR_B_i_0_i_4  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_16 : in    std_logic := 'U';
          ELK_OUT_R_i_0              : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_1  : in    std_logic := 'U';
          ELK_OUT_F_i_0              : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_7  : in    std_logic := 'U';
          CLK_40M_GL                 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_14 : in    std_logic := 'U';
          CCC_160M_FXD               : in    std_logic := 'U'
        );
  end component;

  component DDR_BIDIR_LVDS_DUAL_CLK_1
    port( DCB_SALT_SEL_c_i : in    std_logic := 'U';
          ELK1_DAT_P       : inout   std_logic;
          ELK1_DAT_N       : inout   std_logic;
          ELK_OUT_R_i_0    : in    std_logic := 'U';
          ELK_OUT_F_i_0    : in    std_logic := 'U';
          CCC_160M_FXD     : in    std_logic := 'U';
          CCC_160M_ADJ     : in    std_logic := 'U';
          ELK_IN_DDR_F_i   : out   std_logic;
          ELK_IN_DDR_R_i   : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component SYNC_DAT_SEL_1
    port( ELK_TX_DAT                 : out   std_logic_vector(7 downto 0);
          PATT_ELK_DAT_1             : in    std_logic_vector(7 downto 0) := (others => 'U');
          OP_MODE_c_5_0              : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_11 : in    std_logic := 'U';
          CLK_40M_GL                 : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \ELK_IN_F\, ELK_IN_DDR_F_i, \ELK_IN_R\, 
        ELK_IN_DDR_R_i, \ELK_TX_DAT[0]\, \ELK_TX_DAT[1]\, 
        \ELK_TX_DAT[2]\, \ELK_TX_DAT[3]\, \ELK_TX_DAT[4]\, 
        \ELK_TX_DAT[5]\, \ELK_TX_DAT[6]\, \ELK_TX_DAT[7]\, 
        ELK_OUT_R_i_0, ELK_OUT_F_i_0, \GND\, \VCC\ : std_logic;

    for all : SLAVE_DES320S_1_17
	Use entity work.SLAVE_DES320S_1_17(DEF_ARCH);
    for all : SER320M_3_34_1
	Use entity work.SER320M_3_34_1(DEF_ARCH);
    for all : DDR_BIDIR_LVDS_DUAL_CLK_1
	Use entity work.DDR_BIDIR_LVDS_DUAL_CLK_1(DEF_ARCH);
    for all : SYNC_DAT_SEL_1
	Use entity work.SYNC_DAT_SEL_1(DEF_ARCH);
begin 


    U_SLAVE_1ELK : SLAVE_DES320S_1_17
      port map(ELK_RX_SER_WORD_1(7) => ELK_RX_SER_WORD_1(7), 
        ELK_RX_SER_WORD_1(6) => ELK_RX_SER_WORD_1(6), 
        ELK_RX_SER_WORD_1(5) => ELK_RX_SER_WORD_1(5), 
        ELK_RX_SER_WORD_1(4) => ELK_RX_SER_WORD_1(4), 
        ELK_RX_SER_WORD_1(3) => ELK_RX_SER_WORD_1(3), 
        ELK_RX_SER_WORD_1(2) => ELK_RX_SER_WORD_1(2), 
        ELK_RX_SER_WORD_1(1) => ELK_RX_SER_WORD_1(1), 
        ELK_RX_SER_WORD_1(0) => ELK_RX_SER_WORD_1(0), 
        BIT_OS_SEL_2_0 => BIT_OS_SEL_2_0, BIT_OS_SEL_1(2) => 
        BIT_OS_SEL_1(2), BIT_OS_SEL_1(1) => BIT_OS_SEL_1(1), 
        BIT_OS_SEL_1(0) => BIT_OS_SEL_1(0), BIT_OS_SEL_0_0 => 
        BIT_OS_SEL_0_0, BIT_OS_SEL_0_d0 => BIT_OS_SEL_0_d0, 
        CLK_40M_GL => CLK_40M_GL, CCC_160M_FXD => CCC_160M_FXD, 
        ELK_IN_R => \ELK_IN_R\, ELK_IN_F => \ELK_IN_F\, 
        MASTER_DCB_POR_B_i_0_i => MASTER_DCB_POR_B_i_0_i, 
        CCC_160M_ADJ => CCC_160M_ADJ);
    
    U_ELK1_CMD_TX : SER320M_3_34_1
      port map(ELK_TX_DAT(7) => \ELK_TX_DAT[7]\, ELK_TX_DAT(6)
         => \ELK_TX_DAT[6]\, ELK_TX_DAT(5) => \ELK_TX_DAT[5]\, 
        ELK_TX_DAT(4) => \ELK_TX_DAT[4]\, ELK_TX_DAT(3) => 
        \ELK_TX_DAT[3]\, ELK_TX_DAT(2) => \ELK_TX_DAT[2]\, 
        ELK_TX_DAT(1) => \ELK_TX_DAT[1]\, ELK_TX_DAT(0) => 
        \ELK_TX_DAT[0]\, MASTER_SALT_POR_B_i_0_i_4 => 
        MASTER_SALT_POR_B_i_0_i_4, MASTER_SALT_POR_B_i_0_i_16 => 
        MASTER_SALT_POR_B_i_0_i_16, ELK_OUT_R_i_0 => 
        ELK_OUT_R_i_0, MASTER_SALT_POR_B_i_0_i_1 => 
        MASTER_SALT_POR_B_i_0_i_1, ELK_OUT_F_i_0 => ELK_OUT_F_i_0, 
        MASTER_SALT_POR_B_i_0_i_7 => MASTER_SALT_POR_B_i_0_i_7, 
        CLK_40M_GL => CLK_40M_GL, MASTER_SALT_POR_B_i_0_i_14 => 
        MASTER_SALT_POR_B_i_0_i_14, CCC_160M_FXD => CCC_160M_FXD);
    
    U_DDR_ELK1 : DDR_BIDIR_LVDS_DUAL_CLK_1
      port map(DCB_SALT_SEL_c_i => DCB_SALT_SEL_c_i, ELK1_DAT_P
         => ELK1_DAT_P, ELK1_DAT_N => ELK1_DAT_N, ELK_OUT_R_i_0
         => ELK_OUT_R_i_0, ELK_OUT_F_i_0 => ELK_OUT_F_i_0, 
        CCC_160M_FXD => CCC_160M_FXD, CCC_160M_ADJ => 
        CCC_160M_ADJ, ELK_IN_DDR_F_i => ELK_IN_DDR_F_i, 
        ELK_IN_DDR_R_i => ELK_IN_DDR_R_i);
    
    ELK_IN_F : DFN1C0
      port map(D => ELK_IN_DDR_F_i, CLK => CCC_160M_ADJ, CLR => 
        DEV_RST_B_c_0, Q => \ELK_IN_F\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    U_ELK1_SERDAT_SOURCE : SYNC_DAT_SEL_1
      port map(ELK_TX_DAT(7) => \ELK_TX_DAT[7]\, ELK_TX_DAT(6)
         => \ELK_TX_DAT[6]\, ELK_TX_DAT(5) => \ELK_TX_DAT[5]\, 
        ELK_TX_DAT(4) => \ELK_TX_DAT[4]\, ELK_TX_DAT(3) => 
        \ELK_TX_DAT[3]\, ELK_TX_DAT(2) => \ELK_TX_DAT[2]\, 
        ELK_TX_DAT(1) => \ELK_TX_DAT[1]\, ELK_TX_DAT(0) => 
        \ELK_TX_DAT[0]\, PATT_ELK_DAT_1(7) => PATT_ELK_DAT_1(7), 
        PATT_ELK_DAT_1(6) => PATT_ELK_DAT_1(6), PATT_ELK_DAT_1(5)
         => PATT_ELK_DAT_1(5), PATT_ELK_DAT_1(4) => 
        PATT_ELK_DAT_1(4), PATT_ELK_DAT_1(3) => PATT_ELK_DAT_1(3), 
        PATT_ELK_DAT_1(2) => PATT_ELK_DAT_1(2), PATT_ELK_DAT_1(1)
         => PATT_ELK_DAT_1(1), PATT_ELK_DAT_1(0) => 
        PATT_ELK_DAT_1(0), OP_MODE_c_5_0 => OP_MODE_c_5_0, 
        MASTER_SALT_POR_B_i_0_i_11 => MASTER_SALT_POR_B_i_0_i_11, 
        CLK_40M_GL => CLK_40M_GL);
    
    ELK_IN_R : DFN1C0
      port map(D => ELK_IN_DDR_R_i, CLK => CCC_160M_ADJ, CLR => 
        DEV_RST_B_c_0, Q => \ELK_IN_R\);
    
    GND_i : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SLAVE_DES320S_1_17_1 is

    port( ELK_RX_SER_WORD_3      : out   std_logic_vector(7 downto 0);
          BIT_OS_SEL_1_0         : in    std_logic;
          BIT_OS_SEL_0           : in    std_logic_vector(2 downto 1);
          BIT_OS_SEL_0_d0        : in    std_logic;
          BIT_OS_SEL_6_0         : in    std_logic;
          BIT_OS_SEL_7_0         : in    std_logic;
          CLK_40M_GL             : in    std_logic;
          CCC_160M_FXD           : in    std_logic;
          ELK_IN_R               : in    std_logic;
          ELK_IN_F               : in    std_logic;
          MASTER_DCB_POR_B_i_0_i : in    std_logic;
          CCC_160M_ADJ           : in    std_logic
        );

end SLAVE_DES320S_1_17_1;

architecture DEF_ARCH of SLAVE_DES320S_1_17_1 is 

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal N_17, \ARB_BYTE[0]_net_1\, \ARB_BYTE[4]_net_1\, N_18, 
        \ARB_BYTE[1]_net_1\, \ARB_BYTE[5]_net_1\, N_19, 
        \ARB_BYTE[2]_net_1\, \ARB_BYTE[6]_net_1\, N_20, 
        \ARB_BYTE[3]_net_1\, \ARB_BYTE[7]_net_1\, N_21, 
        \ARB_BYTE[8]_net_1\, N_22, \ARB_BYTE[9]_net_1\, N_23, 
        \ARB_BYTE[10]_net_1\, N_24, \ARB_BYTE[11]_net_1\, N_31, 
        \ARB_BYTE[12]_net_1\, N_32, \ARB_BYTE[13]_net_1\, N_33, 
        N_34, N_35, N_36, N_37, N_38, N_39, N_40, N_56, 
        \ARB_BYTE[14]_net_1\, N_64, \N_RECD_SER_WORD[0]\, 
        \N_RECD_SER_WORD[1]\, \N_RECD_SER_WORD[2]\, 
        \N_RECD_SER_WORD[3]\, \N_RECD_SER_WORD[4]\, 
        \N_RECD_SER_WORD[5]\, \N_RECD_SER_WORD[6]\, 
        \N_RECD_SER_WORD[7]\, \ADJ_SER_IN_F_0DEL\, 
        \ADJ_SER_IN_R_0DEL\, \ADJ_SER_IN_F_1DEL\, 
        \ADJ_SER_IN_R_1DEL\, \Q[0]_net_1\, \ADJ_Q[0]_net_1\, 
        \Q[1]_net_1\, \ADJ_Q[1]_net_1\, \Q[2]_net_1\, 
        \ADJ_Q[2]_net_1\, \Q[3]_net_1\, \ADJ_Q[3]_net_1\, 
        \Q[4]_net_1\, \ADJ_Q[4]_net_1\, \Q[5]_net_1\, 
        \ADJ_Q[5]_net_1\, \Q[6]_net_1\, \ADJ_Q[6]_net_1\, 
        \Q[7]_net_1\, \ADJ_Q[7]_net_1\, \Q[8]_net_1\, 
        \ADJ_Q[8]_net_1\, \Q[9]_net_1\, \ADJ_Q[9]_net_1\, 
        \Q[10]_net_1\, \ADJ_Q[10]_net_1\, \Q[11]_net_1\, 
        \ADJ_Q[11]_net_1\, \Q[12]_net_1\, \ADJ_Q[12]_net_1\, 
        \Q[13]_net_1\, \ADJ_Q[13]_net_1\, \Q[14]_net_1\, 
        \ADJ_Q[14]_net_1\, \ARB_WRD_40M_FIXED[0]_net_1\, 
        \ARB_WRD_40M_FIXED[1]_net_1\, 
        \ARB_WRD_40M_FIXED[2]_net_1\, 
        \ARB_WRD_40M_FIXED[3]_net_1\, 
        \ARB_WRD_40M_FIXED[4]_net_1\, 
        \ARB_WRD_40M_FIXED[5]_net_1\, 
        \ARB_WRD_40M_FIXED[6]_net_1\, 
        \ARB_WRD_40M_FIXED[7]_net_1\, 
        \ARB_WRD_40M_FIXED[8]_net_1\, 
        \ARB_WRD_40M_FIXED[9]_net_1\, 
        \ARB_WRD_40M_FIXED[10]_net_1\, 
        \ARB_WRD_40M_FIXED[11]_net_1\, 
        \ARB_WRD_40M_FIXED[12]_net_1\, 
        \ARB_WRD_40M_FIXED[13]_net_1\, 
        \ARB_WRD_40M_FIXED[14]_net_1\, \GND\, \VCC\ : std_logic;

begin 


    \RECD_SER_WORD_RNO[5]\ : MX2
      port map(A => N_38, B => N_39, S => BIT_OS_SEL_1_0, Y => 
        \N_RECD_SER_WORD[5]\);
    
    \ARB_WRD_40M_FIXED[9]\ : DFN1C0
      port map(D => \Q[9]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[9]_net_1\);
    
    \ADJ_Q[4]\ : DFN1C0
      port map(D => \ADJ_Q[2]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[4]_net_1\);
    
    \ARB_BYTE[6]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[6]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[6]_net_1\);
    
    ADJ_SER_IN_F_1DEL : DFN1C0
      port map(D => \ADJ_SER_IN_F_0DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_F_1DEL\);
    
    \ARB_BYTE[0]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[0]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[0]_net_1\);
    
    \Q[11]\ : DFN1C0
      port map(D => \ADJ_Q[11]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[11]_net_1\);
    
    \ADJ_Q[8]\ : DFN1C0
      port map(D => \ADJ_Q[6]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[8]_net_1\);
    
    \ADJ_Q[6]\ : DFN1C0
      port map(D => \ADJ_Q[4]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[6]_net_1\);
    
    \ARB_BYTE_RNI7K37[4]\ : MX2
      port map(A => \ARB_BYTE[4]_net_1\, B => \ARB_BYTE[8]_net_1\, 
        S => BIT_OS_SEL_7_0, Y => N_21);
    
    \ADJ_Q[12]\ : DFN1C0
      port map(D => \ADJ_Q[10]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[12]_net_1\);
    
    \RECD_SER_WORD_RNO_1[0]\ : MX2
      port map(A => \ARB_BYTE[0]_net_1\, B => \ARB_BYTE[4]_net_1\, 
        S => BIT_OS_SEL_7_0, Y => N_17);
    
    \ARB_BYTE_RNINKVI[1]\ : MX2
      port map(A => N_18, B => N_20, S => BIT_OS_SEL_6_0, Y => 
        N_34);
    
    \Q[1]\ : DFN1C0
      port map(D => \ADJ_Q[1]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[1]_net_1\);
    
    \ARB_BYTE_RNI5I37[3]\ : MX2
      port map(A => \ARB_BYTE[3]_net_1\, B => \ARB_BYTE[7]_net_1\, 
        S => BIT_OS_SEL_7_0, Y => N_20);
    
    \ARB_BYTE_RNI41JT[6]\ : MX2
      port map(A => N_23, B => N_31, S => BIT_OS_SEL_0_d0, Y => 
        N_39);
    
    \ARB_BYTE[4]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[4]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[4]_net_1\);
    
    \ADJ_Q[2]\ : DFN1C0
      port map(D => \ADJ_Q[0]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[2]_net_1\);
    
    \RECD_SER_WORD_RNO_1[7]\ : MX2
      port map(A => \ARB_BYTE[10]_net_1\, B => 
        \ARB_BYTE[14]_net_1\, S => BIT_OS_SEL_0(2), Y => N_56);
    
    \RECD_SER_WORD[4]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[4]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_3(4));
    
    \Q[5]\ : DFN1C0
      port map(D => \ADJ_Q[5]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[5]_net_1\);
    
    \ADJ_Q[11]\ : DFN1C0
      port map(D => \ADJ_Q[9]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[11]_net_1\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \ADJ_Q[3]\ : DFN1C0
      port map(D => \ADJ_Q[1]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[3]_net_1\);
    
    \Q[10]\ : DFN1C0
      port map(D => \ADJ_Q[10]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[10]_net_1\);
    
    \ARB_WRD_40M_FIXED[6]\ : DFN1C0
      port map(D => \Q[6]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[6]_net_1\);
    
    \ARB_BYTE_RNIPSRP[5]\ : MX2
      port map(A => N_22, B => N_24, S => BIT_OS_SEL_0_d0, Y => 
        N_38);
    
    \ARB_WRD_40M_FIXED[1]\ : DFN1C0
      port map(D => \Q[1]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[1]_net_1\);
    
    \RECD_SER_WORD[3]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[3]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_3(3));
    
    \RECD_SER_WORD[0]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[0]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_3(0));
    
    \ARB_BYTE_RNIA1NM[4]\ : MX2
      port map(A => N_21, B => N_23, S => BIT_OS_SEL_6_0, Y => 
        N_37);
    
    \RECD_SER_WORD_RNO[3]\ : MX2
      port map(A => N_36, B => N_37, S => BIT_OS_SEL_1_0, Y => 
        \N_RECD_SER_WORD[3]\);
    
    \Q[0]\ : DFN1C0
      port map(D => \ADJ_Q[0]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[0]_net_1\);
    
    \ARB_BYTE_RNIMSQA[12]\ : MX2
      port map(A => \ARB_BYTE[8]_net_1\, B => 
        \ARB_BYTE[12]_net_1\, S => BIT_OS_SEL_7_0, Y => N_31);
    
    \RECD_SER_WORD_RNO_0[7]\ : MX2
      port map(A => N_31, B => N_56, S => BIT_OS_SEL_0(1), Y => 
        N_64);
    
    \Q[7]\ : DFN1C0
      port map(D => \ADJ_Q[7]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[7]_net_1\);
    
    \ARB_BYTE[14]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[14]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[14]_net_1\);
    
    \ARB_WRD_40M_FIXED[2]\ : DFN1C0
      port map(D => \Q[2]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[2]_net_1\);
    
    \ARB_WRD_40M_FIXED[14]\ : DFN1C0
      port map(D => \Q[14]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[14]_net_1\);
    
    \RECD_SER_WORD_RNO[2]\ : MX2
      port map(A => N_35, B => N_36, S => BIT_OS_SEL_1_0, Y => 
        \N_RECD_SER_WORD[2]\);
    
    \ARB_BYTE[2]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[2]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[2]_net_1\);
    
    \ARB_BYTE_RNI3G37[2]\ : MX2
      port map(A => \ARB_BYTE[2]_net_1\, B => \ARB_BYTE[6]_net_1\, 
        S => BIT_OS_SEL_7_0, Y => N_19);
    
    \ADJ_Q[7]\ : DFN1C0
      port map(D => \ADJ_Q[5]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[7]_net_1\);
    
    \ARB_BYTE[8]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[8]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[8]_net_1\);
    
    \RECD_SER_WORD[5]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[5]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_3(5));
    
    \ARB_BYTE_RNIIOQA[6]\ : MX2
      port map(A => \ARB_BYTE[6]_net_1\, B => 
        \ARB_BYTE[10]_net_1\, S => BIT_OS_SEL_7_0, Y => N_23);
    
    \ARB_BYTE[12]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[12]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[12]_net_1\);
    
    \RECD_SER_WORD[1]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[1]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_3(1));
    
    \Q[3]\ : DFN1C0
      port map(D => \ADJ_Q[3]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[3]_net_1\);
    
    ADJ_SER_IN_F_0DEL : DFN1C0
      port map(D => ELK_IN_F, CLK => CCC_160M_ADJ, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_F_0DEL\);
    
    \RECD_SER_WORD_RNO[7]\ : MX2
      port map(A => N_40, B => N_64, S => BIT_OS_SEL_1_0, Y => 
        \N_RECD_SER_WORD[7]\);
    
    \RECD_SER_WORD_RNO[1]\ : MX2
      port map(A => N_34, B => N_35, S => BIT_OS_SEL_1_0, Y => 
        \N_RECD_SER_WORD[1]\);
    
    \ARB_WRD_40M_FIXED[4]\ : DFN1C0
      port map(D => \Q[4]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[4]_net_1\);
    
    \RECD_SER_WORD_RNO[0]\ : MX2
      port map(A => N_33, B => N_34, S => BIT_OS_SEL_1_0, Y => 
        \N_RECD_SER_WORD[0]\);
    
    \Q[6]\ : DFN1C0
      port map(D => \ADJ_Q[6]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[6]_net_1\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \ARB_WRD_40M_FIXED[8]\ : DFN1C0
      port map(D => \Q[8]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[8]_net_1\);
    
    \ARB_BYTE[11]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[11]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[11]_net_1\);
    
    \Q[9]\ : DFN1C0
      port map(D => \ADJ_Q[9]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[9]_net_1\);
    
    \Q[14]\ : DFN1C0
      port map(D => \ADJ_Q[14]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[14]_net_1\);
    
    \ARB_BYTE_RNI85JT[13]\ : MX2
      port map(A => N_24, B => N_32, S => BIT_OS_SEL_0_d0, Y => 
        N_40);
    
    ADJ_SER_IN_R_0DEL : DFN1C0
      port map(D => ELK_IN_R, CLK => CCC_160M_ADJ, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_R_0DEL\);
    
    \Q[13]\ : DFN1C0
      port map(D => \ADJ_Q[13]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[13]_net_1\);
    
    \ARB_BYTE[9]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[9]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[9]_net_1\);
    
    ADJ_SER_IN_R_1DEL : DFN1C0
      port map(D => \ADJ_SER_IN_R_0DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_R_1DEL\);
    
    \ARB_BYTE[10]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[10]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[10]_net_1\);
    
    \ADJ_Q[9]\ : DFN1C0
      port map(D => \ADJ_Q[7]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[9]_net_1\);
    
    \RECD_SER_WORD[7]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[7]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_3(7));
    
    \ARB_WRD_40M_FIXED[5]\ : DFN1C0
      port map(D => \Q[5]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[5]_net_1\);
    
    \ARB_WRD_40M_FIXED[12]\ : DFN1C0
      port map(D => \Q[12]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[12]_net_1\);
    
    \ARB_WRD_40M_FIXED[11]\ : DFN1C0
      port map(D => \Q[11]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[11]_net_1\);
    
    \ARB_BYTE_RNIVSVI[3]\ : MX2
      port map(A => N_20, B => N_22, S => BIT_OS_SEL_6_0, Y => 
        N_36);
    
    \ARB_BYTE_RNI9M37[5]\ : MX2
      port map(A => \ARB_BYTE[5]_net_1\, B => \ARB_BYTE[9]_net_1\, 
        S => BIT_OS_SEL_7_0, Y => N_22);
    
    \ARB_WRD_40M_FIXED[0]\ : DFN1C0
      port map(D => \Q[0]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[0]_net_1\);
    
    \ADJ_Q[10]\ : DFN1C0
      port map(D => \ADJ_Q[8]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[10]_net_1\);
    
    \Q[2]\ : DFN1C0
      port map(D => \ADJ_Q[2]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[2]_net_1\);
    
    \ARB_BYTE_RNI1E37[1]\ : MX2
      port map(A => \ARB_BYTE[1]_net_1\, B => \ARB_BYTE[5]_net_1\, 
        S => BIT_OS_SEL_7_0, Y => N_18);
    
    \ADJ_Q[1]\ : DFN1C0
      port map(D => \ADJ_SER_IN_F_1DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[1]_net_1\);
    
    \RECD_SER_WORD[6]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[6]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_3(6));
    
    \RECD_SER_WORD[2]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[2]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_3(2));
    
    \ADJ_Q[13]\ : DFN1C0
      port map(D => \ADJ_Q[11]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[13]_net_1\);
    
    \Q[8]\ : DFN1C0
      port map(D => \ADJ_Q[8]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[8]_net_1\);
    
    \ARB_BYTE_RNIOUQA[13]\ : MX2
      port map(A => \ARB_BYTE[9]_net_1\, B => 
        \ARB_BYTE[13]_net_1\, S => BIT_OS_SEL_7_0, Y => N_32);
    
    \ARB_BYTE[5]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[5]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[5]_net_1\);
    
    \ADJ_Q[14]\ : DFN1C0
      port map(D => \ADJ_Q[12]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[14]_net_1\);
    
    \RECD_SER_WORD_RNO[4]\ : MX2
      port map(A => N_37, B => N_38, S => BIT_OS_SEL_1_0, Y => 
        \N_RECD_SER_WORD[4]\);
    
    \Q[12]\ : DFN1C0
      port map(D => \ADJ_Q[12]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[12]_net_1\);
    
    \ARB_BYTE[13]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[13]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[13]_net_1\);
    
    \ARB_WRD_40M_FIXED[3]\ : DFN1C0
      port map(D => \Q[3]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[3]_net_1\);
    
    \ARB_BYTE[7]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[7]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[7]_net_1\);
    
    \RECD_SER_WORD_RNO_0[0]\ : MX2
      port map(A => N_17, B => N_19, S => BIT_OS_SEL_6_0, Y => 
        N_33);
    
    \Q[4]\ : DFN1C0
      port map(D => \ADJ_Q[4]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[4]_net_1\);
    
    \ARB_WRD_40M_FIXED[7]\ : DFN1C0
      port map(D => \Q[7]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[7]_net_1\);
    
    \RECD_SER_WORD_RNO[6]\ : MX2
      port map(A => N_39, B => N_40, S => BIT_OS_SEL_1_0, Y => 
        \N_RECD_SER_WORD[6]\);
    
    \ARB_BYTE[3]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[3]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[3]_net_1\);
    
    \ADJ_Q[5]\ : DFN1C0
      port map(D => \ADJ_Q[3]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[5]_net_1\);
    
    \ARB_BYTE[1]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[1]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[1]_net_1\);
    
    \ARB_BYTE_RNIROVI[2]\ : MX2
      port map(A => N_19, B => N_21, S => BIT_OS_SEL_6_0, Y => 
        N_35);
    
    \ARB_WRD_40M_FIXED[13]\ : DFN1C0
      port map(D => \Q[13]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[13]_net_1\);
    
    \ADJ_Q[0]\ : DFN1C0
      port map(D => \ADJ_SER_IN_R_1DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[0]_net_1\);
    
    \ARB_BYTE_RNIKQQA[11]\ : MX2
      port map(A => \ARB_BYTE[7]_net_1\, B => 
        \ARB_BYTE[11]_net_1\, S => BIT_OS_SEL_7_0, Y => N_24);
    
    \ARB_WRD_40M_FIXED[10]\ : DFN1C0
      port map(D => \Q[10]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[10]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SER320M_3_34_3 is

    port( ELK_TX_DAT                 : in    std_logic_vector(7 downto 0);
          MASTER_SALT_POR_B_i_0_i_12 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_16 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_3  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_2  : in    std_logic;
          ELK_OUT_R_i_0              : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_5  : in    std_logic;
          ELK_OUT_F_i_0              : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_8  : in    std_logic;
          CLK_40M_GL                 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_14 : in    std_logic;
          CCC_160M_FXD               : in    std_logic
        );

end SER320M_3_34_3;

architecture DEF_ARCH of SER320M_3_34_3 is 

  component DFI1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          QN  : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component DFN1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

    signal SER_OUT_RI_i, \SER_CMD_WORD_R[3]_net_1\, SER_OUT_FI_i, 
        \SER_CMD_WORD_F[3]_net_1\, \N_SER_CMD_WORD_R[0]\, 
        \START_RISE\, \N_SER_CMD_WORD_F[0]\, 
        \N_SER_CMD_WORD_R[3]\, \SER_CMD_WORD_R[2]_net_1\, 
        \N_SER_CMD_WORD_R[2]\, \SER_CMD_WORD_R[1]_net_1\, 
        \N_SER_CMD_WORD_R[1]\, \SER_CMD_WORD_R[0]_net_1\, 
        \N_SER_CMD_WORD_F[3]\, \SER_CMD_WORD_F[2]_net_1\, 
        \N_SER_CMD_WORD_F[2]\, \SER_CMD_WORD_F[1]_net_1\, 
        \N_SER_CMD_WORD_F[1]\, \SER_CMD_WORD_F[0]_net_1\, 
        N_START_RISE, \CLK40M_GEN_DEL0\, \GND\, \VCC\
         : std_logic;

begin 


    SER_OUT_FI : DFI1C0
      port map(D => \SER_CMD_WORD_F[3]_net_1\, CLK => 
        CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_14, QN => 
        SER_OUT_FI_i);
    
    \SER_CMD_WORD_F[3]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[3]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_16, Q => 
        \SER_CMD_WORD_F[3]_net_1\);
    
    \SER_CMD_WORD_R[1]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[1]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_12, Q => 
        \SER_CMD_WORD_R[1]_net_1\);
    
    \SER_CMD_WORD_R[2]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[2]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_12, Q => 
        \SER_CMD_WORD_R[2]_net_1\);
    
    \SER_CMD_WORD_R_RNO[3]\ : MX2
      port map(A => \SER_CMD_WORD_R[2]_net_1\, B => ELK_TX_DAT(7), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_R[3]\);
    
    \SER_CMD_WORD_R_RNO[0]\ : NOR2B
      port map(A => \START_RISE\, B => ELK_TX_DAT(1), Y => 
        \N_SER_CMD_WORD_R[0]\);
    
    \SER_CMD_WORD_F[0]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[0]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_16, Q => 
        \SER_CMD_WORD_F[0]_net_1\);
    
    \SER_CMD_WORD_R_RNO[1]\ : MX2
      port map(A => \SER_CMD_WORD_R[0]_net_1\, B => ELK_TX_DAT(3), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_R[1]\);
    
    \SER_CMD_WORD_F_RNO[2]\ : MX2
      port map(A => \SER_CMD_WORD_F[1]_net_1\, B => ELK_TX_DAT(4), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_F[2]\);
    
    \SER_CMD_WORD_F_RNO[3]\ : MX2
      port map(A => \SER_CMD_WORD_F[2]_net_1\, B => ELK_TX_DAT(6), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_F[3]\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    CLK40M_GEN_DEL0 : DFN1C0
      port map(D => CLK_40M_GL, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_8, Q => \CLK40M_GEN_DEL0\);
    
    SER_OUT_RI : DFI1C0
      port map(D => \SER_CMD_WORD_R[3]_net_1\, CLK => 
        CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_14, QN => 
        SER_OUT_RI_i);
    
    \SER_CMD_WORD_F[2]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[2]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_16, Q => 
        \SER_CMD_WORD_F[2]_net_1\);
    
    \SER_CMD_WORD_F_RNO[1]\ : MX2
      port map(A => \SER_CMD_WORD_F[0]_net_1\, B => ELK_TX_DAT(2), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_F[1]\);
    
    \SER_CMD_WORD_R[0]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[0]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_12, Q => 
        \SER_CMD_WORD_R[0]_net_1\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    START_RISE : DFN1C0
      port map(D => N_START_RISE, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_3, Q => \START_RISE\);
    
    \SER_CMD_WORD_R[3]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[3]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_12, Q => 
        \SER_CMD_WORD_R[3]_net_1\);
    
    \SER_CMD_WORD_F_RNO[0]\ : NOR2B
      port map(A => \START_RISE\, B => ELK_TX_DAT(0), Y => 
        \N_SER_CMD_WORD_F[0]\);
    
    SER_OUT_RDEL : DFN1P0
      port map(D => SER_OUT_RI_i, CLK => CCC_160M_FXD, PRE => 
        MASTER_SALT_POR_B_i_0_i_2, Q => ELK_OUT_R_i_0);
    
    \SER_CMD_WORD_F[1]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[1]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_16, Q => 
        \SER_CMD_WORD_F[1]_net_1\);
    
    START_RISE_RNO : NOR2B
      port map(A => \CLK40M_GEN_DEL0\, B => CLK_40M_GL, Y => 
        N_START_RISE);
    
    \SER_CMD_WORD_R_RNO[2]\ : MX2
      port map(A => \SER_CMD_WORD_R[1]_net_1\, B => ELK_TX_DAT(5), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_R[2]\);
    
    SER_OUT_FDEL : DFN1P0
      port map(D => SER_OUT_FI_i, CLK => CCC_160M_FXD, PRE => 
        MASTER_SALT_POR_B_i_0_i_5, Q => ELK_OUT_F_i_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity DDR_BIDIR_LVDS_DUAL_CLK_3 is

    port( DCB_SALT_SEL_c_i : in    std_logic;
          ELK3_DAT_P       : inout std_logic := 'Z';
          ELK3_DAT_N       : inout std_logic := 'Z';
          ELK_OUT_R_i_0    : in    std_logic;
          ELK_OUT_F_i_0    : in    std_logic;
          CCC_160M_FXD     : in    std_logic;
          CCC_160M_ADJ     : in    std_logic;
          ELK_IN_DDR_F_i   : out   std_logic;
          ELK_IN_DDR_R_i   : out   std_logic
        );

end DDR_BIDIR_LVDS_DUAL_CLK_3;

architecture DEF_ARCH of DDR_BIDIR_LVDS_DUAL_CLK_3 is 

  component INV
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DDR_REG
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          QR  : out   std_logic;
          QF  : out   std_logic
        );
  end component;

  component DDR_OUT
    port( DR  : in    std_logic := 'U';
          DF  : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component BIBUF_LVDS
    port( PADP : inout   std_logic;
          PADN : inout   std_logic;
          D    : in    std_logic := 'U';
          E    : in    std_logic := 'U';
          Y    : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal ELK_IN_DDR_R, ELK_IN_DDR_F, 
        DDR_BIDIR_LVDS_DUAL_CLK_3_GND, BIBUF_LVDS_0_Y, 
        DDR_OUT_0_Q, \VCC\ : std_logic;

begin 


    DDR_REG_0_RNI992A_0 : INV
      port map(A => ELK_IN_DDR_R, Y => ELK_IN_DDR_R_i);
    
    DDR_REG_0_RNI992A : INV
      port map(A => ELK_IN_DDR_F, Y => ELK_IN_DDR_F_i);
    
    DDR_REG_0 : DDR_REG
      port map(D => BIBUF_LVDS_0_Y, CLK => CCC_160M_ADJ, CLR => 
        DDR_BIDIR_LVDS_DUAL_CLK_3_GND, QR => ELK_IN_DDR_R, QF => 
        ELK_IN_DDR_F);
    
    DDR_OUT_0 : DDR_OUT
      port map(DR => ELK_OUT_R_i_0, DF => ELK_OUT_F_i_0, CLK => 
        CCC_160M_FXD, CLR => DDR_BIDIR_LVDS_DUAL_CLK_3_GND, Q => 
        DDR_OUT_0_Q);
    
    BIBUF_LVDS_0 : BIBUF_LVDS
      port map(PADP => ELK3_DAT_P, PADN => ELK3_DAT_N, D => 
        DDR_OUT_0_Q, E => DCB_SALT_SEL_c_i, Y => BIBUF_LVDS_0_Y);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    GND_i : GND
      port map(Y => DDR_BIDIR_LVDS_DUAL_CLK_3_GND);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SYNC_DAT_SEL_3 is

    port( ELK_TX_DAT                 : out   std_logic_vector(7 downto 0);
          PATT_ELK_DAT_3             : in    std_logic_vector(7 downto 0);
          OP_MODE_c_5_0              : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_15 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_14 : in    std_logic;
          CLK_40M_GL                 : in    std_logic
        );

end SYNC_DAT_SEL_3;

architecture DEF_ARCH of SYNC_DAT_SEL_3 is 

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \N_SERDAT[0]\, \N_SERDAT[1]\, \N_SERDAT[2]\, 
        \N_SERDAT[3]\, \N_SERDAT[4]\, \N_SERDAT[5]\, 
        \N_SERDAT[6]\, \N_SERDAT[7]\, \GND\, \VCC\ : std_logic;

begin 


    \SERDAT_RNO[4]\ : NOR2A
      port map(A => PATT_ELK_DAT_3(4), B => OP_MODE_c_5_0, Y => 
        \N_SERDAT[4]\);
    
    \SERDAT_RNO[0]\ : NOR2A
      port map(A => PATT_ELK_DAT_3(0), B => OP_MODE_c_5_0, Y => 
        \N_SERDAT[0]\);
    
    \SERDAT[6]\ : DFN1C0
      port map(D => \N_SERDAT[6]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_15, Q => ELK_TX_DAT(6));
    
    \SERDAT[4]\ : DFN1C0
      port map(D => \N_SERDAT[4]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_15, Q => ELK_TX_DAT(4));
    
    \SERDAT_RNO[7]\ : OR2
      port map(A => PATT_ELK_DAT_3(7), B => OP_MODE_c_5_0, Y => 
        \N_SERDAT[7]\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \SERDAT_RNO[3]\ : OR2
      port map(A => PATT_ELK_DAT_3(3), B => OP_MODE_c_5_0, Y => 
        \N_SERDAT[3]\);
    
    \SERDAT_RNO[2]\ : OR2
      port map(A => PATT_ELK_DAT_3(2), B => OP_MODE_c_5_0, Y => 
        \N_SERDAT[2]\);
    
    \SERDAT[5]\ : DFN1C0
      port map(D => \N_SERDAT[5]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_15, Q => ELK_TX_DAT(5));
    
    \SERDAT[7]\ : DFN1C0
      port map(D => \N_SERDAT[7]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_15, Q => ELK_TX_DAT(7));
    
    GND_i : GND
      port map(Y => \GND\);
    
    \SERDAT_RNO[5]\ : NOR2A
      port map(A => PATT_ELK_DAT_3(5), B => OP_MODE_c_5_0, Y => 
        \N_SERDAT[5]\);
    
    \SERDAT[0]\ : DFN1C0
      port map(D => \N_SERDAT[0]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_14, Q => ELK_TX_DAT(0));
    
    \SERDAT_RNO[6]\ : NOR2A
      port map(A => PATT_ELK_DAT_3(6), B => OP_MODE_c_5_0, Y => 
        \N_SERDAT[6]\);
    
    \SERDAT[1]\ : DFN1C0
      port map(D => \N_SERDAT[1]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_15, Q => ELK_TX_DAT(1));
    
    \SERDAT_RNO[1]\ : OR2
      port map(A => PATT_ELK_DAT_3(1), B => OP_MODE_c_5_0, Y => 
        \N_SERDAT[1]\);
    
    \SERDAT[3]\ : DFN1C0
      port map(D => \N_SERDAT[3]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_15, Q => ELK_TX_DAT(3));
    
    \SERDAT[2]\ : DFN1C0
      port map(D => \N_SERDAT[2]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_15, Q => ELK_TX_DAT(2));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity ELINK_SLAVE_INV_2_0 is

    port( BIT_OS_SEL_7_0             : in    std_logic;
          BIT_OS_SEL_6_0             : in    std_logic;
          BIT_OS_SEL_0_d0            : in    std_logic;
          BIT_OS_SEL_0               : in    std_logic_vector(2 downto 1);
          BIT_OS_SEL_1_0             : in    std_logic;
          ELK_RX_SER_WORD_3          : out   std_logic_vector(7 downto 0);
          OP_MODE_c_5_0              : in    std_logic;
          PATT_ELK_DAT_3             : in    std_logic_vector(7 downto 0);
          MASTER_DCB_POR_B_i_0_i     : in    std_logic;
          ELK3_DAT_N                 : inout std_logic := 'Z';
          ELK3_DAT_P                 : inout std_logic := 'Z';
          DCB_SALT_SEL_c_i           : in    std_logic;
          CCC_160M_FXD               : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_8  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_5  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_2  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_3  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_16 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_12 : in    std_logic;
          CLK_40M_GL                 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_14 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_15 : in    std_logic;
          DEV_RST_B_c                : in    std_logic;
          CCC_160M_ADJ               : in    std_logic
        );

end ELINK_SLAVE_INV_2_0;

architecture DEF_ARCH of ELINK_SLAVE_INV_2_0 is 

  component SLAVE_DES320S_1_17_1
    port( ELK_RX_SER_WORD_3      : out   std_logic_vector(7 downto 0);
          BIT_OS_SEL_1_0         : in    std_logic := 'U';
          BIT_OS_SEL_0           : in    std_logic_vector(2 downto 1) := (others => 'U');
          BIT_OS_SEL_0_d0        : in    std_logic := 'U';
          BIT_OS_SEL_6_0         : in    std_logic := 'U';
          BIT_OS_SEL_7_0         : in    std_logic := 'U';
          CLK_40M_GL             : in    std_logic := 'U';
          CCC_160M_FXD           : in    std_logic := 'U';
          ELK_IN_R               : in    std_logic := 'U';
          ELK_IN_F               : in    std_logic := 'U';
          MASTER_DCB_POR_B_i_0_i : in    std_logic := 'U';
          CCC_160M_ADJ           : in    std_logic := 'U'
        );
  end component;

  component SER320M_3_34_3
    port( ELK_TX_DAT                 : in    std_logic_vector(7 downto 0) := (others => 'U');
          MASTER_SALT_POR_B_i_0_i_12 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_16 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_3  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_2  : in    std_logic := 'U';
          ELK_OUT_R_i_0              : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_5  : in    std_logic := 'U';
          ELK_OUT_F_i_0              : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_8  : in    std_logic := 'U';
          CLK_40M_GL                 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_14 : in    std_logic := 'U';
          CCC_160M_FXD               : in    std_logic := 'U'
        );
  end component;

  component DDR_BIDIR_LVDS_DUAL_CLK_3
    port( DCB_SALT_SEL_c_i : in    std_logic := 'U';
          ELK3_DAT_P       : inout   std_logic;
          ELK3_DAT_N       : inout   std_logic;
          ELK_OUT_R_i_0    : in    std_logic := 'U';
          ELK_OUT_F_i_0    : in    std_logic := 'U';
          CCC_160M_FXD     : in    std_logic := 'U';
          CCC_160M_ADJ     : in    std_logic := 'U';
          ELK_IN_DDR_F_i   : out   std_logic;
          ELK_IN_DDR_R_i   : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component SYNC_DAT_SEL_3
    port( ELK_TX_DAT                 : out   std_logic_vector(7 downto 0);
          PATT_ELK_DAT_3             : in    std_logic_vector(7 downto 0) := (others => 'U');
          OP_MODE_c_5_0              : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_15 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_14 : in    std_logic := 'U';
          CLK_40M_GL                 : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \ELK_IN_F\, ELK_IN_DDR_F_i, \ELK_IN_R\, 
        ELK_IN_DDR_R_i, \ELK_TX_DAT[0]\, \ELK_TX_DAT[1]\, 
        \ELK_TX_DAT[2]\, \ELK_TX_DAT[3]\, \ELK_TX_DAT[4]\, 
        \ELK_TX_DAT[5]\, \ELK_TX_DAT[6]\, \ELK_TX_DAT[7]\, 
        ELK_OUT_R_i_0, ELK_OUT_F_i_0, \GND\, \VCC\ : std_logic;

    for all : SLAVE_DES320S_1_17_1
	Use entity work.SLAVE_DES320S_1_17_1(DEF_ARCH);
    for all : SER320M_3_34_3
	Use entity work.SER320M_3_34_3(DEF_ARCH);
    for all : DDR_BIDIR_LVDS_DUAL_CLK_3
	Use entity work.DDR_BIDIR_LVDS_DUAL_CLK_3(DEF_ARCH);
    for all : SYNC_DAT_SEL_3
	Use entity work.SYNC_DAT_SEL_3(DEF_ARCH);
begin 


    U_SLAVE_1ELK : SLAVE_DES320S_1_17_1
      port map(ELK_RX_SER_WORD_3(7) => ELK_RX_SER_WORD_3(7), 
        ELK_RX_SER_WORD_3(6) => ELK_RX_SER_WORD_3(6), 
        ELK_RX_SER_WORD_3(5) => ELK_RX_SER_WORD_3(5), 
        ELK_RX_SER_WORD_3(4) => ELK_RX_SER_WORD_3(4), 
        ELK_RX_SER_WORD_3(3) => ELK_RX_SER_WORD_3(3), 
        ELK_RX_SER_WORD_3(2) => ELK_RX_SER_WORD_3(2), 
        ELK_RX_SER_WORD_3(1) => ELK_RX_SER_WORD_3(1), 
        ELK_RX_SER_WORD_3(0) => ELK_RX_SER_WORD_3(0), 
        BIT_OS_SEL_1_0 => BIT_OS_SEL_1_0, BIT_OS_SEL_0(2) => 
        BIT_OS_SEL_0(2), BIT_OS_SEL_0(1) => BIT_OS_SEL_0(1), 
        BIT_OS_SEL_0_d0 => BIT_OS_SEL_0_d0, BIT_OS_SEL_6_0 => 
        BIT_OS_SEL_6_0, BIT_OS_SEL_7_0 => BIT_OS_SEL_7_0, 
        CLK_40M_GL => CLK_40M_GL, CCC_160M_FXD => CCC_160M_FXD, 
        ELK_IN_R => \ELK_IN_R\, ELK_IN_F => \ELK_IN_F\, 
        MASTER_DCB_POR_B_i_0_i => MASTER_DCB_POR_B_i_0_i, 
        CCC_160M_ADJ => CCC_160M_ADJ);
    
    U_ELK1_CMD_TX : SER320M_3_34_3
      port map(ELK_TX_DAT(7) => \ELK_TX_DAT[7]\, ELK_TX_DAT(6)
         => \ELK_TX_DAT[6]\, ELK_TX_DAT(5) => \ELK_TX_DAT[5]\, 
        ELK_TX_DAT(4) => \ELK_TX_DAT[4]\, ELK_TX_DAT(3) => 
        \ELK_TX_DAT[3]\, ELK_TX_DAT(2) => \ELK_TX_DAT[2]\, 
        ELK_TX_DAT(1) => \ELK_TX_DAT[1]\, ELK_TX_DAT(0) => 
        \ELK_TX_DAT[0]\, MASTER_SALT_POR_B_i_0_i_12 => 
        MASTER_SALT_POR_B_i_0_i_12, MASTER_SALT_POR_B_i_0_i_16
         => MASTER_SALT_POR_B_i_0_i_16, MASTER_SALT_POR_B_i_0_i_3
         => MASTER_SALT_POR_B_i_0_i_3, MASTER_SALT_POR_B_i_0_i_2
         => MASTER_SALT_POR_B_i_0_i_2, ELK_OUT_R_i_0 => 
        ELK_OUT_R_i_0, MASTER_SALT_POR_B_i_0_i_5 => 
        MASTER_SALT_POR_B_i_0_i_5, ELK_OUT_F_i_0 => ELK_OUT_F_i_0, 
        MASTER_SALT_POR_B_i_0_i_8 => MASTER_SALT_POR_B_i_0_i_8, 
        CLK_40M_GL => CLK_40M_GL, MASTER_SALT_POR_B_i_0_i_14 => 
        MASTER_SALT_POR_B_i_0_i_14, CCC_160M_FXD => CCC_160M_FXD);
    
    U_DDR_ELK1 : DDR_BIDIR_LVDS_DUAL_CLK_3
      port map(DCB_SALT_SEL_c_i => DCB_SALT_SEL_c_i, ELK3_DAT_P
         => ELK3_DAT_P, ELK3_DAT_N => ELK3_DAT_N, ELK_OUT_R_i_0
         => ELK_OUT_R_i_0, ELK_OUT_F_i_0 => ELK_OUT_F_i_0, 
        CCC_160M_FXD => CCC_160M_FXD, CCC_160M_ADJ => 
        CCC_160M_ADJ, ELK_IN_DDR_F_i => ELK_IN_DDR_F_i, 
        ELK_IN_DDR_R_i => ELK_IN_DDR_R_i);
    
    ELK_IN_F : DFN1C0
      port map(D => ELK_IN_DDR_F_i, CLK => CCC_160M_ADJ, CLR => 
        DEV_RST_B_c, Q => \ELK_IN_F\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    U_ELK1_SERDAT_SOURCE : SYNC_DAT_SEL_3
      port map(ELK_TX_DAT(7) => \ELK_TX_DAT[7]\, ELK_TX_DAT(6)
         => \ELK_TX_DAT[6]\, ELK_TX_DAT(5) => \ELK_TX_DAT[5]\, 
        ELK_TX_DAT(4) => \ELK_TX_DAT[4]\, ELK_TX_DAT(3) => 
        \ELK_TX_DAT[3]\, ELK_TX_DAT(2) => \ELK_TX_DAT[2]\, 
        ELK_TX_DAT(1) => \ELK_TX_DAT[1]\, ELK_TX_DAT(0) => 
        \ELK_TX_DAT[0]\, PATT_ELK_DAT_3(7) => PATT_ELK_DAT_3(7), 
        PATT_ELK_DAT_3(6) => PATT_ELK_DAT_3(6), PATT_ELK_DAT_3(5)
         => PATT_ELK_DAT_3(5), PATT_ELK_DAT_3(4) => 
        PATT_ELK_DAT_3(4), PATT_ELK_DAT_3(3) => PATT_ELK_DAT_3(3), 
        PATT_ELK_DAT_3(2) => PATT_ELK_DAT_3(2), PATT_ELK_DAT_3(1)
         => PATT_ELK_DAT_3(1), PATT_ELK_DAT_3(0) => 
        PATT_ELK_DAT_3(0), OP_MODE_c_5_0 => OP_MODE_c_5_0, 
        MASTER_SALT_POR_B_i_0_i_15 => MASTER_SALT_POR_B_i_0_i_15, 
        MASTER_SALT_POR_B_i_0_i_14 => MASTER_SALT_POR_B_i_0_i_14, 
        CLK_40M_GL => CLK_40M_GL);
    
    ELK_IN_R : DFN1C0
      port map(D => ELK_IN_DDR_R_i, CLK => CCC_160M_ADJ, CLR => 
        DEV_RST_B_c, Q => \ELK_IN_R\);
    
    GND_i : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity DPRT_512X9_SRAM_0 is

    port( ELINK_RWA_0         : in    std_logic;
          ELK_RX_SER_WORD_0   : in    std_logic_vector(7 downto 0);
          ELINK_DINA_0        : in    std_logic_vector(7 downto 0);
          ELINK_BLKA_0        : in    std_logic;
          ELKS_ADDRB          : in    std_logic_vector(7 downto 0);
          ELINK_ADDRA_0       : in    std_logic_vector(7 downto 0);
          PATT_ELK_DAT_0      : out   std_logic_vector(7 downto 0);
          ELINK_DOUTA_0       : out   std_logic_vector(7 downto 0);
          ELKS_RWB            : in    std_logic;
          P_USB_MASTER_EN_c_0 : in    std_logic;
          CLK_40M_GL          : in    std_logic;
          CLK60MHZ            : in    std_logic;
          ELKS_RAM_BLKB_EN    : in    std_logic
        );

end DPRT_512X9_SRAM_0;

architecture DEF_ARCH of DPRT_512X9_SRAM_0 is 

  component RAM4K9
    generic (MEMORYFILE:string := "");

    port( ADDRA11 : in    std_logic := 'U';
          ADDRA10 : in    std_logic := 'U';
          ADDRA9  : in    std_logic := 'U';
          ADDRA8  : in    std_logic := 'U';
          ADDRA7  : in    std_logic := 'U';
          ADDRA6  : in    std_logic := 'U';
          ADDRA5  : in    std_logic := 'U';
          ADDRA4  : in    std_logic := 'U';
          ADDRA3  : in    std_logic := 'U';
          ADDRA2  : in    std_logic := 'U';
          ADDRA1  : in    std_logic := 'U';
          ADDRA0  : in    std_logic := 'U';
          ADDRB11 : in    std_logic := 'U';
          ADDRB10 : in    std_logic := 'U';
          ADDRB9  : in    std_logic := 'U';
          ADDRB8  : in    std_logic := 'U';
          ADDRB7  : in    std_logic := 'U';
          ADDRB6  : in    std_logic := 'U';
          ADDRB5  : in    std_logic := 'U';
          ADDRB4  : in    std_logic := 'U';
          ADDRB3  : in    std_logic := 'U';
          ADDRB2  : in    std_logic := 'U';
          ADDRB1  : in    std_logic := 'U';
          ADDRB0  : in    std_logic := 'U';
          DINA8   : in    std_logic := 'U';
          DINA7   : in    std_logic := 'U';
          DINA6   : in    std_logic := 'U';
          DINA5   : in    std_logic := 'U';
          DINA4   : in    std_logic := 'U';
          DINA3   : in    std_logic := 'U';
          DINA2   : in    std_logic := 'U';
          DINA1   : in    std_logic := 'U';
          DINA0   : in    std_logic := 'U';
          DINB8   : in    std_logic := 'U';
          DINB7   : in    std_logic := 'U';
          DINB6   : in    std_logic := 'U';
          DINB5   : in    std_logic := 'U';
          DINB4   : in    std_logic := 'U';
          DINB3   : in    std_logic := 'U';
          DINB2   : in    std_logic := 'U';
          DINB1   : in    std_logic := 'U';
          DINB0   : in    std_logic := 'U';
          WIDTHA0 : in    std_logic := 'U';
          WIDTHA1 : in    std_logic := 'U';
          WIDTHB0 : in    std_logic := 'U';
          WIDTHB1 : in    std_logic := 'U';
          PIPEA   : in    std_logic := 'U';
          PIPEB   : in    std_logic := 'U';
          WMODEA  : in    std_logic := 'U';
          WMODEB  : in    std_logic := 'U';
          BLKA    : in    std_logic := 'U';
          BLKB    : in    std_logic := 'U';
          WENA    : in    std_logic := 'U';
          WENB    : in    std_logic := 'U';
          CLKA    : in    std_logic := 'U';
          CLKB    : in    std_logic := 'U';
          RESET   : in    std_logic := 'U';
          DOUTA8  : out   std_logic;
          DOUTA7  : out   std_logic;
          DOUTA6  : out   std_logic;
          DOUTA5  : out   std_logic;
          DOUTA4  : out   std_logic;
          DOUTA3  : out   std_logic;
          DOUTA2  : out   std_logic;
          DOUTA1  : out   std_logic;
          DOUTA0  : out   std_logic;
          DOUTB8  : out   std_logic;
          DOUTB7  : out   std_logic;
          DOUTB6  : out   std_logic;
          DOUTB5  : out   std_logic;
          DOUTB4  : out   std_logic;
          DOUTB3  : out   std_logic;
          DOUTB2  : out   std_logic;
          DOUTB1  : out   std_logic;
          DOUTB0  : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \DOUTA_1[8]\, \DOUTB_1[8]\, DPRT_512X9_SRAM_0_GND, 
        DPRT_512X9_SRAM_0_VCC : std_logic;

begin 


    DPRT_512X9_SRAM_R0C0 : RAM4K9
      generic map(MEMORYFILE => "DPRT_512X9_SRAM_R0C0.mem")

      port map(ADDRA11 => DPRT_512X9_SRAM_0_GND, ADDRA10 => 
        DPRT_512X9_SRAM_0_GND, ADDRA9 => DPRT_512X9_SRAM_0_GND, 
        ADDRA8 => DPRT_512X9_SRAM_0_GND, ADDRA7 => 
        ELINK_ADDRA_0(7), ADDRA6 => ELINK_ADDRA_0(6), ADDRA5 => 
        ELINK_ADDRA_0(5), ADDRA4 => ELINK_ADDRA_0(4), ADDRA3 => 
        ELINK_ADDRA_0(3), ADDRA2 => ELINK_ADDRA_0(2), ADDRA1 => 
        ELINK_ADDRA_0(1), ADDRA0 => ELINK_ADDRA_0(0), ADDRB11 => 
        DPRT_512X9_SRAM_0_GND, ADDRB10 => DPRT_512X9_SRAM_0_GND, 
        ADDRB9 => DPRT_512X9_SRAM_0_GND, ADDRB8 => 
        DPRT_512X9_SRAM_0_GND, ADDRB7 => ELKS_ADDRB(7), ADDRB6
         => ELKS_ADDRB(6), ADDRB5 => ELKS_ADDRB(5), ADDRB4 => 
        ELKS_ADDRB(4), ADDRB3 => ELKS_ADDRB(3), ADDRB2 => 
        ELKS_ADDRB(2), ADDRB1 => ELKS_ADDRB(1), ADDRB0 => 
        ELKS_ADDRB(0), DINA8 => DPRT_512X9_SRAM_0_GND, DINA7 => 
        ELINK_DINA_0(7), DINA6 => ELINK_DINA_0(6), DINA5 => 
        ELINK_DINA_0(5), DINA4 => ELINK_DINA_0(4), DINA3 => 
        ELINK_DINA_0(3), DINA2 => ELINK_DINA_0(2), DINA1 => 
        ELINK_DINA_0(1), DINA0 => ELINK_DINA_0(0), DINB8 => 
        DPRT_512X9_SRAM_0_GND, DINB7 => ELK_RX_SER_WORD_0(7), 
        DINB6 => ELK_RX_SER_WORD_0(6), DINB5 => 
        ELK_RX_SER_WORD_0(5), DINB4 => ELK_RX_SER_WORD_0(4), 
        DINB3 => ELK_RX_SER_WORD_0(3), DINB2 => 
        ELK_RX_SER_WORD_0(2), DINB1 => ELK_RX_SER_WORD_0(1), 
        DINB0 => ELK_RX_SER_WORD_0(0), WIDTHA0 => 
        DPRT_512X9_SRAM_0_VCC, WIDTHA1 => DPRT_512X9_SRAM_0_VCC, 
        WIDTHB0 => DPRT_512X9_SRAM_0_VCC, WIDTHB1 => 
        DPRT_512X9_SRAM_0_VCC, PIPEA => DPRT_512X9_SRAM_0_VCC, 
        PIPEB => DPRT_512X9_SRAM_0_VCC, WMODEA => 
        DPRT_512X9_SRAM_0_GND, WMODEB => DPRT_512X9_SRAM_0_GND, 
        BLKA => ELINK_BLKA_0, BLKB => ELKS_RAM_BLKB_EN, WENA => 
        ELINK_RWA_0, WENB => ELKS_RWB, CLKA => CLK60MHZ, CLKB => 
        CLK_40M_GL, RESET => P_USB_MASTER_EN_c_0, DOUTA8 => 
        \DOUTA_1[8]\, DOUTA7 => ELINK_DOUTA_0(7), DOUTA6 => 
        ELINK_DOUTA_0(6), DOUTA5 => ELINK_DOUTA_0(5), DOUTA4 => 
        ELINK_DOUTA_0(4), DOUTA3 => ELINK_DOUTA_0(3), DOUTA2 => 
        ELINK_DOUTA_0(2), DOUTA1 => ELINK_DOUTA_0(1), DOUTA0 => 
        ELINK_DOUTA_0(0), DOUTB8 => \DOUTB_1[8]\, DOUTB7 => 
        PATT_ELK_DAT_0(7), DOUTB6 => PATT_ELK_DAT_0(6), DOUTB5
         => PATT_ELK_DAT_0(5), DOUTB4 => PATT_ELK_DAT_0(4), 
        DOUTB3 => PATT_ELK_DAT_0(3), DOUTB2 => PATT_ELK_DAT_0(2), 
        DOUTB1 => PATT_ELK_DAT_0(1), DOUTB0 => PATT_ELK_DAT_0(0));
    
    VCC_i : VCC
      port map(Y => DPRT_512X9_SRAM_0_VCC);
    
    GND_i : GND
      port map(Y => DPRT_512X9_SRAM_0_GND);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity DPRT_512X9_SRAM_13 is

    port( ELINK_RWA_0         : in    std_logic;
          ELK_RX_SER_WORD_13  : in    std_logic_vector(7 downto 0);
          ELINK_DINA_13       : in    std_logic_vector(7 downto 0);
          ELINK_BLKA_0        : in    std_logic;
          ELKS_ADDRB_0_d0     : in    std_logic;
          ELKS_ADDRB_1        : in    std_logic;
          ELKS_ADDRB_3        : in    std_logic;
          ELKS_ADDRB_5        : in    std_logic;
          ELKS_ADDRB_7        : in    std_logic;
          ELKS_ADDRB_0_0      : in    std_logic;
          ELKS_ADDRB_0_2      : in    std_logic;
          ELKS_ADDRB_0_4      : in    std_logic;
          ELINK_ADDRA_13      : in    std_logic_vector(7 downto 0);
          PATT_ELK_DAT_13     : out   std_logic_vector(7 downto 0);
          ELINK_DOUTA_13      : out   std_logic_vector(7 downto 0);
          ELKS_RWB            : in    std_logic;
          P_USB_MASTER_EN_c_0 : in    std_logic;
          CLK_40M_GL          : in    std_logic;
          CLK60MHZ            : in    std_logic;
          ELKS_RAM_BLKB_EN    : in    std_logic
        );

end DPRT_512X9_SRAM_13;

architecture DEF_ARCH of DPRT_512X9_SRAM_13 is 

  component RAM4K9
    generic (MEMORYFILE:string := "");

    port( ADDRA11 : in    std_logic := 'U';
          ADDRA10 : in    std_logic := 'U';
          ADDRA9  : in    std_logic := 'U';
          ADDRA8  : in    std_logic := 'U';
          ADDRA7  : in    std_logic := 'U';
          ADDRA6  : in    std_logic := 'U';
          ADDRA5  : in    std_logic := 'U';
          ADDRA4  : in    std_logic := 'U';
          ADDRA3  : in    std_logic := 'U';
          ADDRA2  : in    std_logic := 'U';
          ADDRA1  : in    std_logic := 'U';
          ADDRA0  : in    std_logic := 'U';
          ADDRB11 : in    std_logic := 'U';
          ADDRB10 : in    std_logic := 'U';
          ADDRB9  : in    std_logic := 'U';
          ADDRB8  : in    std_logic := 'U';
          ADDRB7  : in    std_logic := 'U';
          ADDRB6  : in    std_logic := 'U';
          ADDRB5  : in    std_logic := 'U';
          ADDRB4  : in    std_logic := 'U';
          ADDRB3  : in    std_logic := 'U';
          ADDRB2  : in    std_logic := 'U';
          ADDRB1  : in    std_logic := 'U';
          ADDRB0  : in    std_logic := 'U';
          DINA8   : in    std_logic := 'U';
          DINA7   : in    std_logic := 'U';
          DINA6   : in    std_logic := 'U';
          DINA5   : in    std_logic := 'U';
          DINA4   : in    std_logic := 'U';
          DINA3   : in    std_logic := 'U';
          DINA2   : in    std_logic := 'U';
          DINA1   : in    std_logic := 'U';
          DINA0   : in    std_logic := 'U';
          DINB8   : in    std_logic := 'U';
          DINB7   : in    std_logic := 'U';
          DINB6   : in    std_logic := 'U';
          DINB5   : in    std_logic := 'U';
          DINB4   : in    std_logic := 'U';
          DINB3   : in    std_logic := 'U';
          DINB2   : in    std_logic := 'U';
          DINB1   : in    std_logic := 'U';
          DINB0   : in    std_logic := 'U';
          WIDTHA0 : in    std_logic := 'U';
          WIDTHA1 : in    std_logic := 'U';
          WIDTHB0 : in    std_logic := 'U';
          WIDTHB1 : in    std_logic := 'U';
          PIPEA   : in    std_logic := 'U';
          PIPEB   : in    std_logic := 'U';
          WMODEA  : in    std_logic := 'U';
          WMODEB  : in    std_logic := 'U';
          BLKA    : in    std_logic := 'U';
          BLKB    : in    std_logic := 'U';
          WENA    : in    std_logic := 'U';
          WENB    : in    std_logic := 'U';
          CLKA    : in    std_logic := 'U';
          CLKB    : in    std_logic := 'U';
          RESET   : in    std_logic := 'U';
          DOUTA8  : out   std_logic;
          DOUTA7  : out   std_logic;
          DOUTA6  : out   std_logic;
          DOUTA5  : out   std_logic;
          DOUTA4  : out   std_logic;
          DOUTA3  : out   std_logic;
          DOUTA2  : out   std_logic;
          DOUTA1  : out   std_logic;
          DOUTA0  : out   std_logic;
          DOUTB8  : out   std_logic;
          DOUTB7  : out   std_logic;
          DOUTB6  : out   std_logic;
          DOUTB5  : out   std_logic;
          DOUTB4  : out   std_logic;
          DOUTB3  : out   std_logic;
          DOUTB2  : out   std_logic;
          DOUTB1  : out   std_logic;
          DOUTB0  : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \DOUTA_1[8]\, \DOUTB_1[8]\, DPRT_512X9_SRAM_13_GND, 
        DPRT_512X9_SRAM_13_VCC : std_logic;

begin 


    DPRT_512X9_SRAM_R0C0 : RAM4K9
      generic map(MEMORYFILE => "DPRT_512X9_SRAM_R0C0.mem")

      port map(ADDRA11 => DPRT_512X9_SRAM_13_GND, ADDRA10 => 
        DPRT_512X9_SRAM_13_GND, ADDRA9 => DPRT_512X9_SRAM_13_GND, 
        ADDRA8 => DPRT_512X9_SRAM_13_GND, ADDRA7 => 
        ELINK_ADDRA_13(7), ADDRA6 => ELINK_ADDRA_13(6), ADDRA5
         => ELINK_ADDRA_13(5), ADDRA4 => ELINK_ADDRA_13(4), 
        ADDRA3 => ELINK_ADDRA_13(3), ADDRA2 => ELINK_ADDRA_13(2), 
        ADDRA1 => ELINK_ADDRA_13(1), ADDRA0 => ELINK_ADDRA_13(0), 
        ADDRB11 => DPRT_512X9_SRAM_13_GND, ADDRB10 => 
        DPRT_512X9_SRAM_13_GND, ADDRB9 => DPRT_512X9_SRAM_13_GND, 
        ADDRB8 => DPRT_512X9_SRAM_13_GND, ADDRB7 => ELKS_ADDRB_7, 
        ADDRB6 => ELKS_ADDRB_0_4, ADDRB5 => ELKS_ADDRB_5, ADDRB4
         => ELKS_ADDRB_0_2, ADDRB3 => ELKS_ADDRB_3, ADDRB2 => 
        ELKS_ADDRB_0_0, ADDRB1 => ELKS_ADDRB_1, ADDRB0 => 
        ELKS_ADDRB_0_d0, DINA8 => DPRT_512X9_SRAM_13_GND, DINA7
         => ELINK_DINA_13(7), DINA6 => ELINK_DINA_13(6), DINA5
         => ELINK_DINA_13(5), DINA4 => ELINK_DINA_13(4), DINA3
         => ELINK_DINA_13(3), DINA2 => ELINK_DINA_13(2), DINA1
         => ELINK_DINA_13(1), DINA0 => ELINK_DINA_13(0), DINB8
         => DPRT_512X9_SRAM_13_GND, DINB7 => 
        ELK_RX_SER_WORD_13(7), DINB6 => ELK_RX_SER_WORD_13(6), 
        DINB5 => ELK_RX_SER_WORD_13(5), DINB4 => 
        ELK_RX_SER_WORD_13(4), DINB3 => ELK_RX_SER_WORD_13(3), 
        DINB2 => ELK_RX_SER_WORD_13(2), DINB1 => 
        ELK_RX_SER_WORD_13(1), DINB0 => ELK_RX_SER_WORD_13(0), 
        WIDTHA0 => DPRT_512X9_SRAM_13_VCC, WIDTHA1 => 
        DPRT_512X9_SRAM_13_VCC, WIDTHB0 => DPRT_512X9_SRAM_13_VCC, 
        WIDTHB1 => DPRT_512X9_SRAM_13_VCC, PIPEA => 
        DPRT_512X9_SRAM_13_VCC, PIPEB => DPRT_512X9_SRAM_13_VCC, 
        WMODEA => DPRT_512X9_SRAM_13_GND, WMODEB => 
        DPRT_512X9_SRAM_13_GND, BLKA => ELINK_BLKA_0, BLKB => 
        ELKS_RAM_BLKB_EN, WENA => ELINK_RWA_0, WENB => ELKS_RWB, 
        CLKA => CLK60MHZ, CLKB => CLK_40M_GL, RESET => 
        P_USB_MASTER_EN_c_0, DOUTA8 => \DOUTA_1[8]\, DOUTA7 => 
        ELINK_DOUTA_13(7), DOUTA6 => ELINK_DOUTA_13(6), DOUTA5
         => ELINK_DOUTA_13(5), DOUTA4 => ELINK_DOUTA_13(4), 
        DOUTA3 => ELINK_DOUTA_13(3), DOUTA2 => ELINK_DOUTA_13(2), 
        DOUTA1 => ELINK_DOUTA_13(1), DOUTA0 => ELINK_DOUTA_13(0), 
        DOUTB8 => \DOUTB_1[8]\, DOUTB7 => PATT_ELK_DAT_13(7), 
        DOUTB6 => PATT_ELK_DAT_13(6), DOUTB5 => 
        PATT_ELK_DAT_13(5), DOUTB4 => PATT_ELK_DAT_13(4), DOUTB3
         => PATT_ELK_DAT_13(3), DOUTB2 => PATT_ELK_DAT_13(2), 
        DOUTB1 => PATT_ELK_DAT_13(1), DOUTB0 => 
        PATT_ELK_DAT_13(0));
    
    VCC_i : VCC
      port map(Y => DPRT_512X9_SRAM_13_VCC);
    
    GND_i : GND
      port map(Y => DPRT_512X9_SRAM_13_GND);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity DPRT_512X9_SRAM_12 is

    port( ELINK_RWA_0         : in    std_logic;
          ELK_RX_SER_WORD_12  : in    std_logic_vector(7 downto 0);
          ELINK_DINA_12       : in    std_logic_vector(7 downto 0);
          ELINK_BLKA_0        : in    std_logic;
          ELKS_ADDRB_0_d0     : in    std_logic;
          ELKS_ADDRB_1        : in    std_logic;
          ELKS_ADDRB_3        : in    std_logic;
          ELKS_ADDRB_5        : in    std_logic;
          ELKS_ADDRB_7        : in    std_logic;
          ELKS_ADDRB_0_0      : in    std_logic;
          ELKS_ADDRB_0_2      : in    std_logic;
          ELKS_ADDRB_0_4      : in    std_logic;
          ELINK_ADDRA_12      : in    std_logic_vector(7 downto 0);
          PATT_ELK_DAT_12     : out   std_logic_vector(7 downto 0);
          ELINK_DOUTA_12      : out   std_logic_vector(7 downto 0);
          ELKS_RWB            : in    std_logic;
          P_USB_MASTER_EN_c_0 : in    std_logic;
          CLK_40M_GL          : in    std_logic;
          CLK60MHZ            : in    std_logic;
          ELKS_RAM_BLKB_EN    : in    std_logic
        );

end DPRT_512X9_SRAM_12;

architecture DEF_ARCH of DPRT_512X9_SRAM_12 is 

  component RAM4K9
    generic (MEMORYFILE:string := "");

    port( ADDRA11 : in    std_logic := 'U';
          ADDRA10 : in    std_logic := 'U';
          ADDRA9  : in    std_logic := 'U';
          ADDRA8  : in    std_logic := 'U';
          ADDRA7  : in    std_logic := 'U';
          ADDRA6  : in    std_logic := 'U';
          ADDRA5  : in    std_logic := 'U';
          ADDRA4  : in    std_logic := 'U';
          ADDRA3  : in    std_logic := 'U';
          ADDRA2  : in    std_logic := 'U';
          ADDRA1  : in    std_logic := 'U';
          ADDRA0  : in    std_logic := 'U';
          ADDRB11 : in    std_logic := 'U';
          ADDRB10 : in    std_logic := 'U';
          ADDRB9  : in    std_logic := 'U';
          ADDRB8  : in    std_logic := 'U';
          ADDRB7  : in    std_logic := 'U';
          ADDRB6  : in    std_logic := 'U';
          ADDRB5  : in    std_logic := 'U';
          ADDRB4  : in    std_logic := 'U';
          ADDRB3  : in    std_logic := 'U';
          ADDRB2  : in    std_logic := 'U';
          ADDRB1  : in    std_logic := 'U';
          ADDRB0  : in    std_logic := 'U';
          DINA8   : in    std_logic := 'U';
          DINA7   : in    std_logic := 'U';
          DINA6   : in    std_logic := 'U';
          DINA5   : in    std_logic := 'U';
          DINA4   : in    std_logic := 'U';
          DINA3   : in    std_logic := 'U';
          DINA2   : in    std_logic := 'U';
          DINA1   : in    std_logic := 'U';
          DINA0   : in    std_logic := 'U';
          DINB8   : in    std_logic := 'U';
          DINB7   : in    std_logic := 'U';
          DINB6   : in    std_logic := 'U';
          DINB5   : in    std_logic := 'U';
          DINB4   : in    std_logic := 'U';
          DINB3   : in    std_logic := 'U';
          DINB2   : in    std_logic := 'U';
          DINB1   : in    std_logic := 'U';
          DINB0   : in    std_logic := 'U';
          WIDTHA0 : in    std_logic := 'U';
          WIDTHA1 : in    std_logic := 'U';
          WIDTHB0 : in    std_logic := 'U';
          WIDTHB1 : in    std_logic := 'U';
          PIPEA   : in    std_logic := 'U';
          PIPEB   : in    std_logic := 'U';
          WMODEA  : in    std_logic := 'U';
          WMODEB  : in    std_logic := 'U';
          BLKA    : in    std_logic := 'U';
          BLKB    : in    std_logic := 'U';
          WENA    : in    std_logic := 'U';
          WENB    : in    std_logic := 'U';
          CLKA    : in    std_logic := 'U';
          CLKB    : in    std_logic := 'U';
          RESET   : in    std_logic := 'U';
          DOUTA8  : out   std_logic;
          DOUTA7  : out   std_logic;
          DOUTA6  : out   std_logic;
          DOUTA5  : out   std_logic;
          DOUTA4  : out   std_logic;
          DOUTA3  : out   std_logic;
          DOUTA2  : out   std_logic;
          DOUTA1  : out   std_logic;
          DOUTA0  : out   std_logic;
          DOUTB8  : out   std_logic;
          DOUTB7  : out   std_logic;
          DOUTB6  : out   std_logic;
          DOUTB5  : out   std_logic;
          DOUTB4  : out   std_logic;
          DOUTB3  : out   std_logic;
          DOUTB2  : out   std_logic;
          DOUTB1  : out   std_logic;
          DOUTB0  : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \DOUTA_1[8]\, \DOUTB_1[8]\, DPRT_512X9_SRAM_12_GND, 
        DPRT_512X9_SRAM_12_VCC : std_logic;

begin 


    DPRT_512X9_SRAM_R0C0 : RAM4K9
      generic map(MEMORYFILE => "DPRT_512X9_SRAM_R0C0.mem")

      port map(ADDRA11 => DPRT_512X9_SRAM_12_GND, ADDRA10 => 
        DPRT_512X9_SRAM_12_GND, ADDRA9 => DPRT_512X9_SRAM_12_GND, 
        ADDRA8 => DPRT_512X9_SRAM_12_GND, ADDRA7 => 
        ELINK_ADDRA_12(7), ADDRA6 => ELINK_ADDRA_12(6), ADDRA5
         => ELINK_ADDRA_12(5), ADDRA4 => ELINK_ADDRA_12(4), 
        ADDRA3 => ELINK_ADDRA_12(3), ADDRA2 => ELINK_ADDRA_12(2), 
        ADDRA1 => ELINK_ADDRA_12(1), ADDRA0 => ELINK_ADDRA_12(0), 
        ADDRB11 => DPRT_512X9_SRAM_12_GND, ADDRB10 => 
        DPRT_512X9_SRAM_12_GND, ADDRB9 => DPRT_512X9_SRAM_12_GND, 
        ADDRB8 => DPRT_512X9_SRAM_12_GND, ADDRB7 => ELKS_ADDRB_7, 
        ADDRB6 => ELKS_ADDRB_0_4, ADDRB5 => ELKS_ADDRB_5, ADDRB4
         => ELKS_ADDRB_0_2, ADDRB3 => ELKS_ADDRB_3, ADDRB2 => 
        ELKS_ADDRB_0_0, ADDRB1 => ELKS_ADDRB_1, ADDRB0 => 
        ELKS_ADDRB_0_d0, DINA8 => DPRT_512X9_SRAM_12_GND, DINA7
         => ELINK_DINA_12(7), DINA6 => ELINK_DINA_12(6), DINA5
         => ELINK_DINA_12(5), DINA4 => ELINK_DINA_12(4), DINA3
         => ELINK_DINA_12(3), DINA2 => ELINK_DINA_12(2), DINA1
         => ELINK_DINA_12(1), DINA0 => ELINK_DINA_12(0), DINB8
         => DPRT_512X9_SRAM_12_GND, DINB7 => 
        ELK_RX_SER_WORD_12(7), DINB6 => ELK_RX_SER_WORD_12(6), 
        DINB5 => ELK_RX_SER_WORD_12(5), DINB4 => 
        ELK_RX_SER_WORD_12(4), DINB3 => ELK_RX_SER_WORD_12(3), 
        DINB2 => ELK_RX_SER_WORD_12(2), DINB1 => 
        ELK_RX_SER_WORD_12(1), DINB0 => ELK_RX_SER_WORD_12(0), 
        WIDTHA0 => DPRT_512X9_SRAM_12_VCC, WIDTHA1 => 
        DPRT_512X9_SRAM_12_VCC, WIDTHB0 => DPRT_512X9_SRAM_12_VCC, 
        WIDTHB1 => DPRT_512X9_SRAM_12_VCC, PIPEA => 
        DPRT_512X9_SRAM_12_VCC, PIPEB => DPRT_512X9_SRAM_12_VCC, 
        WMODEA => DPRT_512X9_SRAM_12_GND, WMODEB => 
        DPRT_512X9_SRAM_12_GND, BLKA => ELINK_BLKA_0, BLKB => 
        ELKS_RAM_BLKB_EN, WENA => ELINK_RWA_0, WENB => ELKS_RWB, 
        CLKA => CLK60MHZ, CLKB => CLK_40M_GL, RESET => 
        P_USB_MASTER_EN_c_0, DOUTA8 => \DOUTA_1[8]\, DOUTA7 => 
        ELINK_DOUTA_12(7), DOUTA6 => ELINK_DOUTA_12(6), DOUTA5
         => ELINK_DOUTA_12(5), DOUTA4 => ELINK_DOUTA_12(4), 
        DOUTA3 => ELINK_DOUTA_12(3), DOUTA2 => ELINK_DOUTA_12(2), 
        DOUTA1 => ELINK_DOUTA_12(1), DOUTA0 => ELINK_DOUTA_12(0), 
        DOUTB8 => \DOUTB_1[8]\, DOUTB7 => PATT_ELK_DAT_12(7), 
        DOUTB6 => PATT_ELK_DAT_12(6), DOUTB5 => 
        PATT_ELK_DAT_12(5), DOUTB4 => PATT_ELK_DAT_12(4), DOUTB3
         => PATT_ELK_DAT_12(3), DOUTB2 => PATT_ELK_DAT_12(2), 
        DOUTB1 => PATT_ELK_DAT_12(1), DOUTB0 => 
        PATT_ELK_DAT_12(0));
    
    VCC_i : VCC
      port map(Y => DPRT_512X9_SRAM_12_VCC);
    
    GND_i : GND
      port map(Y => DPRT_512X9_SRAM_12_GND);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity DPRT_512X9_SRAM_11 is

    port( ELINK_RWA_0         : in    std_logic;
          ELK_RX_SER_WORD_11  : in    std_logic_vector(7 downto 0);
          ELINK_DINA_11       : in    std_logic_vector(7 downto 0);
          ELINK_BLKA_0        : in    std_logic;
          ELKS_ADDRB_0_d0     : in    std_logic;
          ELKS_ADDRB_1        : in    std_logic;
          ELKS_ADDRB_3        : in    std_logic;
          ELKS_ADDRB_5        : in    std_logic;
          ELKS_ADDRB_7        : in    std_logic;
          ELKS_ADDRB_0_0      : in    std_logic;
          ELKS_ADDRB_0_2      : in    std_logic;
          ELKS_ADDRB_0_4      : in    std_logic;
          ELINK_ADDRA_11      : in    std_logic_vector(7 downto 0);
          PATT_ELK_DAT_11     : out   std_logic_vector(7 downto 0);
          ELINK_DOUTA_11      : out   std_logic_vector(7 downto 0);
          ELKS_RWB            : in    std_logic;
          P_USB_MASTER_EN_c_0 : in    std_logic;
          CLK_40M_GL          : in    std_logic;
          CLK60MHZ            : in    std_logic;
          ELKS_RAM_BLKB_EN    : in    std_logic
        );

end DPRT_512X9_SRAM_11;

architecture DEF_ARCH of DPRT_512X9_SRAM_11 is 

  component RAM4K9
    generic (MEMORYFILE:string := "");

    port( ADDRA11 : in    std_logic := 'U';
          ADDRA10 : in    std_logic := 'U';
          ADDRA9  : in    std_logic := 'U';
          ADDRA8  : in    std_logic := 'U';
          ADDRA7  : in    std_logic := 'U';
          ADDRA6  : in    std_logic := 'U';
          ADDRA5  : in    std_logic := 'U';
          ADDRA4  : in    std_logic := 'U';
          ADDRA3  : in    std_logic := 'U';
          ADDRA2  : in    std_logic := 'U';
          ADDRA1  : in    std_logic := 'U';
          ADDRA0  : in    std_logic := 'U';
          ADDRB11 : in    std_logic := 'U';
          ADDRB10 : in    std_logic := 'U';
          ADDRB9  : in    std_logic := 'U';
          ADDRB8  : in    std_logic := 'U';
          ADDRB7  : in    std_logic := 'U';
          ADDRB6  : in    std_logic := 'U';
          ADDRB5  : in    std_logic := 'U';
          ADDRB4  : in    std_logic := 'U';
          ADDRB3  : in    std_logic := 'U';
          ADDRB2  : in    std_logic := 'U';
          ADDRB1  : in    std_logic := 'U';
          ADDRB0  : in    std_logic := 'U';
          DINA8   : in    std_logic := 'U';
          DINA7   : in    std_logic := 'U';
          DINA6   : in    std_logic := 'U';
          DINA5   : in    std_logic := 'U';
          DINA4   : in    std_logic := 'U';
          DINA3   : in    std_logic := 'U';
          DINA2   : in    std_logic := 'U';
          DINA1   : in    std_logic := 'U';
          DINA0   : in    std_logic := 'U';
          DINB8   : in    std_logic := 'U';
          DINB7   : in    std_logic := 'U';
          DINB6   : in    std_logic := 'U';
          DINB5   : in    std_logic := 'U';
          DINB4   : in    std_logic := 'U';
          DINB3   : in    std_logic := 'U';
          DINB2   : in    std_logic := 'U';
          DINB1   : in    std_logic := 'U';
          DINB0   : in    std_logic := 'U';
          WIDTHA0 : in    std_logic := 'U';
          WIDTHA1 : in    std_logic := 'U';
          WIDTHB0 : in    std_logic := 'U';
          WIDTHB1 : in    std_logic := 'U';
          PIPEA   : in    std_logic := 'U';
          PIPEB   : in    std_logic := 'U';
          WMODEA  : in    std_logic := 'U';
          WMODEB  : in    std_logic := 'U';
          BLKA    : in    std_logic := 'U';
          BLKB    : in    std_logic := 'U';
          WENA    : in    std_logic := 'U';
          WENB    : in    std_logic := 'U';
          CLKA    : in    std_logic := 'U';
          CLKB    : in    std_logic := 'U';
          RESET   : in    std_logic := 'U';
          DOUTA8  : out   std_logic;
          DOUTA7  : out   std_logic;
          DOUTA6  : out   std_logic;
          DOUTA5  : out   std_logic;
          DOUTA4  : out   std_logic;
          DOUTA3  : out   std_logic;
          DOUTA2  : out   std_logic;
          DOUTA1  : out   std_logic;
          DOUTA0  : out   std_logic;
          DOUTB8  : out   std_logic;
          DOUTB7  : out   std_logic;
          DOUTB6  : out   std_logic;
          DOUTB5  : out   std_logic;
          DOUTB4  : out   std_logic;
          DOUTB3  : out   std_logic;
          DOUTB2  : out   std_logic;
          DOUTB1  : out   std_logic;
          DOUTB0  : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \DOUTA_1[8]\, \DOUTB_1[8]\, DPRT_512X9_SRAM_11_GND, 
        DPRT_512X9_SRAM_11_VCC : std_logic;

begin 


    DPRT_512X9_SRAM_R0C0 : RAM4K9
      generic map(MEMORYFILE => "DPRT_512X9_SRAM_R0C0.mem")

      port map(ADDRA11 => DPRT_512X9_SRAM_11_GND, ADDRA10 => 
        DPRT_512X9_SRAM_11_GND, ADDRA9 => DPRT_512X9_SRAM_11_GND, 
        ADDRA8 => DPRT_512X9_SRAM_11_GND, ADDRA7 => 
        ELINK_ADDRA_11(7), ADDRA6 => ELINK_ADDRA_11(6), ADDRA5
         => ELINK_ADDRA_11(5), ADDRA4 => ELINK_ADDRA_11(4), 
        ADDRA3 => ELINK_ADDRA_11(3), ADDRA2 => ELINK_ADDRA_11(2), 
        ADDRA1 => ELINK_ADDRA_11(1), ADDRA0 => ELINK_ADDRA_11(0), 
        ADDRB11 => DPRT_512X9_SRAM_11_GND, ADDRB10 => 
        DPRT_512X9_SRAM_11_GND, ADDRB9 => DPRT_512X9_SRAM_11_GND, 
        ADDRB8 => DPRT_512X9_SRAM_11_GND, ADDRB7 => ELKS_ADDRB_7, 
        ADDRB6 => ELKS_ADDRB_0_4, ADDRB5 => ELKS_ADDRB_5, ADDRB4
         => ELKS_ADDRB_0_2, ADDRB3 => ELKS_ADDRB_3, ADDRB2 => 
        ELKS_ADDRB_0_0, ADDRB1 => ELKS_ADDRB_1, ADDRB0 => 
        ELKS_ADDRB_0_d0, DINA8 => DPRT_512X9_SRAM_11_GND, DINA7
         => ELINK_DINA_11(7), DINA6 => ELINK_DINA_11(6), DINA5
         => ELINK_DINA_11(5), DINA4 => ELINK_DINA_11(4), DINA3
         => ELINK_DINA_11(3), DINA2 => ELINK_DINA_11(2), DINA1
         => ELINK_DINA_11(1), DINA0 => ELINK_DINA_11(0), DINB8
         => DPRT_512X9_SRAM_11_GND, DINB7 => 
        ELK_RX_SER_WORD_11(7), DINB6 => ELK_RX_SER_WORD_11(6), 
        DINB5 => ELK_RX_SER_WORD_11(5), DINB4 => 
        ELK_RX_SER_WORD_11(4), DINB3 => ELK_RX_SER_WORD_11(3), 
        DINB2 => ELK_RX_SER_WORD_11(2), DINB1 => 
        ELK_RX_SER_WORD_11(1), DINB0 => ELK_RX_SER_WORD_11(0), 
        WIDTHA0 => DPRT_512X9_SRAM_11_VCC, WIDTHA1 => 
        DPRT_512X9_SRAM_11_VCC, WIDTHB0 => DPRT_512X9_SRAM_11_VCC, 
        WIDTHB1 => DPRT_512X9_SRAM_11_VCC, PIPEA => 
        DPRT_512X9_SRAM_11_VCC, PIPEB => DPRT_512X9_SRAM_11_VCC, 
        WMODEA => DPRT_512X9_SRAM_11_GND, WMODEB => 
        DPRT_512X9_SRAM_11_GND, BLKA => ELINK_BLKA_0, BLKB => 
        ELKS_RAM_BLKB_EN, WENA => ELINK_RWA_0, WENB => ELKS_RWB, 
        CLKA => CLK60MHZ, CLKB => CLK_40M_GL, RESET => 
        P_USB_MASTER_EN_c_0, DOUTA8 => \DOUTA_1[8]\, DOUTA7 => 
        ELINK_DOUTA_11(7), DOUTA6 => ELINK_DOUTA_11(6), DOUTA5
         => ELINK_DOUTA_11(5), DOUTA4 => ELINK_DOUTA_11(4), 
        DOUTA3 => ELINK_DOUTA_11(3), DOUTA2 => ELINK_DOUTA_11(2), 
        DOUTA1 => ELINK_DOUTA_11(1), DOUTA0 => ELINK_DOUTA_11(0), 
        DOUTB8 => \DOUTB_1[8]\, DOUTB7 => PATT_ELK_DAT_11(7), 
        DOUTB6 => PATT_ELK_DAT_11(6), DOUTB5 => 
        PATT_ELK_DAT_11(5), DOUTB4 => PATT_ELK_DAT_11(4), DOUTB3
         => PATT_ELK_DAT_11(3), DOUTB2 => PATT_ELK_DAT_11(2), 
        DOUTB1 => PATT_ELK_DAT_11(1), DOUTB0 => 
        PATT_ELK_DAT_11(0));
    
    VCC_i : VCC
      port map(Y => DPRT_512X9_SRAM_11_VCC);
    
    GND_i : GND
      port map(Y => DPRT_512X9_SRAM_11_GND);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity DPRT_512X9_SRAM_16 is

    port( ELINK_RWA_0         : in    std_logic;
          ELK_RX_SER_WORD_16  : in    std_logic_vector(7 downto 0);
          ELINK_DINA_16       : in    std_logic_vector(7 downto 0);
          ELINK_BLKA_0        : in    std_logic;
          ELKS_ADDRB_0_d0     : in    std_logic;
          ELKS_ADDRB_1        : in    std_logic;
          ELKS_ADDRB_3        : in    std_logic;
          ELKS_ADDRB_5        : in    std_logic;
          ELKS_ADDRB_7        : in    std_logic;
          ELKS_ADDRB_0_0      : in    std_logic;
          ELKS_ADDRB_0_2      : in    std_logic;
          ELKS_ADDRB_0_4      : in    std_logic;
          ELINK_ADDRA_16      : in    std_logic_vector(7 downto 0);
          PATT_ELK_DAT_16     : out   std_logic_vector(7 downto 0);
          ELINK_DOUTA_16      : out   std_logic_vector(7 downto 0);
          ELKS_RWB            : in    std_logic;
          P_USB_MASTER_EN_c_0 : in    std_logic;
          CLK_40M_GL          : in    std_logic;
          CLK60MHZ            : in    std_logic;
          ELKS_RAM_BLKB_EN    : in    std_logic
        );

end DPRT_512X9_SRAM_16;

architecture DEF_ARCH of DPRT_512X9_SRAM_16 is 

  component RAM4K9
    generic (MEMORYFILE:string := "");

    port( ADDRA11 : in    std_logic := 'U';
          ADDRA10 : in    std_logic := 'U';
          ADDRA9  : in    std_logic := 'U';
          ADDRA8  : in    std_logic := 'U';
          ADDRA7  : in    std_logic := 'U';
          ADDRA6  : in    std_logic := 'U';
          ADDRA5  : in    std_logic := 'U';
          ADDRA4  : in    std_logic := 'U';
          ADDRA3  : in    std_logic := 'U';
          ADDRA2  : in    std_logic := 'U';
          ADDRA1  : in    std_logic := 'U';
          ADDRA0  : in    std_logic := 'U';
          ADDRB11 : in    std_logic := 'U';
          ADDRB10 : in    std_logic := 'U';
          ADDRB9  : in    std_logic := 'U';
          ADDRB8  : in    std_logic := 'U';
          ADDRB7  : in    std_logic := 'U';
          ADDRB6  : in    std_logic := 'U';
          ADDRB5  : in    std_logic := 'U';
          ADDRB4  : in    std_logic := 'U';
          ADDRB3  : in    std_logic := 'U';
          ADDRB2  : in    std_logic := 'U';
          ADDRB1  : in    std_logic := 'U';
          ADDRB0  : in    std_logic := 'U';
          DINA8   : in    std_logic := 'U';
          DINA7   : in    std_logic := 'U';
          DINA6   : in    std_logic := 'U';
          DINA5   : in    std_logic := 'U';
          DINA4   : in    std_logic := 'U';
          DINA3   : in    std_logic := 'U';
          DINA2   : in    std_logic := 'U';
          DINA1   : in    std_logic := 'U';
          DINA0   : in    std_logic := 'U';
          DINB8   : in    std_logic := 'U';
          DINB7   : in    std_logic := 'U';
          DINB6   : in    std_logic := 'U';
          DINB5   : in    std_logic := 'U';
          DINB4   : in    std_logic := 'U';
          DINB3   : in    std_logic := 'U';
          DINB2   : in    std_logic := 'U';
          DINB1   : in    std_logic := 'U';
          DINB0   : in    std_logic := 'U';
          WIDTHA0 : in    std_logic := 'U';
          WIDTHA1 : in    std_logic := 'U';
          WIDTHB0 : in    std_logic := 'U';
          WIDTHB1 : in    std_logic := 'U';
          PIPEA   : in    std_logic := 'U';
          PIPEB   : in    std_logic := 'U';
          WMODEA  : in    std_logic := 'U';
          WMODEB  : in    std_logic := 'U';
          BLKA    : in    std_logic := 'U';
          BLKB    : in    std_logic := 'U';
          WENA    : in    std_logic := 'U';
          WENB    : in    std_logic := 'U';
          CLKA    : in    std_logic := 'U';
          CLKB    : in    std_logic := 'U';
          RESET   : in    std_logic := 'U';
          DOUTA8  : out   std_logic;
          DOUTA7  : out   std_logic;
          DOUTA6  : out   std_logic;
          DOUTA5  : out   std_logic;
          DOUTA4  : out   std_logic;
          DOUTA3  : out   std_logic;
          DOUTA2  : out   std_logic;
          DOUTA1  : out   std_logic;
          DOUTA0  : out   std_logic;
          DOUTB8  : out   std_logic;
          DOUTB7  : out   std_logic;
          DOUTB6  : out   std_logic;
          DOUTB5  : out   std_logic;
          DOUTB4  : out   std_logic;
          DOUTB3  : out   std_logic;
          DOUTB2  : out   std_logic;
          DOUTB1  : out   std_logic;
          DOUTB0  : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \DOUTA_1[8]\, \DOUTB_1[8]\, DPRT_512X9_SRAM_16_GND, 
        DPRT_512X9_SRAM_16_VCC : std_logic;

begin 


    DPRT_512X9_SRAM_R0C0 : RAM4K9
      generic map(MEMORYFILE => "DPRT_512X9_SRAM_R0C0.mem")

      port map(ADDRA11 => DPRT_512X9_SRAM_16_GND, ADDRA10 => 
        DPRT_512X9_SRAM_16_GND, ADDRA9 => DPRT_512X9_SRAM_16_GND, 
        ADDRA8 => DPRT_512X9_SRAM_16_GND, ADDRA7 => 
        ELINK_ADDRA_16(7), ADDRA6 => ELINK_ADDRA_16(6), ADDRA5
         => ELINK_ADDRA_16(5), ADDRA4 => ELINK_ADDRA_16(4), 
        ADDRA3 => ELINK_ADDRA_16(3), ADDRA2 => ELINK_ADDRA_16(2), 
        ADDRA1 => ELINK_ADDRA_16(1), ADDRA0 => ELINK_ADDRA_16(0), 
        ADDRB11 => DPRT_512X9_SRAM_16_GND, ADDRB10 => 
        DPRT_512X9_SRAM_16_GND, ADDRB9 => DPRT_512X9_SRAM_16_GND, 
        ADDRB8 => DPRT_512X9_SRAM_16_GND, ADDRB7 => ELKS_ADDRB_7, 
        ADDRB6 => ELKS_ADDRB_0_4, ADDRB5 => ELKS_ADDRB_5, ADDRB4
         => ELKS_ADDRB_0_2, ADDRB3 => ELKS_ADDRB_3, ADDRB2 => 
        ELKS_ADDRB_0_0, ADDRB1 => ELKS_ADDRB_1, ADDRB0 => 
        ELKS_ADDRB_0_d0, DINA8 => DPRT_512X9_SRAM_16_GND, DINA7
         => ELINK_DINA_16(7), DINA6 => ELINK_DINA_16(6), DINA5
         => ELINK_DINA_16(5), DINA4 => ELINK_DINA_16(4), DINA3
         => ELINK_DINA_16(3), DINA2 => ELINK_DINA_16(2), DINA1
         => ELINK_DINA_16(1), DINA0 => ELINK_DINA_16(0), DINB8
         => DPRT_512X9_SRAM_16_GND, DINB7 => 
        ELK_RX_SER_WORD_16(7), DINB6 => ELK_RX_SER_WORD_16(6), 
        DINB5 => ELK_RX_SER_WORD_16(5), DINB4 => 
        ELK_RX_SER_WORD_16(4), DINB3 => ELK_RX_SER_WORD_16(3), 
        DINB2 => ELK_RX_SER_WORD_16(2), DINB1 => 
        ELK_RX_SER_WORD_16(1), DINB0 => ELK_RX_SER_WORD_16(0), 
        WIDTHA0 => DPRT_512X9_SRAM_16_VCC, WIDTHA1 => 
        DPRT_512X9_SRAM_16_VCC, WIDTHB0 => DPRT_512X9_SRAM_16_VCC, 
        WIDTHB1 => DPRT_512X9_SRAM_16_VCC, PIPEA => 
        DPRT_512X9_SRAM_16_VCC, PIPEB => DPRT_512X9_SRAM_16_VCC, 
        WMODEA => DPRT_512X9_SRAM_16_GND, WMODEB => 
        DPRT_512X9_SRAM_16_GND, BLKA => ELINK_BLKA_0, BLKB => 
        ELKS_RAM_BLKB_EN, WENA => ELINK_RWA_0, WENB => ELKS_RWB, 
        CLKA => CLK60MHZ, CLKB => CLK_40M_GL, RESET => 
        P_USB_MASTER_EN_c_0, DOUTA8 => \DOUTA_1[8]\, DOUTA7 => 
        ELINK_DOUTA_16(7), DOUTA6 => ELINK_DOUTA_16(6), DOUTA5
         => ELINK_DOUTA_16(5), DOUTA4 => ELINK_DOUTA_16(4), 
        DOUTA3 => ELINK_DOUTA_16(3), DOUTA2 => ELINK_DOUTA_16(2), 
        DOUTA1 => ELINK_DOUTA_16(1), DOUTA0 => ELINK_DOUTA_16(0), 
        DOUTB8 => \DOUTB_1[8]\, DOUTB7 => PATT_ELK_DAT_16(7), 
        DOUTB6 => PATT_ELK_DAT_16(6), DOUTB5 => 
        PATT_ELK_DAT_16(5), DOUTB4 => PATT_ELK_DAT_16(4), DOUTB3
         => PATT_ELK_DAT_16(3), DOUTB2 => PATT_ELK_DAT_16(2), 
        DOUTB1 => PATT_ELK_DAT_16(1), DOUTB0 => 
        PATT_ELK_DAT_16(0));
    
    VCC_i : VCC
      port map(Y => DPRT_512X9_SRAM_16_VCC);
    
    GND_i : GND
      port map(Y => DPRT_512X9_SRAM_16_GND);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity CLK60M_TO_40M_4_1 is

    port( ELINKS_STRT_ADDR      : in    std_logic_vector(7 downto 0);
          ELKS_STRT_ADDR        : out   std_logic_vector(7 downto 0);
          P_MASTER_POR_B_c_28   : in    std_logic;
          P_MASTER_POR_B_c_22_0 : in    std_logic;
          P_MASTER_POR_B_c_33   : in    std_logic;
          P_MASTER_POR_B_c_21   : in    std_logic;
          P_MASTER_POR_B_c_32   : in    std_logic;
          CLK_40M_GL            : in    std_logic
        );

end CLK60M_TO_40M_4_1;

architecture DEF_ARCH of CLK60M_TO_40M_4_1 is 

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component XO1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component MX2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal un1_SAMP_TWO_NE_4, un1_SAMP_TWO_5, un1_SAMP_TWO_4, 
        un1_SAMP_TWO_NE_1, un1_SAMP_TWO_NE_3, \ELKS_STRT_ADDR[2]\, 
        \SAMP_TWO[2]_net_1\, un1_SAMP_TWO_3, un1_SAMP_TWO_NE_2, 
        \ELKS_STRT_ADDR[0]\, \SAMP_TWO[0]_net_1\, un1_SAMP_TWO_1, 
        \ELKS_STRT_ADDR[6]\, \SAMP_TWO[6]_net_1\, un1_SAMP_TWO_7, 
        n_sync_sm3, \N_DELCNT[0]\, \SYNC_SM[0]_net_1\, 
        \DELCNT[0]_net_1\, un7_delcnt, \DELCNT[1]_net_1\, 
        \N_SYNC_SM[0]\, \SAMP_TWO[7]_net_1\, \ELKS_STRT_ADDR[7]\, 
        \SAMP_TWO[5]_net_1\, \ELKS_STRT_ADDR[5]\, 
        \SAMP_TWO[4]_net_1\, \ELKS_STRT_ADDR[4]\, 
        \SAMP_TWO[3]_net_1\, \ELKS_STRT_ADDR[3]\, 
        \SAMP_TWO[1]_net_1\, \ELKS_STRT_ADDR[1]\, SUM1_2, 
        \SAMP_ONE[0]_net_1\, \SAMP_ONE[1]_net_1\, 
        \SAMP_ONE[2]_net_1\, \SAMP_ONE[3]_net_1\, 
        \SAMP_ONE[4]_net_1\, \SAMP_ONE[5]_net_1\, 
        \SAMP_ONE[6]_net_1\, \SAMP_ONE[7]_net_1\, \GND\, \VCC\
         : std_logic;

begin 

    ELKS_STRT_ADDR(7) <= \ELKS_STRT_ADDR[7]\;
    ELKS_STRT_ADDR(6) <= \ELKS_STRT_ADDR[6]\;
    ELKS_STRT_ADDR(5) <= \ELKS_STRT_ADDR[5]\;
    ELKS_STRT_ADDR(4) <= \ELKS_STRT_ADDR[4]\;
    ELKS_STRT_ADDR(3) <= \ELKS_STRT_ADDR[3]\;
    ELKS_STRT_ADDR(2) <= \ELKS_STRT_ADDR[2]\;
    ELKS_STRT_ADDR(1) <= \ELKS_STRT_ADDR[1]\;
    ELKS_STRT_ADDR(0) <= \ELKS_STRT_ADDR[0]\;

    \SAMP_ONE[2]\ : DFN1C0
      port map(D => ELINKS_STRT_ADDR(2), CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_33, Q => \SAMP_ONE[2]_net_1\);
    
    \SYNC_SM_RNO_6[0]\ : XOR2
      port map(A => \SAMP_TWO[5]_net_1\, B => \ELKS_STRT_ADDR[5]\, 
        Y => un1_SAMP_TWO_5);
    
    \LOCAL_REG_VAL[3]\ : DFN1E1C0
      port map(D => \SAMP_TWO[3]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_21, E => un7_delcnt, Q => 
        \ELKS_STRT_ADDR[3]\);
    
    \SYNC_SM[0]\ : DFN1C0
      port map(D => \N_SYNC_SM[0]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_32, Q => \SYNC_SM[0]_net_1\);
    
    \SYNC_SM_RNO_5[0]\ : XOR2
      port map(A => \SAMP_TWO[1]_net_1\, B => \ELKS_STRT_ADDR[1]\, 
        Y => un1_SAMP_TWO_1);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \DELCNT[1]\ : DFN1C0
      port map(D => SUM1_2, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_28, Q => \DELCNT[1]_net_1\);
    
    \LOCAL_REG_VAL[5]\ : DFN1E1C0
      port map(D => \SAMP_TWO[5]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_21, E => un7_delcnt, Q => 
        \ELKS_STRT_ADDR[5]\);
    
    \SYNC_SM_RNO_1[0]\ : XO1
      port map(A => \ELKS_STRT_ADDR[2]\, B => \SAMP_TWO[2]_net_1\, 
        C => un1_SAMP_TWO_3, Y => un1_SAMP_TWO_NE_3);
    
    \SAMP_TWO[0]\ : DFN1C0
      port map(D => \SAMP_ONE[0]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_22_0, Q => \SAMP_TWO[0]_net_1\);
    
    \SAMP_ONE[1]\ : DFN1C0
      port map(D => ELINKS_STRT_ADDR(1), CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_33, Q => \SAMP_ONE[1]_net_1\);
    
    \SAMP_TWO[1]\ : DFN1C0
      port map(D => \SAMP_ONE[1]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_22_0, Q => \SAMP_TWO[1]_net_1\);
    
    \SYNC_SM_RNO_3[0]\ : OR3
      port map(A => un1_SAMP_TWO_5, B => un1_SAMP_TWO_4, C => 
        un1_SAMP_TWO_NE_1, Y => un1_SAMP_TWO_NE_4);
    
    \SYNC_SM_RNO_9[0]\ : XOR2
      port map(A => \SAMP_TWO[7]_net_1\, B => \ELKS_STRT_ADDR[7]\, 
        Y => un1_SAMP_TWO_7);
    
    un2_n_delcnt_1_1_SUM1 : XOR2
      port map(A => \DELCNT[1]_net_1\, B => \DELCNT[0]_net_1\, Y
         => SUM1_2);
    
    \SAMP_TWO[3]\ : DFN1C0
      port map(D => \SAMP_ONE[3]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_22_0, Q => \SAMP_TWO[3]_net_1\);
    
    \SYNC_SM_RNO_8[0]\ : XO1
      port map(A => \ELKS_STRT_ADDR[6]\, B => \SAMP_TWO[6]_net_1\, 
        C => un1_SAMP_TWO_7, Y => un1_SAMP_TWO_NE_1);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \SYNC_SM_RNO_4[0]\ : XOR2
      port map(A => \SAMP_TWO[3]_net_1\, B => \ELKS_STRT_ADDR[3]\, 
        Y => un1_SAMP_TWO_3);
    
    \SYNC_SM_RNO[0]\ : MX2B
      port map(A => n_sync_sm3, B => un7_delcnt, S => 
        \SYNC_SM[0]_net_1\, Y => \N_SYNC_SM[0]\);
    
    \SAMP_ONE[4]\ : DFN1C0
      port map(D => ELINKS_STRT_ADDR(4), CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_33, Q => \SAMP_ONE[4]_net_1\);
    
    \LOCAL_REG_VAL[2]\ : DFN1E1C0
      port map(D => \SAMP_TWO[2]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_21, E => un7_delcnt, Q => 
        \ELKS_STRT_ADDR[2]\);
    
    \SAMP_TWO[5]\ : DFN1C0
      port map(D => \SAMP_ONE[5]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_22_0, Q => \SAMP_TWO[5]_net_1\);
    
    \SAMP_TWO[4]\ : DFN1C0
      port map(D => \SAMP_ONE[4]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_22_0, Q => \SAMP_TWO[4]_net_1\);
    
    \SAMP_TWO[2]\ : DFN1C0
      port map(D => \SAMP_ONE[2]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_22_0, Q => \SAMP_TWO[2]_net_1\);
    
    \DELCNT_RNO[0]\ : NOR2A
      port map(A => \SYNC_SM[0]_net_1\, B => \DELCNT[0]_net_1\, Y
         => \N_DELCNT[0]\);
    
    \LOCAL_REG_VAL[0]\ : DFN1E1C0
      port map(D => \SAMP_TWO[0]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_21, E => un7_delcnt, Q => 
        \ELKS_STRT_ADDR[0]\);
    
    \LOCAL_REG_VAL[7]\ : DFN1E1C0
      port map(D => \SAMP_TWO[7]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_21, E => un7_delcnt, Q => 
        \ELKS_STRT_ADDR[7]\);
    
    \SYNC_SM_RNO_0[0]\ : OR3
      port map(A => un1_SAMP_TWO_NE_3, B => un1_SAMP_TWO_NE_2, C
         => un1_SAMP_TWO_NE_4, Y => n_sync_sm3);
    
    \DELCNT[0]\ : DFN1C0
      port map(D => \N_DELCNT[0]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_28, Q => \DELCNT[0]_net_1\);
    
    \LOCAL_REG_VAL[4]\ : DFN1E1C0
      port map(D => \SAMP_TWO[4]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_21, E => un7_delcnt, Q => 
        \ELKS_STRT_ADDR[4]\);
    
    \SAMP_ONE[7]\ : DFN1C0
      port map(D => ELINKS_STRT_ADDR(7), CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_33, Q => \SAMP_ONE[7]_net_1\);
    
    \SYNC_SM_RNO_2[0]\ : XO1
      port map(A => \ELKS_STRT_ADDR[0]\, B => \SAMP_TWO[0]_net_1\, 
        C => un1_SAMP_TWO_1, Y => un1_SAMP_TWO_NE_2);
    
    \SAMP_TWO[7]\ : DFN1C0
      port map(D => \SAMP_ONE[7]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_22_0, Q => \SAMP_TWO[7]_net_1\);
    
    \DELCNT_RNINMVG[1]\ : NOR2B
      port map(A => \DELCNT[1]_net_1\, B => \DELCNT[0]_net_1\, Y
         => un7_delcnt);
    
    \SAMP_ONE[5]\ : DFN1C0
      port map(D => ELINKS_STRT_ADDR(5), CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_33, Q => \SAMP_ONE[5]_net_1\);
    
    \LOCAL_REG_VAL[6]\ : DFN1E1C0
      port map(D => \SAMP_TWO[6]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_21, E => un7_delcnt, Q => 
        \ELKS_STRT_ADDR[6]\);
    
    \SYNC_SM_RNO_7[0]\ : XOR2
      port map(A => \SAMP_TWO[4]_net_1\, B => \ELKS_STRT_ADDR[4]\, 
        Y => un1_SAMP_TWO_4);
    
    \SAMP_ONE[6]\ : DFN1C0
      port map(D => ELINKS_STRT_ADDR(6), CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_33, Q => \SAMP_ONE[6]_net_1\);
    
    \SAMP_ONE[0]\ : DFN1C0
      port map(D => ELINKS_STRT_ADDR(0), CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_33, Q => \SAMP_ONE[0]_net_1\);
    
    \LOCAL_REG_VAL[1]\ : DFN1E1C0
      port map(D => \SAMP_TWO[1]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_21, E => un7_delcnt, Q => 
        \ELKS_STRT_ADDR[1]\);
    
    \SAMP_TWO[6]\ : DFN1C0
      port map(D => \SAMP_ONE[6]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_22_0, Q => \SAMP_TWO[6]_net_1\);
    
    \SAMP_ONE[3]\ : DFN1C0
      port map(D => ELINKS_STRT_ADDR(3), CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_33, Q => \SAMP_ONE[3]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity DPRT_512X9_SRAM_3 is

    port( ELINK_RWA_0         : in    std_logic;
          ELK_RX_SER_WORD_3   : in    std_logic_vector(7 downto 0);
          ELINK_DINA_3        : in    std_logic_vector(7 downto 0);
          ELINK_BLKA_0        : in    std_logic;
          ELKS_ADDRB_0_d0     : in    std_logic;
          ELKS_ADDRB_1        : in    std_logic;
          ELKS_ADDRB_3        : in    std_logic;
          ELKS_ADDRB_5        : in    std_logic;
          ELKS_ADDRB_7        : in    std_logic;
          ELKS_ADDRB_0_0      : in    std_logic;
          ELKS_ADDRB_0_2      : in    std_logic;
          ELKS_ADDRB_0_4      : in    std_logic;
          ELINK_ADDRA_3       : in    std_logic_vector(7 downto 0);
          PATT_ELK_DAT_3      : out   std_logic_vector(7 downto 0);
          ELINK_DOUTA_3       : out   std_logic_vector(7 downto 0);
          ELKS_RWB            : in    std_logic;
          P_USB_MASTER_EN_c_0 : in    std_logic;
          CLK_40M_GL          : in    std_logic;
          CLK60MHZ            : in    std_logic;
          ELKS_RAM_BLKB_EN    : in    std_logic
        );

end DPRT_512X9_SRAM_3;

architecture DEF_ARCH of DPRT_512X9_SRAM_3 is 

  component RAM4K9
    generic (MEMORYFILE:string := "");

    port( ADDRA11 : in    std_logic := 'U';
          ADDRA10 : in    std_logic := 'U';
          ADDRA9  : in    std_logic := 'U';
          ADDRA8  : in    std_logic := 'U';
          ADDRA7  : in    std_logic := 'U';
          ADDRA6  : in    std_logic := 'U';
          ADDRA5  : in    std_logic := 'U';
          ADDRA4  : in    std_logic := 'U';
          ADDRA3  : in    std_logic := 'U';
          ADDRA2  : in    std_logic := 'U';
          ADDRA1  : in    std_logic := 'U';
          ADDRA0  : in    std_logic := 'U';
          ADDRB11 : in    std_logic := 'U';
          ADDRB10 : in    std_logic := 'U';
          ADDRB9  : in    std_logic := 'U';
          ADDRB8  : in    std_logic := 'U';
          ADDRB7  : in    std_logic := 'U';
          ADDRB6  : in    std_logic := 'U';
          ADDRB5  : in    std_logic := 'U';
          ADDRB4  : in    std_logic := 'U';
          ADDRB3  : in    std_logic := 'U';
          ADDRB2  : in    std_logic := 'U';
          ADDRB1  : in    std_logic := 'U';
          ADDRB0  : in    std_logic := 'U';
          DINA8   : in    std_logic := 'U';
          DINA7   : in    std_logic := 'U';
          DINA6   : in    std_logic := 'U';
          DINA5   : in    std_logic := 'U';
          DINA4   : in    std_logic := 'U';
          DINA3   : in    std_logic := 'U';
          DINA2   : in    std_logic := 'U';
          DINA1   : in    std_logic := 'U';
          DINA0   : in    std_logic := 'U';
          DINB8   : in    std_logic := 'U';
          DINB7   : in    std_logic := 'U';
          DINB6   : in    std_logic := 'U';
          DINB5   : in    std_logic := 'U';
          DINB4   : in    std_logic := 'U';
          DINB3   : in    std_logic := 'U';
          DINB2   : in    std_logic := 'U';
          DINB1   : in    std_logic := 'U';
          DINB0   : in    std_logic := 'U';
          WIDTHA0 : in    std_logic := 'U';
          WIDTHA1 : in    std_logic := 'U';
          WIDTHB0 : in    std_logic := 'U';
          WIDTHB1 : in    std_logic := 'U';
          PIPEA   : in    std_logic := 'U';
          PIPEB   : in    std_logic := 'U';
          WMODEA  : in    std_logic := 'U';
          WMODEB  : in    std_logic := 'U';
          BLKA    : in    std_logic := 'U';
          BLKB    : in    std_logic := 'U';
          WENA    : in    std_logic := 'U';
          WENB    : in    std_logic := 'U';
          CLKA    : in    std_logic := 'U';
          CLKB    : in    std_logic := 'U';
          RESET   : in    std_logic := 'U';
          DOUTA8  : out   std_logic;
          DOUTA7  : out   std_logic;
          DOUTA6  : out   std_logic;
          DOUTA5  : out   std_logic;
          DOUTA4  : out   std_logic;
          DOUTA3  : out   std_logic;
          DOUTA2  : out   std_logic;
          DOUTA1  : out   std_logic;
          DOUTA0  : out   std_logic;
          DOUTB8  : out   std_logic;
          DOUTB7  : out   std_logic;
          DOUTB6  : out   std_logic;
          DOUTB5  : out   std_logic;
          DOUTB4  : out   std_logic;
          DOUTB3  : out   std_logic;
          DOUTB2  : out   std_logic;
          DOUTB1  : out   std_logic;
          DOUTB0  : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \DOUTA_1[8]\, \DOUTB_1[8]\, DPRT_512X9_SRAM_3_GND, 
        DPRT_512X9_SRAM_3_VCC : std_logic;

begin 


    DPRT_512X9_SRAM_R0C0 : RAM4K9
      generic map(MEMORYFILE => "DPRT_512X9_SRAM_R0C0.mem")

      port map(ADDRA11 => DPRT_512X9_SRAM_3_GND, ADDRA10 => 
        DPRT_512X9_SRAM_3_GND, ADDRA9 => DPRT_512X9_SRAM_3_GND, 
        ADDRA8 => DPRT_512X9_SRAM_3_GND, ADDRA7 => 
        ELINK_ADDRA_3(7), ADDRA6 => ELINK_ADDRA_3(6), ADDRA5 => 
        ELINK_ADDRA_3(5), ADDRA4 => ELINK_ADDRA_3(4), ADDRA3 => 
        ELINK_ADDRA_3(3), ADDRA2 => ELINK_ADDRA_3(2), ADDRA1 => 
        ELINK_ADDRA_3(1), ADDRA0 => ELINK_ADDRA_3(0), ADDRB11 => 
        DPRT_512X9_SRAM_3_GND, ADDRB10 => DPRT_512X9_SRAM_3_GND, 
        ADDRB9 => DPRT_512X9_SRAM_3_GND, ADDRB8 => 
        DPRT_512X9_SRAM_3_GND, ADDRB7 => ELKS_ADDRB_7, ADDRB6 => 
        ELKS_ADDRB_0_4, ADDRB5 => ELKS_ADDRB_5, ADDRB4 => 
        ELKS_ADDRB_0_2, ADDRB3 => ELKS_ADDRB_3, ADDRB2 => 
        ELKS_ADDRB_0_0, ADDRB1 => ELKS_ADDRB_1, ADDRB0 => 
        ELKS_ADDRB_0_d0, DINA8 => DPRT_512X9_SRAM_3_GND, DINA7
         => ELINK_DINA_3(7), DINA6 => ELINK_DINA_3(6), DINA5 => 
        ELINK_DINA_3(5), DINA4 => ELINK_DINA_3(4), DINA3 => 
        ELINK_DINA_3(3), DINA2 => ELINK_DINA_3(2), DINA1 => 
        ELINK_DINA_3(1), DINA0 => ELINK_DINA_3(0), DINB8 => 
        DPRT_512X9_SRAM_3_GND, DINB7 => ELK_RX_SER_WORD_3(7), 
        DINB6 => ELK_RX_SER_WORD_3(6), DINB5 => 
        ELK_RX_SER_WORD_3(5), DINB4 => ELK_RX_SER_WORD_3(4), 
        DINB3 => ELK_RX_SER_WORD_3(3), DINB2 => 
        ELK_RX_SER_WORD_3(2), DINB1 => ELK_RX_SER_WORD_3(1), 
        DINB0 => ELK_RX_SER_WORD_3(0), WIDTHA0 => 
        DPRT_512X9_SRAM_3_VCC, WIDTHA1 => DPRT_512X9_SRAM_3_VCC, 
        WIDTHB0 => DPRT_512X9_SRAM_3_VCC, WIDTHB1 => 
        DPRT_512X9_SRAM_3_VCC, PIPEA => DPRT_512X9_SRAM_3_VCC, 
        PIPEB => DPRT_512X9_SRAM_3_VCC, WMODEA => 
        DPRT_512X9_SRAM_3_GND, WMODEB => DPRT_512X9_SRAM_3_GND, 
        BLKA => ELINK_BLKA_0, BLKB => ELKS_RAM_BLKB_EN, WENA => 
        ELINK_RWA_0, WENB => ELKS_RWB, CLKA => CLK60MHZ, CLKB => 
        CLK_40M_GL, RESET => P_USB_MASTER_EN_c_0, DOUTA8 => 
        \DOUTA_1[8]\, DOUTA7 => ELINK_DOUTA_3(7), DOUTA6 => 
        ELINK_DOUTA_3(6), DOUTA5 => ELINK_DOUTA_3(5), DOUTA4 => 
        ELINK_DOUTA_3(4), DOUTA3 => ELINK_DOUTA_3(3), DOUTA2 => 
        ELINK_DOUTA_3(2), DOUTA1 => ELINK_DOUTA_3(1), DOUTA0 => 
        ELINK_DOUTA_3(0), DOUTB8 => \DOUTB_1[8]\, DOUTB7 => 
        PATT_ELK_DAT_3(7), DOUTB6 => PATT_ELK_DAT_3(6), DOUTB5
         => PATT_ELK_DAT_3(5), DOUTB4 => PATT_ELK_DAT_3(4), 
        DOUTB3 => PATT_ELK_DAT_3(3), DOUTB2 => PATT_ELK_DAT_3(2), 
        DOUTB1 => PATT_ELK_DAT_3(1), DOUTB0 => PATT_ELK_DAT_3(0));
    
    VCC_i : VCC
      port map(Y => DPRT_512X9_SRAM_3_VCC);
    
    GND_i : GND
      port map(Y => DPRT_512X9_SRAM_3_GND);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity DPRT_512X9_SRAM_2 is

    port( ELINK_RWA_0         : in    std_logic;
          ELK_RX_SER_WORD_2   : in    std_logic_vector(7 downto 0);
          ELINK_DINA_2        : in    std_logic_vector(7 downto 0);
          ELINK_BLKA_0        : in    std_logic;
          ELKS_ADDRB          : in    std_logic_vector(7 downto 0);
          ELINK_ADDRA_2       : in    std_logic_vector(7 downto 0);
          PATT_ELK_DAT_2      : out   std_logic_vector(7 downto 0);
          ELINK_DOUTA_2       : out   std_logic_vector(7 downto 0);
          ELKS_RWB            : in    std_logic;
          P_USB_MASTER_EN_c_0 : in    std_logic;
          CLK_40M_GL          : in    std_logic;
          CLK60MHZ            : in    std_logic;
          ELKS_RAM_BLKB_EN    : in    std_logic
        );

end DPRT_512X9_SRAM_2;

architecture DEF_ARCH of DPRT_512X9_SRAM_2 is 

  component RAM4K9
    generic (MEMORYFILE:string := "");

    port( ADDRA11 : in    std_logic := 'U';
          ADDRA10 : in    std_logic := 'U';
          ADDRA9  : in    std_logic := 'U';
          ADDRA8  : in    std_logic := 'U';
          ADDRA7  : in    std_logic := 'U';
          ADDRA6  : in    std_logic := 'U';
          ADDRA5  : in    std_logic := 'U';
          ADDRA4  : in    std_logic := 'U';
          ADDRA3  : in    std_logic := 'U';
          ADDRA2  : in    std_logic := 'U';
          ADDRA1  : in    std_logic := 'U';
          ADDRA0  : in    std_logic := 'U';
          ADDRB11 : in    std_logic := 'U';
          ADDRB10 : in    std_logic := 'U';
          ADDRB9  : in    std_logic := 'U';
          ADDRB8  : in    std_logic := 'U';
          ADDRB7  : in    std_logic := 'U';
          ADDRB6  : in    std_logic := 'U';
          ADDRB5  : in    std_logic := 'U';
          ADDRB4  : in    std_logic := 'U';
          ADDRB3  : in    std_logic := 'U';
          ADDRB2  : in    std_logic := 'U';
          ADDRB1  : in    std_logic := 'U';
          ADDRB0  : in    std_logic := 'U';
          DINA8   : in    std_logic := 'U';
          DINA7   : in    std_logic := 'U';
          DINA6   : in    std_logic := 'U';
          DINA5   : in    std_logic := 'U';
          DINA4   : in    std_logic := 'U';
          DINA3   : in    std_logic := 'U';
          DINA2   : in    std_logic := 'U';
          DINA1   : in    std_logic := 'U';
          DINA0   : in    std_logic := 'U';
          DINB8   : in    std_logic := 'U';
          DINB7   : in    std_logic := 'U';
          DINB6   : in    std_logic := 'U';
          DINB5   : in    std_logic := 'U';
          DINB4   : in    std_logic := 'U';
          DINB3   : in    std_logic := 'U';
          DINB2   : in    std_logic := 'U';
          DINB1   : in    std_logic := 'U';
          DINB0   : in    std_logic := 'U';
          WIDTHA0 : in    std_logic := 'U';
          WIDTHA1 : in    std_logic := 'U';
          WIDTHB0 : in    std_logic := 'U';
          WIDTHB1 : in    std_logic := 'U';
          PIPEA   : in    std_logic := 'U';
          PIPEB   : in    std_logic := 'U';
          WMODEA  : in    std_logic := 'U';
          WMODEB  : in    std_logic := 'U';
          BLKA    : in    std_logic := 'U';
          BLKB    : in    std_logic := 'U';
          WENA    : in    std_logic := 'U';
          WENB    : in    std_logic := 'U';
          CLKA    : in    std_logic := 'U';
          CLKB    : in    std_logic := 'U';
          RESET   : in    std_logic := 'U';
          DOUTA8  : out   std_logic;
          DOUTA7  : out   std_logic;
          DOUTA6  : out   std_logic;
          DOUTA5  : out   std_logic;
          DOUTA4  : out   std_logic;
          DOUTA3  : out   std_logic;
          DOUTA2  : out   std_logic;
          DOUTA1  : out   std_logic;
          DOUTA0  : out   std_logic;
          DOUTB8  : out   std_logic;
          DOUTB7  : out   std_logic;
          DOUTB6  : out   std_logic;
          DOUTB5  : out   std_logic;
          DOUTB4  : out   std_logic;
          DOUTB3  : out   std_logic;
          DOUTB2  : out   std_logic;
          DOUTB1  : out   std_logic;
          DOUTB0  : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \DOUTA_1[8]\, \DOUTB_1[8]\, DPRT_512X9_SRAM_2_GND, 
        DPRT_512X9_SRAM_2_VCC : std_logic;

begin 


    DPRT_512X9_SRAM_R0C0 : RAM4K9
      generic map(MEMORYFILE => "DPRT_512X9_SRAM_R0C0.mem")

      port map(ADDRA11 => DPRT_512X9_SRAM_2_GND, ADDRA10 => 
        DPRT_512X9_SRAM_2_GND, ADDRA9 => DPRT_512X9_SRAM_2_GND, 
        ADDRA8 => DPRT_512X9_SRAM_2_GND, ADDRA7 => 
        ELINK_ADDRA_2(7), ADDRA6 => ELINK_ADDRA_2(6), ADDRA5 => 
        ELINK_ADDRA_2(5), ADDRA4 => ELINK_ADDRA_2(4), ADDRA3 => 
        ELINK_ADDRA_2(3), ADDRA2 => ELINK_ADDRA_2(2), ADDRA1 => 
        ELINK_ADDRA_2(1), ADDRA0 => ELINK_ADDRA_2(0), ADDRB11 => 
        DPRT_512X9_SRAM_2_GND, ADDRB10 => DPRT_512X9_SRAM_2_GND, 
        ADDRB9 => DPRT_512X9_SRAM_2_GND, ADDRB8 => 
        DPRT_512X9_SRAM_2_GND, ADDRB7 => ELKS_ADDRB(7), ADDRB6
         => ELKS_ADDRB(6), ADDRB5 => ELKS_ADDRB(5), ADDRB4 => 
        ELKS_ADDRB(4), ADDRB3 => ELKS_ADDRB(3), ADDRB2 => 
        ELKS_ADDRB(2), ADDRB1 => ELKS_ADDRB(1), ADDRB0 => 
        ELKS_ADDRB(0), DINA8 => DPRT_512X9_SRAM_2_GND, DINA7 => 
        ELINK_DINA_2(7), DINA6 => ELINK_DINA_2(6), DINA5 => 
        ELINK_DINA_2(5), DINA4 => ELINK_DINA_2(4), DINA3 => 
        ELINK_DINA_2(3), DINA2 => ELINK_DINA_2(2), DINA1 => 
        ELINK_DINA_2(1), DINA0 => ELINK_DINA_2(0), DINB8 => 
        DPRT_512X9_SRAM_2_GND, DINB7 => ELK_RX_SER_WORD_2(7), 
        DINB6 => ELK_RX_SER_WORD_2(6), DINB5 => 
        ELK_RX_SER_WORD_2(5), DINB4 => ELK_RX_SER_WORD_2(4), 
        DINB3 => ELK_RX_SER_WORD_2(3), DINB2 => 
        ELK_RX_SER_WORD_2(2), DINB1 => ELK_RX_SER_WORD_2(1), 
        DINB0 => ELK_RX_SER_WORD_2(0), WIDTHA0 => 
        DPRT_512X9_SRAM_2_VCC, WIDTHA1 => DPRT_512X9_SRAM_2_VCC, 
        WIDTHB0 => DPRT_512X9_SRAM_2_VCC, WIDTHB1 => 
        DPRT_512X9_SRAM_2_VCC, PIPEA => DPRT_512X9_SRAM_2_VCC, 
        PIPEB => DPRT_512X9_SRAM_2_VCC, WMODEA => 
        DPRT_512X9_SRAM_2_GND, WMODEB => DPRT_512X9_SRAM_2_GND, 
        BLKA => ELINK_BLKA_0, BLKB => ELKS_RAM_BLKB_EN, WENA => 
        ELINK_RWA_0, WENB => ELKS_RWB, CLKA => CLK60MHZ, CLKB => 
        CLK_40M_GL, RESET => P_USB_MASTER_EN_c_0, DOUTA8 => 
        \DOUTA_1[8]\, DOUTA7 => ELINK_DOUTA_2(7), DOUTA6 => 
        ELINK_DOUTA_2(6), DOUTA5 => ELINK_DOUTA_2(5), DOUTA4 => 
        ELINK_DOUTA_2(4), DOUTA3 => ELINK_DOUTA_2(3), DOUTA2 => 
        ELINK_DOUTA_2(2), DOUTA1 => ELINK_DOUTA_2(1), DOUTA0 => 
        ELINK_DOUTA_2(0), DOUTB8 => \DOUTB_1[8]\, DOUTB7 => 
        PATT_ELK_DAT_2(7), DOUTB6 => PATT_ELK_DAT_2(6), DOUTB5
         => PATT_ELK_DAT_2(5), DOUTB4 => PATT_ELK_DAT_2(4), 
        DOUTB3 => PATT_ELK_DAT_2(3), DOUTB2 => PATT_ELK_DAT_2(2), 
        DOUTB1 => PATT_ELK_DAT_2(1), DOUTB0 => PATT_ELK_DAT_2(0));
    
    VCC_i : VCC
      port map(Y => DPRT_512X9_SRAM_2_VCC);
    
    GND_i : GND
      port map(Y => DPRT_512X9_SRAM_2_GND);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity DPRT_512X9_SRAM_1 is

    port( ELINK_RWA_0         : in    std_logic;
          ELK_RX_SER_WORD_1   : in    std_logic_vector(7 downto 0);
          ELINK_DINA_1        : in    std_logic_vector(7 downto 0);
          ELINK_BLKA_0        : in    std_logic;
          ELKS_ADDRB_0_d0     : in    std_logic;
          ELKS_ADDRB_1        : in    std_logic;
          ELKS_ADDRB_3        : in    std_logic;
          ELKS_ADDRB_5        : in    std_logic;
          ELKS_ADDRB_7        : in    std_logic;
          ELKS_ADDRB_0_0      : in    std_logic;
          ELKS_ADDRB_0_2      : in    std_logic;
          ELKS_ADDRB_0_4      : in    std_logic;
          ELINK_ADDRA_1       : in    std_logic_vector(7 downto 0);
          PATT_ELK_DAT_1      : out   std_logic_vector(7 downto 0);
          ELINK_DOUTA_1       : out   std_logic_vector(7 downto 0);
          ELKS_RWB            : in    std_logic;
          P_USB_MASTER_EN_c_0 : in    std_logic;
          CLK_40M_GL          : in    std_logic;
          CLK60MHZ            : in    std_logic;
          ELKS_RAM_BLKB_EN    : in    std_logic
        );

end DPRT_512X9_SRAM_1;

architecture DEF_ARCH of DPRT_512X9_SRAM_1 is 

  component RAM4K9
    generic (MEMORYFILE:string := "");

    port( ADDRA11 : in    std_logic := 'U';
          ADDRA10 : in    std_logic := 'U';
          ADDRA9  : in    std_logic := 'U';
          ADDRA8  : in    std_logic := 'U';
          ADDRA7  : in    std_logic := 'U';
          ADDRA6  : in    std_logic := 'U';
          ADDRA5  : in    std_logic := 'U';
          ADDRA4  : in    std_logic := 'U';
          ADDRA3  : in    std_logic := 'U';
          ADDRA2  : in    std_logic := 'U';
          ADDRA1  : in    std_logic := 'U';
          ADDRA0  : in    std_logic := 'U';
          ADDRB11 : in    std_logic := 'U';
          ADDRB10 : in    std_logic := 'U';
          ADDRB9  : in    std_logic := 'U';
          ADDRB8  : in    std_logic := 'U';
          ADDRB7  : in    std_logic := 'U';
          ADDRB6  : in    std_logic := 'U';
          ADDRB5  : in    std_logic := 'U';
          ADDRB4  : in    std_logic := 'U';
          ADDRB3  : in    std_logic := 'U';
          ADDRB2  : in    std_logic := 'U';
          ADDRB1  : in    std_logic := 'U';
          ADDRB0  : in    std_logic := 'U';
          DINA8   : in    std_logic := 'U';
          DINA7   : in    std_logic := 'U';
          DINA6   : in    std_logic := 'U';
          DINA5   : in    std_logic := 'U';
          DINA4   : in    std_logic := 'U';
          DINA3   : in    std_logic := 'U';
          DINA2   : in    std_logic := 'U';
          DINA1   : in    std_logic := 'U';
          DINA0   : in    std_logic := 'U';
          DINB8   : in    std_logic := 'U';
          DINB7   : in    std_logic := 'U';
          DINB6   : in    std_logic := 'U';
          DINB5   : in    std_logic := 'U';
          DINB4   : in    std_logic := 'U';
          DINB3   : in    std_logic := 'U';
          DINB2   : in    std_logic := 'U';
          DINB1   : in    std_logic := 'U';
          DINB0   : in    std_logic := 'U';
          WIDTHA0 : in    std_logic := 'U';
          WIDTHA1 : in    std_logic := 'U';
          WIDTHB0 : in    std_logic := 'U';
          WIDTHB1 : in    std_logic := 'U';
          PIPEA   : in    std_logic := 'U';
          PIPEB   : in    std_logic := 'U';
          WMODEA  : in    std_logic := 'U';
          WMODEB  : in    std_logic := 'U';
          BLKA    : in    std_logic := 'U';
          BLKB    : in    std_logic := 'U';
          WENA    : in    std_logic := 'U';
          WENB    : in    std_logic := 'U';
          CLKA    : in    std_logic := 'U';
          CLKB    : in    std_logic := 'U';
          RESET   : in    std_logic := 'U';
          DOUTA8  : out   std_logic;
          DOUTA7  : out   std_logic;
          DOUTA6  : out   std_logic;
          DOUTA5  : out   std_logic;
          DOUTA4  : out   std_logic;
          DOUTA3  : out   std_logic;
          DOUTA2  : out   std_logic;
          DOUTA1  : out   std_logic;
          DOUTA0  : out   std_logic;
          DOUTB8  : out   std_logic;
          DOUTB7  : out   std_logic;
          DOUTB6  : out   std_logic;
          DOUTB5  : out   std_logic;
          DOUTB4  : out   std_logic;
          DOUTB3  : out   std_logic;
          DOUTB2  : out   std_logic;
          DOUTB1  : out   std_logic;
          DOUTB0  : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \DOUTA_1[8]\, \DOUTB_1[8]\, DPRT_512X9_SRAM_1_GND, 
        DPRT_512X9_SRAM_1_VCC : std_logic;

begin 


    DPRT_512X9_SRAM_R0C0 : RAM4K9
      generic map(MEMORYFILE => "DPRT_512X9_SRAM_R0C0.mem")

      port map(ADDRA11 => DPRT_512X9_SRAM_1_GND, ADDRA10 => 
        DPRT_512X9_SRAM_1_GND, ADDRA9 => DPRT_512X9_SRAM_1_GND, 
        ADDRA8 => DPRT_512X9_SRAM_1_GND, ADDRA7 => 
        ELINK_ADDRA_1(7), ADDRA6 => ELINK_ADDRA_1(6), ADDRA5 => 
        ELINK_ADDRA_1(5), ADDRA4 => ELINK_ADDRA_1(4), ADDRA3 => 
        ELINK_ADDRA_1(3), ADDRA2 => ELINK_ADDRA_1(2), ADDRA1 => 
        ELINK_ADDRA_1(1), ADDRA0 => ELINK_ADDRA_1(0), ADDRB11 => 
        DPRT_512X9_SRAM_1_GND, ADDRB10 => DPRT_512X9_SRAM_1_GND, 
        ADDRB9 => DPRT_512X9_SRAM_1_GND, ADDRB8 => 
        DPRT_512X9_SRAM_1_GND, ADDRB7 => ELKS_ADDRB_7, ADDRB6 => 
        ELKS_ADDRB_0_4, ADDRB5 => ELKS_ADDRB_5, ADDRB4 => 
        ELKS_ADDRB_0_2, ADDRB3 => ELKS_ADDRB_3, ADDRB2 => 
        ELKS_ADDRB_0_0, ADDRB1 => ELKS_ADDRB_1, ADDRB0 => 
        ELKS_ADDRB_0_d0, DINA8 => DPRT_512X9_SRAM_1_GND, DINA7
         => ELINK_DINA_1(7), DINA6 => ELINK_DINA_1(6), DINA5 => 
        ELINK_DINA_1(5), DINA4 => ELINK_DINA_1(4), DINA3 => 
        ELINK_DINA_1(3), DINA2 => ELINK_DINA_1(2), DINA1 => 
        ELINK_DINA_1(1), DINA0 => ELINK_DINA_1(0), DINB8 => 
        DPRT_512X9_SRAM_1_GND, DINB7 => ELK_RX_SER_WORD_1(7), 
        DINB6 => ELK_RX_SER_WORD_1(6), DINB5 => 
        ELK_RX_SER_WORD_1(5), DINB4 => ELK_RX_SER_WORD_1(4), 
        DINB3 => ELK_RX_SER_WORD_1(3), DINB2 => 
        ELK_RX_SER_WORD_1(2), DINB1 => ELK_RX_SER_WORD_1(1), 
        DINB0 => ELK_RX_SER_WORD_1(0), WIDTHA0 => 
        DPRT_512X9_SRAM_1_VCC, WIDTHA1 => DPRT_512X9_SRAM_1_VCC, 
        WIDTHB0 => DPRT_512X9_SRAM_1_VCC, WIDTHB1 => 
        DPRT_512X9_SRAM_1_VCC, PIPEA => DPRT_512X9_SRAM_1_VCC, 
        PIPEB => DPRT_512X9_SRAM_1_VCC, WMODEA => 
        DPRT_512X9_SRAM_1_GND, WMODEB => DPRT_512X9_SRAM_1_GND, 
        BLKA => ELINK_BLKA_0, BLKB => ELKS_RAM_BLKB_EN, WENA => 
        ELINK_RWA_0, WENB => ELKS_RWB, CLKA => CLK60MHZ, CLKB => 
        CLK_40M_GL, RESET => P_USB_MASTER_EN_c_0, DOUTA8 => 
        \DOUTA_1[8]\, DOUTA7 => ELINK_DOUTA_1(7), DOUTA6 => 
        ELINK_DOUTA_1(6), DOUTA5 => ELINK_DOUTA_1(5), DOUTA4 => 
        ELINK_DOUTA_1(4), DOUTA3 => ELINK_DOUTA_1(3), DOUTA2 => 
        ELINK_DOUTA_1(2), DOUTA1 => ELINK_DOUTA_1(1), DOUTA0 => 
        ELINK_DOUTA_1(0), DOUTB8 => \DOUTB_1[8]\, DOUTB7 => 
        PATT_ELK_DAT_1(7), DOUTB6 => PATT_ELK_DAT_1(6), DOUTB5
         => PATT_ELK_DAT_1(5), DOUTB4 => PATT_ELK_DAT_1(4), 
        DOUTB3 => PATT_ELK_DAT_1(3), DOUTB2 => PATT_ELK_DAT_1(2), 
        DOUTB1 => PATT_ELK_DAT_1(1), DOUTB0 => PATT_ELK_DAT_1(0));
    
    VCC_i : VCC
      port map(Y => DPRT_512X9_SRAM_1_VCC);
    
    GND_i : GND
      port map(Y => DPRT_512X9_SRAM_1_GND);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity DPRT_512X9_SRAM_6 is

    port( ELINK_RWA_0         : in    std_logic;
          ELK_RX_SER_WORD_6   : in    std_logic_vector(7 downto 0);
          ELINK_DINA_6        : in    std_logic_vector(7 downto 0);
          ELINK_BLKA_0        : in    std_logic;
          ELKS_ADDRB_0_d0     : in    std_logic;
          ELKS_ADDRB_1        : in    std_logic;
          ELKS_ADDRB_3        : in    std_logic;
          ELKS_ADDRB_5        : in    std_logic;
          ELKS_ADDRB_7        : in    std_logic;
          ELKS_ADDRB_0_0      : in    std_logic;
          ELKS_ADDRB_0_2      : in    std_logic;
          ELKS_ADDRB_0_4      : in    std_logic;
          ELINK_ADDRA_6       : in    std_logic_vector(7 downto 0);
          PATT_ELK_DAT_6      : out   std_logic_vector(7 downto 0);
          ELINK_DOUTA_6       : out   std_logic_vector(7 downto 0);
          ELKS_RWB            : in    std_logic;
          P_USB_MASTER_EN_c_0 : in    std_logic;
          CLK_40M_GL          : in    std_logic;
          CLK60MHZ            : in    std_logic;
          ELKS_RAM_BLKB_EN    : in    std_logic
        );

end DPRT_512X9_SRAM_6;

architecture DEF_ARCH of DPRT_512X9_SRAM_6 is 

  component RAM4K9
    generic (MEMORYFILE:string := "");

    port( ADDRA11 : in    std_logic := 'U';
          ADDRA10 : in    std_logic := 'U';
          ADDRA9  : in    std_logic := 'U';
          ADDRA8  : in    std_logic := 'U';
          ADDRA7  : in    std_logic := 'U';
          ADDRA6  : in    std_logic := 'U';
          ADDRA5  : in    std_logic := 'U';
          ADDRA4  : in    std_logic := 'U';
          ADDRA3  : in    std_logic := 'U';
          ADDRA2  : in    std_logic := 'U';
          ADDRA1  : in    std_logic := 'U';
          ADDRA0  : in    std_logic := 'U';
          ADDRB11 : in    std_logic := 'U';
          ADDRB10 : in    std_logic := 'U';
          ADDRB9  : in    std_logic := 'U';
          ADDRB8  : in    std_logic := 'U';
          ADDRB7  : in    std_logic := 'U';
          ADDRB6  : in    std_logic := 'U';
          ADDRB5  : in    std_logic := 'U';
          ADDRB4  : in    std_logic := 'U';
          ADDRB3  : in    std_logic := 'U';
          ADDRB2  : in    std_logic := 'U';
          ADDRB1  : in    std_logic := 'U';
          ADDRB0  : in    std_logic := 'U';
          DINA8   : in    std_logic := 'U';
          DINA7   : in    std_logic := 'U';
          DINA6   : in    std_logic := 'U';
          DINA5   : in    std_logic := 'U';
          DINA4   : in    std_logic := 'U';
          DINA3   : in    std_logic := 'U';
          DINA2   : in    std_logic := 'U';
          DINA1   : in    std_logic := 'U';
          DINA0   : in    std_logic := 'U';
          DINB8   : in    std_logic := 'U';
          DINB7   : in    std_logic := 'U';
          DINB6   : in    std_logic := 'U';
          DINB5   : in    std_logic := 'U';
          DINB4   : in    std_logic := 'U';
          DINB3   : in    std_logic := 'U';
          DINB2   : in    std_logic := 'U';
          DINB1   : in    std_logic := 'U';
          DINB0   : in    std_logic := 'U';
          WIDTHA0 : in    std_logic := 'U';
          WIDTHA1 : in    std_logic := 'U';
          WIDTHB0 : in    std_logic := 'U';
          WIDTHB1 : in    std_logic := 'U';
          PIPEA   : in    std_logic := 'U';
          PIPEB   : in    std_logic := 'U';
          WMODEA  : in    std_logic := 'U';
          WMODEB  : in    std_logic := 'U';
          BLKA    : in    std_logic := 'U';
          BLKB    : in    std_logic := 'U';
          WENA    : in    std_logic := 'U';
          WENB    : in    std_logic := 'U';
          CLKA    : in    std_logic := 'U';
          CLKB    : in    std_logic := 'U';
          RESET   : in    std_logic := 'U';
          DOUTA8  : out   std_logic;
          DOUTA7  : out   std_logic;
          DOUTA6  : out   std_logic;
          DOUTA5  : out   std_logic;
          DOUTA4  : out   std_logic;
          DOUTA3  : out   std_logic;
          DOUTA2  : out   std_logic;
          DOUTA1  : out   std_logic;
          DOUTA0  : out   std_logic;
          DOUTB8  : out   std_logic;
          DOUTB7  : out   std_logic;
          DOUTB6  : out   std_logic;
          DOUTB5  : out   std_logic;
          DOUTB4  : out   std_logic;
          DOUTB3  : out   std_logic;
          DOUTB2  : out   std_logic;
          DOUTB1  : out   std_logic;
          DOUTB0  : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \DOUTA_1[8]\, \DOUTB_1[8]\, DPRT_512X9_SRAM_6_GND, 
        DPRT_512X9_SRAM_6_VCC : std_logic;

begin 


    DPRT_512X9_SRAM_R0C0 : RAM4K9
      generic map(MEMORYFILE => "DPRT_512X9_SRAM_R0C0.mem")

      port map(ADDRA11 => DPRT_512X9_SRAM_6_GND, ADDRA10 => 
        DPRT_512X9_SRAM_6_GND, ADDRA9 => DPRT_512X9_SRAM_6_GND, 
        ADDRA8 => DPRT_512X9_SRAM_6_GND, ADDRA7 => 
        ELINK_ADDRA_6(7), ADDRA6 => ELINK_ADDRA_6(6), ADDRA5 => 
        ELINK_ADDRA_6(5), ADDRA4 => ELINK_ADDRA_6(4), ADDRA3 => 
        ELINK_ADDRA_6(3), ADDRA2 => ELINK_ADDRA_6(2), ADDRA1 => 
        ELINK_ADDRA_6(1), ADDRA0 => ELINK_ADDRA_6(0), ADDRB11 => 
        DPRT_512X9_SRAM_6_GND, ADDRB10 => DPRT_512X9_SRAM_6_GND, 
        ADDRB9 => DPRT_512X9_SRAM_6_GND, ADDRB8 => 
        DPRT_512X9_SRAM_6_GND, ADDRB7 => ELKS_ADDRB_7, ADDRB6 => 
        ELKS_ADDRB_0_4, ADDRB5 => ELKS_ADDRB_5, ADDRB4 => 
        ELKS_ADDRB_0_2, ADDRB3 => ELKS_ADDRB_3, ADDRB2 => 
        ELKS_ADDRB_0_0, ADDRB1 => ELKS_ADDRB_1, ADDRB0 => 
        ELKS_ADDRB_0_d0, DINA8 => DPRT_512X9_SRAM_6_GND, DINA7
         => ELINK_DINA_6(7), DINA6 => ELINK_DINA_6(6), DINA5 => 
        ELINK_DINA_6(5), DINA4 => ELINK_DINA_6(4), DINA3 => 
        ELINK_DINA_6(3), DINA2 => ELINK_DINA_6(2), DINA1 => 
        ELINK_DINA_6(1), DINA0 => ELINK_DINA_6(0), DINB8 => 
        DPRT_512X9_SRAM_6_GND, DINB7 => ELK_RX_SER_WORD_6(7), 
        DINB6 => ELK_RX_SER_WORD_6(6), DINB5 => 
        ELK_RX_SER_WORD_6(5), DINB4 => ELK_RX_SER_WORD_6(4), 
        DINB3 => ELK_RX_SER_WORD_6(3), DINB2 => 
        ELK_RX_SER_WORD_6(2), DINB1 => ELK_RX_SER_WORD_6(1), 
        DINB0 => ELK_RX_SER_WORD_6(0), WIDTHA0 => 
        DPRT_512X9_SRAM_6_VCC, WIDTHA1 => DPRT_512X9_SRAM_6_VCC, 
        WIDTHB0 => DPRT_512X9_SRAM_6_VCC, WIDTHB1 => 
        DPRT_512X9_SRAM_6_VCC, PIPEA => DPRT_512X9_SRAM_6_VCC, 
        PIPEB => DPRT_512X9_SRAM_6_VCC, WMODEA => 
        DPRT_512X9_SRAM_6_GND, WMODEB => DPRT_512X9_SRAM_6_GND, 
        BLKA => ELINK_BLKA_0, BLKB => ELKS_RAM_BLKB_EN, WENA => 
        ELINK_RWA_0, WENB => ELKS_RWB, CLKA => CLK60MHZ, CLKB => 
        CLK_40M_GL, RESET => P_USB_MASTER_EN_c_0, DOUTA8 => 
        \DOUTA_1[8]\, DOUTA7 => ELINK_DOUTA_6(7), DOUTA6 => 
        ELINK_DOUTA_6(6), DOUTA5 => ELINK_DOUTA_6(5), DOUTA4 => 
        ELINK_DOUTA_6(4), DOUTA3 => ELINK_DOUTA_6(3), DOUTA2 => 
        ELINK_DOUTA_6(2), DOUTA1 => ELINK_DOUTA_6(1), DOUTA0 => 
        ELINK_DOUTA_6(0), DOUTB8 => \DOUTB_1[8]\, DOUTB7 => 
        PATT_ELK_DAT_6(7), DOUTB6 => PATT_ELK_DAT_6(6), DOUTB5
         => PATT_ELK_DAT_6(5), DOUTB4 => PATT_ELK_DAT_6(4), 
        DOUTB3 => PATT_ELK_DAT_6(3), DOUTB2 => PATT_ELK_DAT_6(2), 
        DOUTB1 => PATT_ELK_DAT_6(1), DOUTB0 => PATT_ELK_DAT_6(0));
    
    VCC_i : VCC
      port map(Y => DPRT_512X9_SRAM_6_VCC);
    
    GND_i : GND
      port map(Y => DPRT_512X9_SRAM_6_GND);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity CLK60M_TO_40M_0 is

    port( OP_MODE              : inout std_logic_vector(7 downto 0) := (others => 'Z');
          OP_MODE_0_0          : in    std_logic;
          OP_MODE_0_4          : in    std_logic;
          OP_MODE_c_1_d0       : out   std_logic;
          OP_MODE_c_5_d0       : out   std_logic;
          OP_MODE_c_4_d0       : out   std_logic;
          OP_MODE_c_0_d0       : out   std_logic;
          OP_MODE_c_0_0        : out   std_logic;
          OP_MODE_c_1_0        : out   std_logic;
          OP_MODE_c_2_0        : out   std_logic;
          OP_MODE_c_3_0        : out   std_logic;
          OP_MODE_c_4_0        : out   std_logic;
          OP_MODE_c_5_0        : out   std_logic;
          OP_MODE_c_6_0        : out   std_logic;
          P_MASTER_POR_B_c_25  : in    std_logic;
          P_MASTER_POR_B_c_24  : in    std_logic;
          P_MASTER_POR_B_c_23  : in    std_logic;
          P_MASTER_POR_B_c_6   : in    std_logic;
          P_MASTER_POR_B_c     : in    std_logic;
          P_MASTER_POR_B_c_1   : in    std_logic;
          P_MASTER_POR_B_c_0_0 : in    std_logic;
          CLK_40M_GL           : in    std_logic
        );

end CLK60M_TO_40M_0;

architecture DEF_ARCH of CLK60M_TO_40M_0 is 

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XO1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component OR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component MX2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \OP_MODE_c_6[1]\, \SAMP_TWO[1]_net_1\, un7_delcnt, 
        un1_SAMP_TWO_NE_4, un1_SAMP_TWO_0, un1_SAMP_TWO_NE_0, 
        un1_SAMP_TWO_NE_2, un1_SAMP_TWO_NE_3, \OP_MODE_c[2]\, 
        \SAMP_TWO[2]_net_1\, un1_SAMP_TWO_6, \SAMP_TWO[4]_net_1\, 
        un1_SAMP_TWO_5, \SAMP_TWO[3]_net_1\, 
        \LOCAL_REG_VAL[3]_net_1\, un1_SAMP_TWO_7, n_sync_sm3, 
        un1_SAMP_TWO_1, \N_DELCNT[0]\, \SYNC_SM[0]_net_1\, 
        \DELCNT[0]_net_1\, \DELCNT[1]_net_1\, \N_SYNC_SM[0]\, 
        \LOCAL_REG_VAL[7]_net_1\, \SAMP_TWO[7]_net_1\, 
        \SAMP_TWO[6]_net_1\, \OP_MODE_c[6]\, \SAMP_TWO[5]_net_1\, 
        \OP_MODE_c[5]\, \SAMP_TWO[0]_net_1\, SUM1_4, 
        \SAMP_ONE[0]_net_1\, \SAMP_ONE[1]_net_1\, 
        \SAMP_ONE[2]_net_1\, \SAMP_ONE[3]_net_1\, 
        \SAMP_ONE[4]_net_1\, \SAMP_ONE[5]_net_1\, 
        \SAMP_ONE[6]_net_1\, \SAMP_ONE[7]_net_1\, \GND\, \VCC\
         : std_logic;

begin 

    OP_MODE_c_1_d0 <= \OP_MODE_c[2]\;
    OP_MODE_c_5_d0 <= \OP_MODE_c[6]\;
    OP_MODE_c_4_d0 <= \OP_MODE_c[5]\;
    OP_MODE_c_6_0 <= \OP_MODE_c_6[1]\;

    \SAMP_ONE[2]\ : DFN1C0
      port map(D => OP_MODE(2), CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c, Q => \SAMP_ONE[2]_net_1\);
    
    \DELCNT_RNIR2EA[1]\ : NOR2B
      port map(A => \DELCNT[1]_net_1\, B => \DELCNT[0]_net_1\, Y
         => un7_delcnt);
    
    \SYNC_SM_RNO_6[0]\ : XO1
      port map(A => OP_MODE(4), B => \SAMP_TWO[4]_net_1\, C => 
        un1_SAMP_TWO_5, Y => un1_SAMP_TWO_NE_2);
    
    \LOCAL_REG_VAL[3]\ : DFN1E1C0
      port map(D => \SAMP_TWO[3]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_6, E => un7_delcnt, Q => 
        \LOCAL_REG_VAL[3]_net_1\);
    
    \SYNC_SM[0]\ : DFN1C0
      port map(D => \N_SYNC_SM[0]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c, Q => \SYNC_SM[0]_net_1\);
    
    \SYNC_SM_RNO_5[0]\ : XO1
      port map(A => \SAMP_TWO[3]_net_1\, B => 
        \LOCAL_REG_VAL[3]_net_1\, C => un1_SAMP_TWO_7, Y => 
        un1_SAMP_TWO_NE_0);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \DELCNT[1]\ : DFN1C0
      port map(D => SUM1_4, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_25, Q => \DELCNT[1]_net_1\);
    
    \LOCAL_REG_VAL_6[1]\ : DFN1E1C0
      port map(D => \SAMP_TWO[1]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_0_0, E => un7_delcnt, Q => 
        \OP_MODE_c_6[1]\);
    
    \LOCAL_REG_VAL[5]\ : DFN1E1C0
      port map(D => \SAMP_TWO[5]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_6, E => un7_delcnt, Q => 
        \OP_MODE_c[5]\);
    
    \SYNC_SM_RNO_1[0]\ : OR3
      port map(A => un1_SAMP_TWO_0, B => un1_SAMP_TWO_NE_0, C => 
        un1_SAMP_TWO_NE_2, Y => un1_SAMP_TWO_NE_4);
    
    \SAMP_TWO[0]\ : DFN1C0
      port map(D => \SAMP_ONE[0]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_23, Q => \SAMP_TWO[0]_net_1\);
    
    \SAMP_ONE[1]\ : DFN1C0
      port map(D => OP_MODE(1), CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c, Q => \SAMP_ONE[1]_net_1\);
    
    \SAMP_TWO[1]\ : DFN1C0
      port map(D => \SAMP_ONE[1]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_23, Q => \SAMP_TWO[1]_net_1\);
    
    \SYNC_SM_RNO_3[0]\ : XOR2
      port map(A => \SAMP_TWO[1]_net_1\, B => \OP_MODE_c_6[1]\, Y
         => un1_SAMP_TWO_1);
    
    \LOCAL_REG_VAL_5[1]\ : DFN1E1C0
      port map(D => \SAMP_TWO[1]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_1, E => un7_delcnt, Q => 
        OP_MODE_c_5_0);
    
    \SYNC_SM_RNO_9[0]\ : XOR2
      port map(A => \SAMP_TWO[5]_net_1\, B => \OP_MODE_c[5]\, Y
         => un1_SAMP_TWO_5);
    
    \LOCAL_REG_VAL_1[1]\ : DFN1E1C0
      port map(D => \SAMP_TWO[1]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_1, E => un7_delcnt, Q => 
        OP_MODE_c_1_0);
    
    un2_n_delcnt_1_1_SUM1 : XOR2
      port map(A => \DELCNT[1]_net_1\, B => \DELCNT[0]_net_1\, Y
         => SUM1_4);
    
    \SAMP_TWO[3]\ : DFN1C0
      port map(D => \SAMP_ONE[3]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_23, Q => \SAMP_TWO[3]_net_1\);
    
    \SYNC_SM_RNO_8[0]\ : XOR2
      port map(A => \LOCAL_REG_VAL[7]_net_1\, B => 
        \SAMP_TWO[7]_net_1\, Y => un1_SAMP_TWO_7);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \SYNC_SM_RNO_4[0]\ : XOR2
      port map(A => \SAMP_TWO[0]_net_1\, B => OP_MODE(0), Y => 
        un1_SAMP_TWO_0);
    
    \SYNC_SM_RNO[0]\ : MX2B
      port map(A => n_sync_sm3, B => un7_delcnt, S => 
        \SYNC_SM[0]_net_1\, Y => \N_SYNC_SM[0]\);
    
    \SAMP_ONE[4]\ : DFN1C0
      port map(D => OP_MODE_0_4, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c, Q => \SAMP_ONE[4]_net_1\);
    
    \LOCAL_REG_VAL[2]\ : DFN1E1C0
      port map(D => \SAMP_TWO[2]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_6, E => un7_delcnt, Q => 
        \OP_MODE_c[2]\);
    
    \SAMP_TWO[5]\ : DFN1C0
      port map(D => \SAMP_ONE[5]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_24, Q => \SAMP_TWO[5]_net_1\);
    
    \SAMP_TWO[4]\ : DFN1C0
      port map(D => \SAMP_ONE[4]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_23, Q => \SAMP_TWO[4]_net_1\);
    
    \SAMP_TWO[2]\ : DFN1C0
      port map(D => \SAMP_ONE[2]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_23, Q => \SAMP_TWO[2]_net_1\);
    
    \DELCNT_RNO[0]\ : NOR2A
      port map(A => \SYNC_SM[0]_net_1\, B => \DELCNT[0]_net_1\, Y
         => \N_DELCNT[0]\);
    
    \LOCAL_REG_VAL_4[1]\ : DFN1E1C0
      port map(D => \SAMP_TWO[1]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_1, E => un7_delcnt, Q => 
        OP_MODE_c_4_0);
    
    \LOCAL_REG_VAL[0]\ : DFN1E1C0
      port map(D => \SAMP_TWO[0]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_6, E => un7_delcnt, Q => OP_MODE(0));
    
    \LOCAL_REG_VAL[7]\ : DFN1E1C0
      port map(D => \SAMP_TWO[7]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_6, E => un7_delcnt, Q => 
        \LOCAL_REG_VAL[7]_net_1\);
    
    \SYNC_SM_RNO_0[0]\ : OR3
      port map(A => un1_SAMP_TWO_NE_4, B => un1_SAMP_TWO_NE_3, C
         => un1_SAMP_TWO_1, Y => n_sync_sm3);
    
    \DELCNT[0]\ : DFN1C0
      port map(D => \N_DELCNT[0]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_25, Q => \DELCNT[0]_net_1\);
    
    \LOCAL_REG_VAL_2[1]\ : DFN1E1C0
      port map(D => \SAMP_TWO[1]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_1, E => un7_delcnt, Q => 
        OP_MODE_c_2_0);
    
    \LOCAL_REG_VAL[4]\ : DFN1E1C0
      port map(D => \SAMP_TWO[4]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_6, E => un7_delcnt, Q => OP_MODE(4));
    
    \SAMP_ONE[7]\ : DFN1C0
      port map(D => OP_MODE(7), CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c, Q => \SAMP_ONE[7]_net_1\);
    
    \SYNC_SM_RNO_2[0]\ : XO1
      port map(A => \OP_MODE_c[2]\, B => \SAMP_TWO[2]_net_1\, C
         => un1_SAMP_TWO_6, Y => un1_SAMP_TWO_NE_3);
    
    \SAMP_TWO[7]\ : DFN1C0
      port map(D => \SAMP_ONE[7]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_24, Q => \SAMP_TWO[7]_net_1\);
    
    \SAMP_ONE[5]\ : DFN1C0
      port map(D => OP_MODE(5), CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c, Q => \SAMP_ONE[5]_net_1\);
    
    \LOCAL_REG_VAL[6]\ : DFN1E1C0
      port map(D => \SAMP_TWO[6]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_6, E => un7_delcnt, Q => 
        \OP_MODE_c[6]\);
    
    \SYNC_SM_RNO_7[0]\ : XOR2
      port map(A => \SAMP_TWO[6]_net_1\, B => \OP_MODE_c[6]\, Y
         => un1_SAMP_TWO_6);
    
    \SAMP_ONE[6]\ : DFN1C0
      port map(D => OP_MODE(6), CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c, Q => \SAMP_ONE[6]_net_1\);
    
    \SAMP_ONE[0]\ : DFN1C0
      port map(D => OP_MODE_0_0, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c, Q => \SAMP_ONE[0]_net_1\);
    
    \LOCAL_REG_VAL_3[1]\ : DFN1E1C0
      port map(D => \SAMP_TWO[1]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_1, E => un7_delcnt, Q => 
        OP_MODE_c_3_0);
    
    \LOCAL_REG_VAL[1]\ : DFN1E1C0
      port map(D => \SAMP_TWO[1]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_6, E => un7_delcnt, Q => 
        OP_MODE_c_0_d0);
    
    \SAMP_TWO[6]\ : DFN1C0
      port map(D => \SAMP_ONE[6]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_24, Q => \SAMP_TWO[6]_net_1\);
    
    \SAMP_ONE[3]\ : DFN1C0
      port map(D => OP_MODE(3), CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c, Q => \SAMP_ONE[3]_net_1\);
    
    \LOCAL_REG_VAL_0[1]\ : DFN1E1C0
      port map(D => \SAMP_TWO[1]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_1, E => un7_delcnt, Q => 
        OP_MODE_c_0_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity BIDIR_LVTTL is

    port( WR_USB_ADBUS    : in    std_logic_vector(7 downto 0);
          N_RD_USB_ADBUS  : out   std_logic_vector(7 downto 0);
          BIDIR_USB_ADBUS : inout std_logic_vector(7 downto 0) := (others => 'Z');
          TrienAux        : in    std_logic
        );

end BIDIR_LVTTL;

architecture DEF_ARCH of BIDIR_LVTTL is 

  component BIBUF_F_24U
    port( PAD : inout   std_logic;
          D   : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \GND\, \VCC\ : std_logic;

begin 


    \BIBUF_F_24U[6]\ : BIBUF_F_24U
      port map(PAD => BIDIR_USB_ADBUS(6), D => WR_USB_ADBUS(6), E
         => TrienAux, Y => N_RD_USB_ADBUS(6));
    
    \BIBUF_F_24U[7]\ : BIBUF_F_24U
      port map(PAD => BIDIR_USB_ADBUS(7), D => WR_USB_ADBUS(7), E
         => TrienAux, Y => N_RD_USB_ADBUS(7));
    
    \BIBUF_F_24U[4]\ : BIBUF_F_24U
      port map(PAD => BIDIR_USB_ADBUS(4), D => WR_USB_ADBUS(4), E
         => TrienAux, Y => N_RD_USB_ADBUS(4));
    
    \BIBUF_F_24U[2]\ : BIBUF_F_24U
      port map(PAD => BIDIR_USB_ADBUS(2), D => WR_USB_ADBUS(2), E
         => TrienAux, Y => N_RD_USB_ADBUS(2));
    
    \BIBUF_F_24U[1]\ : BIBUF_F_24U
      port map(PAD => BIDIR_USB_ADBUS(1), D => WR_USB_ADBUS(1), E
         => TrienAux, Y => N_RD_USB_ADBUS(1));
    
    \BIBUF_F_24U[3]\ : BIBUF_F_24U
      port map(PAD => BIDIR_USB_ADBUS(3), D => WR_USB_ADBUS(3), E
         => TrienAux, Y => N_RD_USB_ADBUS(3));
    
    \BIBUF_F_24U[0]\ : BIBUF_F_24U
      port map(PAD => BIDIR_USB_ADBUS(0), D => WR_USB_ADBUS(0), E
         => TrienAux, Y => N_RD_USB_ADBUS(0));
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \BIBUF_F_24U[5]\ : BIBUF_F_24U
      port map(PAD => BIDIR_USB_ADBUS(5), D => WR_USB_ADBUS(5), E
         => TrienAux, Y => N_RD_USB_ADBUS(5));
    
    GND_i : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity DPRT_512X9_SRAM_14 is

    port( ELINK_RWA_0         : in    std_logic;
          ELK_RX_SER_WORD_14  : in    std_logic_vector(7 downto 0);
          ELINK_DINA_14       : in    std_logic_vector(7 downto 0);
          ELINK_BLKA_0        : in    std_logic;
          ELKS_ADDRB_0_d0     : in    std_logic;
          ELKS_ADDRB_1        : in    std_logic;
          ELKS_ADDRB_3        : in    std_logic;
          ELKS_ADDRB_5        : in    std_logic;
          ELKS_ADDRB_7        : in    std_logic;
          ELKS_ADDRB_0_0      : in    std_logic;
          ELKS_ADDRB_0_2      : in    std_logic;
          ELKS_ADDRB_0_4      : in    std_logic;
          ELINK_ADDRA_14      : in    std_logic_vector(7 downto 0);
          PATT_ELK_DAT_14     : out   std_logic_vector(7 downto 0);
          ELINK_DOUTA_14      : out   std_logic_vector(7 downto 0);
          ELKS_RWB            : in    std_logic;
          P_USB_MASTER_EN_c_0 : in    std_logic;
          CLK_40M_GL          : in    std_logic;
          CLK60MHZ            : in    std_logic;
          ELKS_RAM_BLKB_EN    : in    std_logic
        );

end DPRT_512X9_SRAM_14;

architecture DEF_ARCH of DPRT_512X9_SRAM_14 is 

  component RAM4K9
    generic (MEMORYFILE:string := "");

    port( ADDRA11 : in    std_logic := 'U';
          ADDRA10 : in    std_logic := 'U';
          ADDRA9  : in    std_logic := 'U';
          ADDRA8  : in    std_logic := 'U';
          ADDRA7  : in    std_logic := 'U';
          ADDRA6  : in    std_logic := 'U';
          ADDRA5  : in    std_logic := 'U';
          ADDRA4  : in    std_logic := 'U';
          ADDRA3  : in    std_logic := 'U';
          ADDRA2  : in    std_logic := 'U';
          ADDRA1  : in    std_logic := 'U';
          ADDRA0  : in    std_logic := 'U';
          ADDRB11 : in    std_logic := 'U';
          ADDRB10 : in    std_logic := 'U';
          ADDRB9  : in    std_logic := 'U';
          ADDRB8  : in    std_logic := 'U';
          ADDRB7  : in    std_logic := 'U';
          ADDRB6  : in    std_logic := 'U';
          ADDRB5  : in    std_logic := 'U';
          ADDRB4  : in    std_logic := 'U';
          ADDRB3  : in    std_logic := 'U';
          ADDRB2  : in    std_logic := 'U';
          ADDRB1  : in    std_logic := 'U';
          ADDRB0  : in    std_logic := 'U';
          DINA8   : in    std_logic := 'U';
          DINA7   : in    std_logic := 'U';
          DINA6   : in    std_logic := 'U';
          DINA5   : in    std_logic := 'U';
          DINA4   : in    std_logic := 'U';
          DINA3   : in    std_logic := 'U';
          DINA2   : in    std_logic := 'U';
          DINA1   : in    std_logic := 'U';
          DINA0   : in    std_logic := 'U';
          DINB8   : in    std_logic := 'U';
          DINB7   : in    std_logic := 'U';
          DINB6   : in    std_logic := 'U';
          DINB5   : in    std_logic := 'U';
          DINB4   : in    std_logic := 'U';
          DINB3   : in    std_logic := 'U';
          DINB2   : in    std_logic := 'U';
          DINB1   : in    std_logic := 'U';
          DINB0   : in    std_logic := 'U';
          WIDTHA0 : in    std_logic := 'U';
          WIDTHA1 : in    std_logic := 'U';
          WIDTHB0 : in    std_logic := 'U';
          WIDTHB1 : in    std_logic := 'U';
          PIPEA   : in    std_logic := 'U';
          PIPEB   : in    std_logic := 'U';
          WMODEA  : in    std_logic := 'U';
          WMODEB  : in    std_logic := 'U';
          BLKA    : in    std_logic := 'U';
          BLKB    : in    std_logic := 'U';
          WENA    : in    std_logic := 'U';
          WENB    : in    std_logic := 'U';
          CLKA    : in    std_logic := 'U';
          CLKB    : in    std_logic := 'U';
          RESET   : in    std_logic := 'U';
          DOUTA8  : out   std_logic;
          DOUTA7  : out   std_logic;
          DOUTA6  : out   std_logic;
          DOUTA5  : out   std_logic;
          DOUTA4  : out   std_logic;
          DOUTA3  : out   std_logic;
          DOUTA2  : out   std_logic;
          DOUTA1  : out   std_logic;
          DOUTA0  : out   std_logic;
          DOUTB8  : out   std_logic;
          DOUTB7  : out   std_logic;
          DOUTB6  : out   std_logic;
          DOUTB5  : out   std_logic;
          DOUTB4  : out   std_logic;
          DOUTB3  : out   std_logic;
          DOUTB2  : out   std_logic;
          DOUTB1  : out   std_logic;
          DOUTB0  : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \DOUTA_1[8]\, \DOUTB_1[8]\, DPRT_512X9_SRAM_14_GND, 
        DPRT_512X9_SRAM_14_VCC : std_logic;

begin 


    DPRT_512X9_SRAM_R0C0 : RAM4K9
      generic map(MEMORYFILE => "DPRT_512X9_SRAM_R0C0.mem")

      port map(ADDRA11 => DPRT_512X9_SRAM_14_GND, ADDRA10 => 
        DPRT_512X9_SRAM_14_GND, ADDRA9 => DPRT_512X9_SRAM_14_GND, 
        ADDRA8 => DPRT_512X9_SRAM_14_GND, ADDRA7 => 
        ELINK_ADDRA_14(7), ADDRA6 => ELINK_ADDRA_14(6), ADDRA5
         => ELINK_ADDRA_14(5), ADDRA4 => ELINK_ADDRA_14(4), 
        ADDRA3 => ELINK_ADDRA_14(3), ADDRA2 => ELINK_ADDRA_14(2), 
        ADDRA1 => ELINK_ADDRA_14(1), ADDRA0 => ELINK_ADDRA_14(0), 
        ADDRB11 => DPRT_512X9_SRAM_14_GND, ADDRB10 => 
        DPRT_512X9_SRAM_14_GND, ADDRB9 => DPRT_512X9_SRAM_14_GND, 
        ADDRB8 => DPRT_512X9_SRAM_14_GND, ADDRB7 => ELKS_ADDRB_7, 
        ADDRB6 => ELKS_ADDRB_0_4, ADDRB5 => ELKS_ADDRB_5, ADDRB4
         => ELKS_ADDRB_0_2, ADDRB3 => ELKS_ADDRB_3, ADDRB2 => 
        ELKS_ADDRB_0_0, ADDRB1 => ELKS_ADDRB_1, ADDRB0 => 
        ELKS_ADDRB_0_d0, DINA8 => DPRT_512X9_SRAM_14_GND, DINA7
         => ELINK_DINA_14(7), DINA6 => ELINK_DINA_14(6), DINA5
         => ELINK_DINA_14(5), DINA4 => ELINK_DINA_14(4), DINA3
         => ELINK_DINA_14(3), DINA2 => ELINK_DINA_14(2), DINA1
         => ELINK_DINA_14(1), DINA0 => ELINK_DINA_14(0), DINB8
         => DPRT_512X9_SRAM_14_GND, DINB7 => 
        ELK_RX_SER_WORD_14(7), DINB6 => ELK_RX_SER_WORD_14(6), 
        DINB5 => ELK_RX_SER_WORD_14(5), DINB4 => 
        ELK_RX_SER_WORD_14(4), DINB3 => ELK_RX_SER_WORD_14(3), 
        DINB2 => ELK_RX_SER_WORD_14(2), DINB1 => 
        ELK_RX_SER_WORD_14(1), DINB0 => ELK_RX_SER_WORD_14(0), 
        WIDTHA0 => DPRT_512X9_SRAM_14_VCC, WIDTHA1 => 
        DPRT_512X9_SRAM_14_VCC, WIDTHB0 => DPRT_512X9_SRAM_14_VCC, 
        WIDTHB1 => DPRT_512X9_SRAM_14_VCC, PIPEA => 
        DPRT_512X9_SRAM_14_VCC, PIPEB => DPRT_512X9_SRAM_14_VCC, 
        WMODEA => DPRT_512X9_SRAM_14_GND, WMODEB => 
        DPRT_512X9_SRAM_14_GND, BLKA => ELINK_BLKA_0, BLKB => 
        ELKS_RAM_BLKB_EN, WENA => ELINK_RWA_0, WENB => ELKS_RWB, 
        CLKA => CLK60MHZ, CLKB => CLK_40M_GL, RESET => 
        P_USB_MASTER_EN_c_0, DOUTA8 => \DOUTA_1[8]\, DOUTA7 => 
        ELINK_DOUTA_14(7), DOUTA6 => ELINK_DOUTA_14(6), DOUTA5
         => ELINK_DOUTA_14(5), DOUTA4 => ELINK_DOUTA_14(4), 
        DOUTA3 => ELINK_DOUTA_14(3), DOUTA2 => ELINK_DOUTA_14(2), 
        DOUTA1 => ELINK_DOUTA_14(1), DOUTA0 => ELINK_DOUTA_14(0), 
        DOUTB8 => \DOUTB_1[8]\, DOUTB7 => PATT_ELK_DAT_14(7), 
        DOUTB6 => PATT_ELK_DAT_14(6), DOUTB5 => 
        PATT_ELK_DAT_14(5), DOUTB4 => PATT_ELK_DAT_14(4), DOUTB3
         => PATT_ELK_DAT_14(3), DOUTB2 => PATT_ELK_DAT_14(2), 
        DOUTB1 => PATT_ELK_DAT_14(1), DOUTB0 => 
        PATT_ELK_DAT_14(0));
    
    VCC_i : VCC
      port map(Y => DPRT_512X9_SRAM_14_VCC);
    
    GND_i : GND
      port map(Y => DPRT_512X9_SRAM_14_GND);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity DPRT_512X9_SRAM_17 is

    port( ELINK_RWA_0         : in    std_logic;
          ELK_RX_SER_WORD_17  : in    std_logic_vector(7 downto 0);
          ELINK_DINA_17       : in    std_logic_vector(7 downto 0);
          ELINK_BLKA_0        : in    std_logic;
          ELKS_ADDRB          : in    std_logic_vector(7 downto 0);
          ELINK_ADDRA_17      : in    std_logic_vector(7 downto 0);
          PATT_ELK_DAT_17     : out   std_logic_vector(7 downto 0);
          ELINK_DOUTA_17      : out   std_logic_vector(7 downto 0);
          ELKS_RWB            : in    std_logic;
          P_USB_MASTER_EN_c_0 : in    std_logic;
          CLK_40M_GL          : in    std_logic;
          CLK60MHZ            : in    std_logic;
          ELKS_RAM_BLKB_EN    : in    std_logic
        );

end DPRT_512X9_SRAM_17;

architecture DEF_ARCH of DPRT_512X9_SRAM_17 is 

  component RAM4K9
    generic (MEMORYFILE:string := "");

    port( ADDRA11 : in    std_logic := 'U';
          ADDRA10 : in    std_logic := 'U';
          ADDRA9  : in    std_logic := 'U';
          ADDRA8  : in    std_logic := 'U';
          ADDRA7  : in    std_logic := 'U';
          ADDRA6  : in    std_logic := 'U';
          ADDRA5  : in    std_logic := 'U';
          ADDRA4  : in    std_logic := 'U';
          ADDRA3  : in    std_logic := 'U';
          ADDRA2  : in    std_logic := 'U';
          ADDRA1  : in    std_logic := 'U';
          ADDRA0  : in    std_logic := 'U';
          ADDRB11 : in    std_logic := 'U';
          ADDRB10 : in    std_logic := 'U';
          ADDRB9  : in    std_logic := 'U';
          ADDRB8  : in    std_logic := 'U';
          ADDRB7  : in    std_logic := 'U';
          ADDRB6  : in    std_logic := 'U';
          ADDRB5  : in    std_logic := 'U';
          ADDRB4  : in    std_logic := 'U';
          ADDRB3  : in    std_logic := 'U';
          ADDRB2  : in    std_logic := 'U';
          ADDRB1  : in    std_logic := 'U';
          ADDRB0  : in    std_logic := 'U';
          DINA8   : in    std_logic := 'U';
          DINA7   : in    std_logic := 'U';
          DINA6   : in    std_logic := 'U';
          DINA5   : in    std_logic := 'U';
          DINA4   : in    std_logic := 'U';
          DINA3   : in    std_logic := 'U';
          DINA2   : in    std_logic := 'U';
          DINA1   : in    std_logic := 'U';
          DINA0   : in    std_logic := 'U';
          DINB8   : in    std_logic := 'U';
          DINB7   : in    std_logic := 'U';
          DINB6   : in    std_logic := 'U';
          DINB5   : in    std_logic := 'U';
          DINB4   : in    std_logic := 'U';
          DINB3   : in    std_logic := 'U';
          DINB2   : in    std_logic := 'U';
          DINB1   : in    std_logic := 'U';
          DINB0   : in    std_logic := 'U';
          WIDTHA0 : in    std_logic := 'U';
          WIDTHA1 : in    std_logic := 'U';
          WIDTHB0 : in    std_logic := 'U';
          WIDTHB1 : in    std_logic := 'U';
          PIPEA   : in    std_logic := 'U';
          PIPEB   : in    std_logic := 'U';
          WMODEA  : in    std_logic := 'U';
          WMODEB  : in    std_logic := 'U';
          BLKA    : in    std_logic := 'U';
          BLKB    : in    std_logic := 'U';
          WENA    : in    std_logic := 'U';
          WENB    : in    std_logic := 'U';
          CLKA    : in    std_logic := 'U';
          CLKB    : in    std_logic := 'U';
          RESET   : in    std_logic := 'U';
          DOUTA8  : out   std_logic;
          DOUTA7  : out   std_logic;
          DOUTA6  : out   std_logic;
          DOUTA5  : out   std_logic;
          DOUTA4  : out   std_logic;
          DOUTA3  : out   std_logic;
          DOUTA2  : out   std_logic;
          DOUTA1  : out   std_logic;
          DOUTA0  : out   std_logic;
          DOUTB8  : out   std_logic;
          DOUTB7  : out   std_logic;
          DOUTB6  : out   std_logic;
          DOUTB5  : out   std_logic;
          DOUTB4  : out   std_logic;
          DOUTB3  : out   std_logic;
          DOUTB2  : out   std_logic;
          DOUTB1  : out   std_logic;
          DOUTB0  : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \DOUTA_1[8]\, \DOUTB_1[8]\, DPRT_512X9_SRAM_17_GND, 
        DPRT_512X9_SRAM_17_VCC : std_logic;

begin 


    DPRT_512X9_SRAM_R0C0 : RAM4K9
      generic map(MEMORYFILE => "DPRT_512X9_SRAM_R0C0.mem")

      port map(ADDRA11 => DPRT_512X9_SRAM_17_GND, ADDRA10 => 
        DPRT_512X9_SRAM_17_GND, ADDRA9 => DPRT_512X9_SRAM_17_GND, 
        ADDRA8 => DPRT_512X9_SRAM_17_GND, ADDRA7 => 
        ELINK_ADDRA_17(7), ADDRA6 => ELINK_ADDRA_17(6), ADDRA5
         => ELINK_ADDRA_17(5), ADDRA4 => ELINK_ADDRA_17(4), 
        ADDRA3 => ELINK_ADDRA_17(3), ADDRA2 => ELINK_ADDRA_17(2), 
        ADDRA1 => ELINK_ADDRA_17(1), ADDRA0 => ELINK_ADDRA_17(0), 
        ADDRB11 => DPRT_512X9_SRAM_17_GND, ADDRB10 => 
        DPRT_512X9_SRAM_17_GND, ADDRB9 => DPRT_512X9_SRAM_17_GND, 
        ADDRB8 => DPRT_512X9_SRAM_17_GND, ADDRB7 => ELKS_ADDRB(7), 
        ADDRB6 => ELKS_ADDRB(6), ADDRB5 => ELKS_ADDRB(5), ADDRB4
         => ELKS_ADDRB(4), ADDRB3 => ELKS_ADDRB(3), ADDRB2 => 
        ELKS_ADDRB(2), ADDRB1 => ELKS_ADDRB(1), ADDRB0 => 
        ELKS_ADDRB(0), DINA8 => DPRT_512X9_SRAM_17_GND, DINA7 => 
        ELINK_DINA_17(7), DINA6 => ELINK_DINA_17(6), DINA5 => 
        ELINK_DINA_17(5), DINA4 => ELINK_DINA_17(4), DINA3 => 
        ELINK_DINA_17(3), DINA2 => ELINK_DINA_17(2), DINA1 => 
        ELINK_DINA_17(1), DINA0 => ELINK_DINA_17(0), DINB8 => 
        DPRT_512X9_SRAM_17_GND, DINB7 => ELK_RX_SER_WORD_17(7), 
        DINB6 => ELK_RX_SER_WORD_17(6), DINB5 => 
        ELK_RX_SER_WORD_17(5), DINB4 => ELK_RX_SER_WORD_17(4), 
        DINB3 => ELK_RX_SER_WORD_17(3), DINB2 => 
        ELK_RX_SER_WORD_17(2), DINB1 => ELK_RX_SER_WORD_17(1), 
        DINB0 => ELK_RX_SER_WORD_17(0), WIDTHA0 => 
        DPRT_512X9_SRAM_17_VCC, WIDTHA1 => DPRT_512X9_SRAM_17_VCC, 
        WIDTHB0 => DPRT_512X9_SRAM_17_VCC, WIDTHB1 => 
        DPRT_512X9_SRAM_17_VCC, PIPEA => DPRT_512X9_SRAM_17_VCC, 
        PIPEB => DPRT_512X9_SRAM_17_VCC, WMODEA => 
        DPRT_512X9_SRAM_17_GND, WMODEB => DPRT_512X9_SRAM_17_GND, 
        BLKA => ELINK_BLKA_0, BLKB => ELKS_RAM_BLKB_EN, WENA => 
        ELINK_RWA_0, WENB => ELKS_RWB, CLKA => CLK60MHZ, CLKB => 
        CLK_40M_GL, RESET => P_USB_MASTER_EN_c_0, DOUTA8 => 
        \DOUTA_1[8]\, DOUTA7 => ELINK_DOUTA_17(7), DOUTA6 => 
        ELINK_DOUTA_17(6), DOUTA5 => ELINK_DOUTA_17(5), DOUTA4
         => ELINK_DOUTA_17(4), DOUTA3 => ELINK_DOUTA_17(3), 
        DOUTA2 => ELINK_DOUTA_17(2), DOUTA1 => ELINK_DOUTA_17(1), 
        DOUTA0 => ELINK_DOUTA_17(0), DOUTB8 => \DOUTB_1[8]\, 
        DOUTB7 => PATT_ELK_DAT_17(7), DOUTB6 => 
        PATT_ELK_DAT_17(6), DOUTB5 => PATT_ELK_DAT_17(5), DOUTB4
         => PATT_ELK_DAT_17(4), DOUTB3 => PATT_ELK_DAT_17(3), 
        DOUTB2 => PATT_ELK_DAT_17(2), DOUTB1 => 
        PATT_ELK_DAT_17(1), DOUTB0 => PATT_ELK_DAT_17(0));
    
    VCC_i : VCC
      port map(Y => DPRT_512X9_SRAM_17_VCC);
    
    GND_i : GND
      port map(Y => DPRT_512X9_SRAM_17_GND);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity CLK60M_TO_40M_4_2 is

    port( ELINKS_STOP_ADDR    : in    std_logic_vector(7 downto 0);
          ELKS_STOP_ADDR      : out   std_logic_vector(7 downto 0);
          P_MASTER_POR_B_c_26 : in    std_logic;
          P_MASTER_POR_B_c_30 : in    std_logic;
          P_MASTER_POR_B_c_3  : in    std_logic;
          P_MASTER_POR_B_c_25 : in    std_logic;
          CLK_40M_GL          : in    std_logic
        );

end CLK60M_TO_40M_4_2;

architecture DEF_ARCH of CLK60M_TO_40M_4_2 is 

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component XO1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component MX2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal un1_SAMP_TWO_NE_4, un1_SAMP_TWO_5, un1_SAMP_TWO_4, 
        un1_SAMP_TWO_NE_1, un1_SAMP_TWO_NE_3, \ELKS_STOP_ADDR[2]\, 
        \SAMP_TWO[2]_net_1\, un1_SAMP_TWO_3, un1_SAMP_TWO_NE_2, 
        \ELKS_STOP_ADDR[0]\, \SAMP_TWO[0]_net_1\, un1_SAMP_TWO_1, 
        \ELKS_STOP_ADDR[6]\, \SAMP_TWO[6]_net_1\, un1_SAMP_TWO_7, 
        n_sync_sm3, \N_DELCNT[0]\, \SYNC_SM[0]_net_1\, 
        \DELCNT[0]_net_1\, un7_delcnt, \DELCNT[1]_net_1\, 
        \N_SYNC_SM[0]\, \SAMP_TWO[7]_net_1\, \ELKS_STOP_ADDR[7]\, 
        \SAMP_TWO[5]_net_1\, \ELKS_STOP_ADDR[5]\, 
        \SAMP_TWO[4]_net_1\, \ELKS_STOP_ADDR[4]\, 
        \SAMP_TWO[3]_net_1\, \ELKS_STOP_ADDR[3]\, 
        \SAMP_TWO[1]_net_1\, \ELKS_STOP_ADDR[1]\, SUM1_3, 
        \SAMP_ONE[0]_net_1\, \SAMP_ONE[1]_net_1\, 
        \SAMP_ONE[2]_net_1\, \SAMP_ONE[3]_net_1\, 
        \SAMP_ONE[4]_net_1\, \SAMP_ONE[5]_net_1\, 
        \SAMP_ONE[6]_net_1\, \SAMP_ONE[7]_net_1\, \GND\, \VCC\
         : std_logic;

begin 

    ELKS_STOP_ADDR(7) <= \ELKS_STOP_ADDR[7]\;
    ELKS_STOP_ADDR(6) <= \ELKS_STOP_ADDR[6]\;
    ELKS_STOP_ADDR(5) <= \ELKS_STOP_ADDR[5]\;
    ELKS_STOP_ADDR(4) <= \ELKS_STOP_ADDR[4]\;
    ELKS_STOP_ADDR(3) <= \ELKS_STOP_ADDR[3]\;
    ELKS_STOP_ADDR(2) <= \ELKS_STOP_ADDR[2]\;
    ELKS_STOP_ADDR(1) <= \ELKS_STOP_ADDR[1]\;
    ELKS_STOP_ADDR(0) <= \ELKS_STOP_ADDR[0]\;

    \SAMP_ONE[2]\ : DFN1C0
      port map(D => ELINKS_STOP_ADDR(2), CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_25, Q => \SAMP_ONE[2]_net_1\);
    
    \SYNC_SM_RNO_6[0]\ : XOR2
      port map(A => \SAMP_TWO[5]_net_1\, B => \ELKS_STOP_ADDR[5]\, 
        Y => un1_SAMP_TWO_5);
    
    \LOCAL_REG_VAL[3]\ : DFN1E1C0
      port map(D => \SAMP_TWO[3]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_3, E => un7_delcnt, Q => 
        \ELKS_STOP_ADDR[3]\);
    
    \DELCNT_RNIPSMD[1]\ : NOR2B
      port map(A => \DELCNT[1]_net_1\, B => \DELCNT[0]_net_1\, Y
         => un7_delcnt);
    
    \SYNC_SM[0]\ : DFN1C0
      port map(D => \N_SYNC_SM[0]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_25, Q => \SYNC_SM[0]_net_1\);
    
    \SYNC_SM_RNO_5[0]\ : XOR2
      port map(A => \SAMP_TWO[1]_net_1\, B => \ELKS_STOP_ADDR[1]\, 
        Y => un1_SAMP_TWO_1);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \DELCNT[1]\ : DFN1C0
      port map(D => SUM1_3, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_26, Q => \DELCNT[1]_net_1\);
    
    \LOCAL_REG_VAL[5]\ : DFN1E1C0
      port map(D => \SAMP_TWO[5]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_3, E => un7_delcnt, Q => 
        \ELKS_STOP_ADDR[5]\);
    
    \SYNC_SM_RNO_1[0]\ : XO1
      port map(A => \ELKS_STOP_ADDR[2]\, B => \SAMP_TWO[2]_net_1\, 
        C => un1_SAMP_TWO_3, Y => un1_SAMP_TWO_NE_3);
    
    \SAMP_TWO[0]\ : DFN1C0
      port map(D => \SAMP_ONE[0]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_30, Q => \SAMP_TWO[0]_net_1\);
    
    \SAMP_ONE[1]\ : DFN1C0
      port map(D => ELINKS_STOP_ADDR(1), CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_25, Q => \SAMP_ONE[1]_net_1\);
    
    \SAMP_TWO[1]\ : DFN1C0
      port map(D => \SAMP_ONE[1]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_30, Q => \SAMP_TWO[1]_net_1\);
    
    \SYNC_SM_RNO_3[0]\ : OR3
      port map(A => un1_SAMP_TWO_5, B => un1_SAMP_TWO_4, C => 
        un1_SAMP_TWO_NE_1, Y => un1_SAMP_TWO_NE_4);
    
    \SYNC_SM_RNO_9[0]\ : XOR2
      port map(A => \SAMP_TWO[7]_net_1\, B => \ELKS_STOP_ADDR[7]\, 
        Y => un1_SAMP_TWO_7);
    
    un2_n_delcnt_1_1_SUM1 : XOR2
      port map(A => \DELCNT[1]_net_1\, B => \DELCNT[0]_net_1\, Y
         => SUM1_3);
    
    \SAMP_TWO[3]\ : DFN1C0
      port map(D => \SAMP_ONE[3]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_30, Q => \SAMP_TWO[3]_net_1\);
    
    \SYNC_SM_RNO_8[0]\ : XO1
      port map(A => \ELKS_STOP_ADDR[6]\, B => \SAMP_TWO[6]_net_1\, 
        C => un1_SAMP_TWO_7, Y => un1_SAMP_TWO_NE_1);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \SYNC_SM_RNO_4[0]\ : XOR2
      port map(A => \SAMP_TWO[3]_net_1\, B => \ELKS_STOP_ADDR[3]\, 
        Y => un1_SAMP_TWO_3);
    
    \SYNC_SM_RNO[0]\ : MX2B
      port map(A => n_sync_sm3, B => un7_delcnt, S => 
        \SYNC_SM[0]_net_1\, Y => \N_SYNC_SM[0]\);
    
    \SAMP_ONE[4]\ : DFN1C0
      port map(D => ELINKS_STOP_ADDR(4), CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_25, Q => \SAMP_ONE[4]_net_1\);
    
    \LOCAL_REG_VAL[2]\ : DFN1E1C0
      port map(D => \SAMP_TWO[2]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_3, E => un7_delcnt, Q => 
        \ELKS_STOP_ADDR[2]\);
    
    \SAMP_TWO[5]\ : DFN1C0
      port map(D => \SAMP_ONE[5]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_30, Q => \SAMP_TWO[5]_net_1\);
    
    \SAMP_TWO[4]\ : DFN1C0
      port map(D => \SAMP_ONE[4]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_30, Q => \SAMP_TWO[4]_net_1\);
    
    \SAMP_TWO[2]\ : DFN1C0
      port map(D => \SAMP_ONE[2]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_30, Q => \SAMP_TWO[2]_net_1\);
    
    \DELCNT_RNO[0]\ : NOR2A
      port map(A => \SYNC_SM[0]_net_1\, B => \DELCNT[0]_net_1\, Y
         => \N_DELCNT[0]\);
    
    \LOCAL_REG_VAL[0]\ : DFN1E1C0
      port map(D => \SAMP_TWO[0]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_3, E => un7_delcnt, Q => 
        \ELKS_STOP_ADDR[0]\);
    
    \LOCAL_REG_VAL[7]\ : DFN1E1C0
      port map(D => \SAMP_TWO[7]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_3, E => un7_delcnt, Q => 
        \ELKS_STOP_ADDR[7]\);
    
    \SYNC_SM_RNO_0[0]\ : OR3
      port map(A => un1_SAMP_TWO_NE_3, B => un1_SAMP_TWO_NE_2, C
         => un1_SAMP_TWO_NE_4, Y => n_sync_sm3);
    
    \DELCNT[0]\ : DFN1C0
      port map(D => \N_DELCNT[0]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_26, Q => \DELCNT[0]_net_1\);
    
    \LOCAL_REG_VAL[4]\ : DFN1E1C0
      port map(D => \SAMP_TWO[4]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_3, E => un7_delcnt, Q => 
        \ELKS_STOP_ADDR[4]\);
    
    \SAMP_ONE[7]\ : DFN1C0
      port map(D => ELINKS_STOP_ADDR(7), CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_25, Q => \SAMP_ONE[7]_net_1\);
    
    \SYNC_SM_RNO_2[0]\ : XO1
      port map(A => \ELKS_STOP_ADDR[0]\, B => \SAMP_TWO[0]_net_1\, 
        C => un1_SAMP_TWO_1, Y => un1_SAMP_TWO_NE_2);
    
    \SAMP_TWO[7]\ : DFN1C0
      port map(D => \SAMP_ONE[7]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_30, Q => \SAMP_TWO[7]_net_1\);
    
    \SAMP_ONE[5]\ : DFN1C0
      port map(D => ELINKS_STOP_ADDR(5), CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_25, Q => \SAMP_ONE[5]_net_1\);
    
    \LOCAL_REG_VAL[6]\ : DFN1E1C0
      port map(D => \SAMP_TWO[6]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_3, E => un7_delcnt, Q => 
        \ELKS_STOP_ADDR[6]\);
    
    \SYNC_SM_RNO_7[0]\ : XOR2
      port map(A => \SAMP_TWO[4]_net_1\, B => \ELKS_STOP_ADDR[4]\, 
        Y => un1_SAMP_TWO_4);
    
    \SAMP_ONE[6]\ : DFN1C0
      port map(D => ELINKS_STOP_ADDR(6), CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_25, Q => \SAMP_ONE[6]_net_1\);
    
    \SAMP_ONE[0]\ : DFN1C0
      port map(D => ELINKS_STOP_ADDR(0), CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_25, Q => \SAMP_ONE[0]_net_1\);
    
    \LOCAL_REG_VAL[1]\ : DFN1E1C0
      port map(D => \SAMP_TWO[1]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_3, E => un7_delcnt, Q => 
        \ELKS_STOP_ADDR[1]\);
    
    \SAMP_TWO[6]\ : DFN1C0
      port map(D => \SAMP_ONE[6]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_30, Q => \SAMP_TWO[6]_net_1\);
    
    \SAMP_ONE[3]\ : DFN1C0
      port map(D => ELINKS_STOP_ADDR(3), CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_25, Q => \SAMP_ONE[3]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity CLK60M_TO_40M_4_0 is

    port( TFC_STOP_ADDR_0       : in    std_logic_vector(7 downto 0);
          TFC_STOP_ADDR         : out   std_logic_vector(7 downto 0);
          P_MASTER_POR_B_c_30   : in    std_logic;
          P_MASTER_POR_B_c_29   : in    std_logic;
          P_MASTER_POR_B_c_25   : in    std_logic;
          P_MASTER_POR_B_c_24_0 : in    std_logic;
          P_MASTER_POR_B_c_19   : in    std_logic;
          P_MASTER_POR_B_c_23   : in    std_logic;
          CLK_40M_GL            : in    std_logic
        );

end CLK60M_TO_40M_4_0;

architecture DEF_ARCH of CLK60M_TO_40M_4_0 is 

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component XO1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component MX2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal un1_SAMP_TWO_NE_4, un1_SAMP_TWO_5, un1_SAMP_TWO_4, 
        un1_SAMP_TWO_NE_1, un1_SAMP_TWO_NE_3, \TFC_STOP_ADDR[2]\, 
        \SAMP_TWO[2]_net_1\, un1_SAMP_TWO_3, un1_SAMP_TWO_NE_2, 
        \TFC_STOP_ADDR[0]\, \SAMP_TWO[0]_net_1\, un1_SAMP_TWO_1, 
        \TFC_STOP_ADDR[6]\, \SAMP_TWO[6]_net_1\, un1_SAMP_TWO_7, 
        n_sync_sm3, \N_DELCNT[0]\, \SYNC_SM[0]_net_1\, 
        \DELCNT[0]_net_1\, un7_delcnt, \DELCNT[1]_net_1\, 
        \N_SYNC_SM[0]\, \SAMP_TWO[7]_net_1\, \TFC_STOP_ADDR[7]\, 
        \SAMP_TWO[5]_net_1\, \TFC_STOP_ADDR[5]\, 
        \SAMP_TWO[4]_net_1\, \TFC_STOP_ADDR[4]\, 
        \SAMP_TWO[3]_net_1\, \TFC_STOP_ADDR[3]\, 
        \SAMP_TWO[1]_net_1\, \TFC_STOP_ADDR[1]\, SUM1_1, 
        \SAMP_ONE[0]_net_1\, \SAMP_ONE[1]_net_1\, 
        \SAMP_ONE[2]_net_1\, \SAMP_ONE[3]_net_1\, 
        \SAMP_ONE[4]_net_1\, \SAMP_ONE[5]_net_1\, 
        \SAMP_ONE[6]_net_1\, \SAMP_ONE[7]_net_1\, \GND\, \VCC\
         : std_logic;

begin 

    TFC_STOP_ADDR(7) <= \TFC_STOP_ADDR[7]\;
    TFC_STOP_ADDR(6) <= \TFC_STOP_ADDR[6]\;
    TFC_STOP_ADDR(5) <= \TFC_STOP_ADDR[5]\;
    TFC_STOP_ADDR(4) <= \TFC_STOP_ADDR[4]\;
    TFC_STOP_ADDR(3) <= \TFC_STOP_ADDR[3]\;
    TFC_STOP_ADDR(2) <= \TFC_STOP_ADDR[2]\;
    TFC_STOP_ADDR(1) <= \TFC_STOP_ADDR[1]\;
    TFC_STOP_ADDR(0) <= \TFC_STOP_ADDR[0]\;

    \SAMP_ONE[2]\ : DFN1C0
      port map(D => TFC_STOP_ADDR_0(2), CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_25, Q => \SAMP_ONE[2]_net_1\);
    
    \SYNC_SM_RNO_6[0]\ : XOR2
      port map(A => \SAMP_TWO[5]_net_1\, B => \TFC_STOP_ADDR[5]\, 
        Y => un1_SAMP_TWO_5);
    
    \LOCAL_REG_VAL[3]\ : DFN1E1C0
      port map(D => \SAMP_TWO[3]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_19, E => un7_delcnt, Q => 
        \TFC_STOP_ADDR[3]\);
    
    \SYNC_SM[0]\ : DFN1C0
      port map(D => \N_SYNC_SM[0]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_23, Q => \SYNC_SM[0]_net_1\);
    
    \SYNC_SM_RNO_5[0]\ : XOR2
      port map(A => \SAMP_TWO[1]_net_1\, B => \TFC_STOP_ADDR[1]\, 
        Y => un1_SAMP_TWO_1);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \DELCNT[1]\ : DFN1C0
      port map(D => SUM1_1, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_30, Q => \DELCNT[1]_net_1\);
    
    \LOCAL_REG_VAL[5]\ : DFN1E1C0
      port map(D => \SAMP_TWO[5]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_19, E => un7_delcnt, Q => 
        \TFC_STOP_ADDR[5]\);
    
    \SYNC_SM_RNO_1[0]\ : XO1
      port map(A => \TFC_STOP_ADDR[2]\, B => \SAMP_TWO[2]_net_1\, 
        C => un1_SAMP_TWO_3, Y => un1_SAMP_TWO_NE_3);
    
    \SAMP_TWO[0]\ : DFN1C0
      port map(D => \SAMP_ONE[0]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_29, Q => \SAMP_TWO[0]_net_1\);
    
    \SAMP_ONE[1]\ : DFN1C0
      port map(D => TFC_STOP_ADDR_0(1), CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_24_0, Q => \SAMP_ONE[1]_net_1\);
    
    \SAMP_TWO[1]\ : DFN1C0
      port map(D => \SAMP_ONE[1]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_29, Q => \SAMP_TWO[1]_net_1\);
    
    \SYNC_SM_RNO_3[0]\ : OR3
      port map(A => un1_SAMP_TWO_5, B => un1_SAMP_TWO_4, C => 
        un1_SAMP_TWO_NE_1, Y => un1_SAMP_TWO_NE_4);
    
    \SYNC_SM_RNO_9[0]\ : XOR2
      port map(A => \SAMP_TWO[7]_net_1\, B => \TFC_STOP_ADDR[7]\, 
        Y => un1_SAMP_TWO_7);
    
    un2_n_delcnt_1_1_SUM1 : XOR2
      port map(A => \DELCNT[1]_net_1\, B => \DELCNT[0]_net_1\, Y
         => SUM1_1);
    
    \SAMP_TWO[3]\ : DFN1C0
      port map(D => \SAMP_ONE[3]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_29, Q => \SAMP_TWO[3]_net_1\);
    
    \SYNC_SM_RNO_8[0]\ : XO1
      port map(A => \TFC_STOP_ADDR[6]\, B => \SAMP_TWO[6]_net_1\, 
        C => un1_SAMP_TWO_7, Y => un1_SAMP_TWO_NE_1);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \SYNC_SM_RNO_4[0]\ : XOR2
      port map(A => \SAMP_TWO[3]_net_1\, B => \TFC_STOP_ADDR[3]\, 
        Y => un1_SAMP_TWO_3);
    
    \SYNC_SM_RNO[0]\ : MX2B
      port map(A => n_sync_sm3, B => un7_delcnt, S => 
        \SYNC_SM[0]_net_1\, Y => \N_SYNC_SM[0]\);
    
    \SAMP_ONE[4]\ : DFN1C0
      port map(D => TFC_STOP_ADDR_0(4), CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_25, Q => \SAMP_ONE[4]_net_1\);
    
    \LOCAL_REG_VAL[2]\ : DFN1E1C0
      port map(D => \SAMP_TWO[2]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_19, E => un7_delcnt, Q => 
        \TFC_STOP_ADDR[2]\);
    
    \SAMP_TWO[5]\ : DFN1C0
      port map(D => \SAMP_ONE[5]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_29, Q => \SAMP_TWO[5]_net_1\);
    
    \SAMP_TWO[4]\ : DFN1C0
      port map(D => \SAMP_ONE[4]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_29, Q => \SAMP_TWO[4]_net_1\);
    
    \SAMP_TWO[2]\ : DFN1C0
      port map(D => \SAMP_ONE[2]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_29, Q => \SAMP_TWO[2]_net_1\);
    
    \DELCNT_RNO[0]\ : NOR2A
      port map(A => \SYNC_SM[0]_net_1\, B => \DELCNT[0]_net_1\, Y
         => \N_DELCNT[0]\);
    
    \LOCAL_REG_VAL[0]\ : DFN1E1C0
      port map(D => \SAMP_TWO[0]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_19, E => un7_delcnt, Q => 
        \TFC_STOP_ADDR[0]\);
    
    \LOCAL_REG_VAL[7]\ : DFN1E1C0
      port map(D => \SAMP_TWO[7]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_19, E => un7_delcnt, Q => 
        \TFC_STOP_ADDR[7]\);
    
    \SYNC_SM_RNO_0[0]\ : OR3
      port map(A => un1_SAMP_TWO_NE_3, B => un1_SAMP_TWO_NE_2, C
         => un1_SAMP_TWO_NE_4, Y => n_sync_sm3);
    
    \DELCNT[0]\ : DFN1C0
      port map(D => \N_DELCNT[0]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_30, Q => \DELCNT[0]_net_1\);
    
    \LOCAL_REG_VAL[4]\ : DFN1E1C0
      port map(D => \SAMP_TWO[4]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_19, E => un7_delcnt, Q => 
        \TFC_STOP_ADDR[4]\);
    
    \SAMP_ONE[7]\ : DFN1C0
      port map(D => TFC_STOP_ADDR_0(7), CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_25, Q => \SAMP_ONE[7]_net_1\);
    
    \SYNC_SM_RNO_2[0]\ : XO1
      port map(A => \TFC_STOP_ADDR[0]\, B => \SAMP_TWO[0]_net_1\, 
        C => un1_SAMP_TWO_1, Y => un1_SAMP_TWO_NE_2);
    
    \SAMP_TWO[7]\ : DFN1C0
      port map(D => \SAMP_ONE[7]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_29, Q => \SAMP_TWO[7]_net_1\);
    
    \SAMP_ONE[5]\ : DFN1C0
      port map(D => TFC_STOP_ADDR_0(5), CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_25, Q => \SAMP_ONE[5]_net_1\);
    
    \LOCAL_REG_VAL[6]\ : DFN1E1C0
      port map(D => \SAMP_TWO[6]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_19, E => un7_delcnt, Q => 
        \TFC_STOP_ADDR[6]\);
    
    \SYNC_SM_RNO_7[0]\ : XOR2
      port map(A => \SAMP_TWO[4]_net_1\, B => \TFC_STOP_ADDR[4]\, 
        Y => un1_SAMP_TWO_4);
    
    \SAMP_ONE[6]\ : DFN1C0
      port map(D => TFC_STOP_ADDR_0(6), CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_25, Q => \SAMP_ONE[6]_net_1\);
    
    \SAMP_ONE[0]\ : DFN1C0
      port map(D => TFC_STOP_ADDR_0(0), CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_24_0, Q => \SAMP_ONE[0]_net_1\);
    
    \LOCAL_REG_VAL[1]\ : DFN1E1C0
      port map(D => \SAMP_TWO[1]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_19, E => un7_delcnt, Q => 
        \TFC_STOP_ADDR[1]\);
    
    \SAMP_TWO[6]\ : DFN1C0
      port map(D => \SAMP_ONE[6]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_29, Q => \SAMP_TWO[6]_net_1\);
    
    \SAMP_ONE[3]\ : DFN1C0
      port map(D => TFC_STOP_ADDR_0(3), CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_25, Q => \SAMP_ONE[3]_net_1\);
    
    \DELCNT_RNILG8K[1]\ : NOR2B
      port map(A => \DELCNT[1]_net_1\, B => \DELCNT[0]_net_1\, Y
         => un7_delcnt);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity DPRT_512X9_SRAM_4 is

    port( ELINK_RWA_0         : in    std_logic;
          ELK_RX_SER_WORD_4   : in    std_logic_vector(7 downto 0);
          ELINK_DINA_4        : in    std_logic_vector(7 downto 0);
          ELINK_BLKA_0        : in    std_logic;
          ELKS_ADDRB          : in    std_logic_vector(7 downto 0);
          ELINK_ADDRA_4       : in    std_logic_vector(7 downto 0);
          PATT_ELK_DAT_4      : out   std_logic_vector(7 downto 0);
          ELINK_DOUTA_4       : out   std_logic_vector(7 downto 0);
          ELKS_RWB            : in    std_logic;
          P_USB_MASTER_EN_c_0 : in    std_logic;
          CLK_40M_GL          : in    std_logic;
          CLK60MHZ            : in    std_logic;
          ELKS_RAM_BLKB_EN    : in    std_logic
        );

end DPRT_512X9_SRAM_4;

architecture DEF_ARCH of DPRT_512X9_SRAM_4 is 

  component RAM4K9
    generic (MEMORYFILE:string := "");

    port( ADDRA11 : in    std_logic := 'U';
          ADDRA10 : in    std_logic := 'U';
          ADDRA9  : in    std_logic := 'U';
          ADDRA8  : in    std_logic := 'U';
          ADDRA7  : in    std_logic := 'U';
          ADDRA6  : in    std_logic := 'U';
          ADDRA5  : in    std_logic := 'U';
          ADDRA4  : in    std_logic := 'U';
          ADDRA3  : in    std_logic := 'U';
          ADDRA2  : in    std_logic := 'U';
          ADDRA1  : in    std_logic := 'U';
          ADDRA0  : in    std_logic := 'U';
          ADDRB11 : in    std_logic := 'U';
          ADDRB10 : in    std_logic := 'U';
          ADDRB9  : in    std_logic := 'U';
          ADDRB8  : in    std_logic := 'U';
          ADDRB7  : in    std_logic := 'U';
          ADDRB6  : in    std_logic := 'U';
          ADDRB5  : in    std_logic := 'U';
          ADDRB4  : in    std_logic := 'U';
          ADDRB3  : in    std_logic := 'U';
          ADDRB2  : in    std_logic := 'U';
          ADDRB1  : in    std_logic := 'U';
          ADDRB0  : in    std_logic := 'U';
          DINA8   : in    std_logic := 'U';
          DINA7   : in    std_logic := 'U';
          DINA6   : in    std_logic := 'U';
          DINA5   : in    std_logic := 'U';
          DINA4   : in    std_logic := 'U';
          DINA3   : in    std_logic := 'U';
          DINA2   : in    std_logic := 'U';
          DINA1   : in    std_logic := 'U';
          DINA0   : in    std_logic := 'U';
          DINB8   : in    std_logic := 'U';
          DINB7   : in    std_logic := 'U';
          DINB6   : in    std_logic := 'U';
          DINB5   : in    std_logic := 'U';
          DINB4   : in    std_logic := 'U';
          DINB3   : in    std_logic := 'U';
          DINB2   : in    std_logic := 'U';
          DINB1   : in    std_logic := 'U';
          DINB0   : in    std_logic := 'U';
          WIDTHA0 : in    std_logic := 'U';
          WIDTHA1 : in    std_logic := 'U';
          WIDTHB0 : in    std_logic := 'U';
          WIDTHB1 : in    std_logic := 'U';
          PIPEA   : in    std_logic := 'U';
          PIPEB   : in    std_logic := 'U';
          WMODEA  : in    std_logic := 'U';
          WMODEB  : in    std_logic := 'U';
          BLKA    : in    std_logic := 'U';
          BLKB    : in    std_logic := 'U';
          WENA    : in    std_logic := 'U';
          WENB    : in    std_logic := 'U';
          CLKA    : in    std_logic := 'U';
          CLKB    : in    std_logic := 'U';
          RESET   : in    std_logic := 'U';
          DOUTA8  : out   std_logic;
          DOUTA7  : out   std_logic;
          DOUTA6  : out   std_logic;
          DOUTA5  : out   std_logic;
          DOUTA4  : out   std_logic;
          DOUTA3  : out   std_logic;
          DOUTA2  : out   std_logic;
          DOUTA1  : out   std_logic;
          DOUTA0  : out   std_logic;
          DOUTB8  : out   std_logic;
          DOUTB7  : out   std_logic;
          DOUTB6  : out   std_logic;
          DOUTB5  : out   std_logic;
          DOUTB4  : out   std_logic;
          DOUTB3  : out   std_logic;
          DOUTB2  : out   std_logic;
          DOUTB1  : out   std_logic;
          DOUTB0  : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \DOUTA_1[8]\, \DOUTB_1[8]\, DPRT_512X9_SRAM_4_GND, 
        DPRT_512X9_SRAM_4_VCC : std_logic;

begin 


    DPRT_512X9_SRAM_R0C0 : RAM4K9
      generic map(MEMORYFILE => "DPRT_512X9_SRAM_R0C0.mem")

      port map(ADDRA11 => DPRT_512X9_SRAM_4_GND, ADDRA10 => 
        DPRT_512X9_SRAM_4_GND, ADDRA9 => DPRT_512X9_SRAM_4_GND, 
        ADDRA8 => DPRT_512X9_SRAM_4_GND, ADDRA7 => 
        ELINK_ADDRA_4(7), ADDRA6 => ELINK_ADDRA_4(6), ADDRA5 => 
        ELINK_ADDRA_4(5), ADDRA4 => ELINK_ADDRA_4(4), ADDRA3 => 
        ELINK_ADDRA_4(3), ADDRA2 => ELINK_ADDRA_4(2), ADDRA1 => 
        ELINK_ADDRA_4(1), ADDRA0 => ELINK_ADDRA_4(0), ADDRB11 => 
        DPRT_512X9_SRAM_4_GND, ADDRB10 => DPRT_512X9_SRAM_4_GND, 
        ADDRB9 => DPRT_512X9_SRAM_4_GND, ADDRB8 => 
        DPRT_512X9_SRAM_4_GND, ADDRB7 => ELKS_ADDRB(7), ADDRB6
         => ELKS_ADDRB(6), ADDRB5 => ELKS_ADDRB(5), ADDRB4 => 
        ELKS_ADDRB(4), ADDRB3 => ELKS_ADDRB(3), ADDRB2 => 
        ELKS_ADDRB(2), ADDRB1 => ELKS_ADDRB(1), ADDRB0 => 
        ELKS_ADDRB(0), DINA8 => DPRT_512X9_SRAM_4_GND, DINA7 => 
        ELINK_DINA_4(7), DINA6 => ELINK_DINA_4(6), DINA5 => 
        ELINK_DINA_4(5), DINA4 => ELINK_DINA_4(4), DINA3 => 
        ELINK_DINA_4(3), DINA2 => ELINK_DINA_4(2), DINA1 => 
        ELINK_DINA_4(1), DINA0 => ELINK_DINA_4(0), DINB8 => 
        DPRT_512X9_SRAM_4_GND, DINB7 => ELK_RX_SER_WORD_4(7), 
        DINB6 => ELK_RX_SER_WORD_4(6), DINB5 => 
        ELK_RX_SER_WORD_4(5), DINB4 => ELK_RX_SER_WORD_4(4), 
        DINB3 => ELK_RX_SER_WORD_4(3), DINB2 => 
        ELK_RX_SER_WORD_4(2), DINB1 => ELK_RX_SER_WORD_4(1), 
        DINB0 => ELK_RX_SER_WORD_4(0), WIDTHA0 => 
        DPRT_512X9_SRAM_4_VCC, WIDTHA1 => DPRT_512X9_SRAM_4_VCC, 
        WIDTHB0 => DPRT_512X9_SRAM_4_VCC, WIDTHB1 => 
        DPRT_512X9_SRAM_4_VCC, PIPEA => DPRT_512X9_SRAM_4_VCC, 
        PIPEB => DPRT_512X9_SRAM_4_VCC, WMODEA => 
        DPRT_512X9_SRAM_4_GND, WMODEB => DPRT_512X9_SRAM_4_GND, 
        BLKA => ELINK_BLKA_0, BLKB => ELKS_RAM_BLKB_EN, WENA => 
        ELINK_RWA_0, WENB => ELKS_RWB, CLKA => CLK60MHZ, CLKB => 
        CLK_40M_GL, RESET => P_USB_MASTER_EN_c_0, DOUTA8 => 
        \DOUTA_1[8]\, DOUTA7 => ELINK_DOUTA_4(7), DOUTA6 => 
        ELINK_DOUTA_4(6), DOUTA5 => ELINK_DOUTA_4(5), DOUTA4 => 
        ELINK_DOUTA_4(4), DOUTA3 => ELINK_DOUTA_4(3), DOUTA2 => 
        ELINK_DOUTA_4(2), DOUTA1 => ELINK_DOUTA_4(1), DOUTA0 => 
        ELINK_DOUTA_4(0), DOUTB8 => \DOUTB_1[8]\, DOUTB7 => 
        PATT_ELK_DAT_4(7), DOUTB6 => PATT_ELK_DAT_4(6), DOUTB5
         => PATT_ELK_DAT_4(5), DOUTB4 => PATT_ELK_DAT_4(4), 
        DOUTB3 => PATT_ELK_DAT_4(3), DOUTB2 => PATT_ELK_DAT_4(2), 
        DOUTB1 => PATT_ELK_DAT_4(1), DOUTB0 => PATT_ELK_DAT_4(0));
    
    VCC_i : VCC
      port map(Y => DPRT_512X9_SRAM_4_VCC);
    
    GND_i : GND
      port map(Y => DPRT_512X9_SRAM_4_GND);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity DPRT_512X9_SRAM_19 is

    port( ELINK_RWA_0         : in    std_logic;
          ELK_RX_SER_WORD_19  : in    std_logic_vector(7 downto 0);
          ELINK_DINA_19       : in    std_logic_vector(7 downto 0);
          ELINK_BLKA_0        : in    std_logic;
          ELKS_ADDRB          : in    std_logic_vector(7 downto 0);
          ELINK_ADDRA_19      : in    std_logic_vector(7 downto 0);
          PATT_ELK_DAT_19     : out   std_logic_vector(7 downto 0);
          ELINK_DOUTA_19      : out   std_logic_vector(7 downto 0);
          ELKS_RWB            : in    std_logic;
          P_USB_MASTER_EN_c_0 : in    std_logic;
          CLK_40M_GL          : in    std_logic;
          CLK60MHZ            : in    std_logic;
          ELKS_RAM_BLKB_EN    : in    std_logic
        );

end DPRT_512X9_SRAM_19;

architecture DEF_ARCH of DPRT_512X9_SRAM_19 is 

  component RAM4K9
    generic (MEMORYFILE:string := "");

    port( ADDRA11 : in    std_logic := 'U';
          ADDRA10 : in    std_logic := 'U';
          ADDRA9  : in    std_logic := 'U';
          ADDRA8  : in    std_logic := 'U';
          ADDRA7  : in    std_logic := 'U';
          ADDRA6  : in    std_logic := 'U';
          ADDRA5  : in    std_logic := 'U';
          ADDRA4  : in    std_logic := 'U';
          ADDRA3  : in    std_logic := 'U';
          ADDRA2  : in    std_logic := 'U';
          ADDRA1  : in    std_logic := 'U';
          ADDRA0  : in    std_logic := 'U';
          ADDRB11 : in    std_logic := 'U';
          ADDRB10 : in    std_logic := 'U';
          ADDRB9  : in    std_logic := 'U';
          ADDRB8  : in    std_logic := 'U';
          ADDRB7  : in    std_logic := 'U';
          ADDRB6  : in    std_logic := 'U';
          ADDRB5  : in    std_logic := 'U';
          ADDRB4  : in    std_logic := 'U';
          ADDRB3  : in    std_logic := 'U';
          ADDRB2  : in    std_logic := 'U';
          ADDRB1  : in    std_logic := 'U';
          ADDRB0  : in    std_logic := 'U';
          DINA8   : in    std_logic := 'U';
          DINA7   : in    std_logic := 'U';
          DINA6   : in    std_logic := 'U';
          DINA5   : in    std_logic := 'U';
          DINA4   : in    std_logic := 'U';
          DINA3   : in    std_logic := 'U';
          DINA2   : in    std_logic := 'U';
          DINA1   : in    std_logic := 'U';
          DINA0   : in    std_logic := 'U';
          DINB8   : in    std_logic := 'U';
          DINB7   : in    std_logic := 'U';
          DINB6   : in    std_logic := 'U';
          DINB5   : in    std_logic := 'U';
          DINB4   : in    std_logic := 'U';
          DINB3   : in    std_logic := 'U';
          DINB2   : in    std_logic := 'U';
          DINB1   : in    std_logic := 'U';
          DINB0   : in    std_logic := 'U';
          WIDTHA0 : in    std_logic := 'U';
          WIDTHA1 : in    std_logic := 'U';
          WIDTHB0 : in    std_logic := 'U';
          WIDTHB1 : in    std_logic := 'U';
          PIPEA   : in    std_logic := 'U';
          PIPEB   : in    std_logic := 'U';
          WMODEA  : in    std_logic := 'U';
          WMODEB  : in    std_logic := 'U';
          BLKA    : in    std_logic := 'U';
          BLKB    : in    std_logic := 'U';
          WENA    : in    std_logic := 'U';
          WENB    : in    std_logic := 'U';
          CLKA    : in    std_logic := 'U';
          CLKB    : in    std_logic := 'U';
          RESET   : in    std_logic := 'U';
          DOUTA8  : out   std_logic;
          DOUTA7  : out   std_logic;
          DOUTA6  : out   std_logic;
          DOUTA5  : out   std_logic;
          DOUTA4  : out   std_logic;
          DOUTA3  : out   std_logic;
          DOUTA2  : out   std_logic;
          DOUTA1  : out   std_logic;
          DOUTA0  : out   std_logic;
          DOUTB8  : out   std_logic;
          DOUTB7  : out   std_logic;
          DOUTB6  : out   std_logic;
          DOUTB5  : out   std_logic;
          DOUTB4  : out   std_logic;
          DOUTB3  : out   std_logic;
          DOUTB2  : out   std_logic;
          DOUTB1  : out   std_logic;
          DOUTB0  : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \DOUTA_1[8]\, \DOUTB_1[8]\, DPRT_512X9_SRAM_19_GND, 
        DPRT_512X9_SRAM_19_VCC : std_logic;

begin 


    DPRT_512X9_SRAM_R0C0 : RAM4K9
      generic map(MEMORYFILE => "DPRT_512X9_SRAM_R0C0.mem")

      port map(ADDRA11 => DPRT_512X9_SRAM_19_GND, ADDRA10 => 
        DPRT_512X9_SRAM_19_GND, ADDRA9 => DPRT_512X9_SRAM_19_GND, 
        ADDRA8 => DPRT_512X9_SRAM_19_GND, ADDRA7 => 
        ELINK_ADDRA_19(7), ADDRA6 => ELINK_ADDRA_19(6), ADDRA5
         => ELINK_ADDRA_19(5), ADDRA4 => ELINK_ADDRA_19(4), 
        ADDRA3 => ELINK_ADDRA_19(3), ADDRA2 => ELINK_ADDRA_19(2), 
        ADDRA1 => ELINK_ADDRA_19(1), ADDRA0 => ELINK_ADDRA_19(0), 
        ADDRB11 => DPRT_512X9_SRAM_19_GND, ADDRB10 => 
        DPRT_512X9_SRAM_19_GND, ADDRB9 => DPRT_512X9_SRAM_19_GND, 
        ADDRB8 => DPRT_512X9_SRAM_19_GND, ADDRB7 => ELKS_ADDRB(7), 
        ADDRB6 => ELKS_ADDRB(6), ADDRB5 => ELKS_ADDRB(5), ADDRB4
         => ELKS_ADDRB(4), ADDRB3 => ELKS_ADDRB(3), ADDRB2 => 
        ELKS_ADDRB(2), ADDRB1 => ELKS_ADDRB(1), ADDRB0 => 
        ELKS_ADDRB(0), DINA8 => DPRT_512X9_SRAM_19_GND, DINA7 => 
        ELINK_DINA_19(7), DINA6 => ELINK_DINA_19(6), DINA5 => 
        ELINK_DINA_19(5), DINA4 => ELINK_DINA_19(4), DINA3 => 
        ELINK_DINA_19(3), DINA2 => ELINK_DINA_19(2), DINA1 => 
        ELINK_DINA_19(1), DINA0 => ELINK_DINA_19(0), DINB8 => 
        DPRT_512X9_SRAM_19_GND, DINB7 => ELK_RX_SER_WORD_19(7), 
        DINB6 => ELK_RX_SER_WORD_19(6), DINB5 => 
        ELK_RX_SER_WORD_19(5), DINB4 => ELK_RX_SER_WORD_19(4), 
        DINB3 => ELK_RX_SER_WORD_19(3), DINB2 => 
        ELK_RX_SER_WORD_19(2), DINB1 => ELK_RX_SER_WORD_19(1), 
        DINB0 => ELK_RX_SER_WORD_19(0), WIDTHA0 => 
        DPRT_512X9_SRAM_19_VCC, WIDTHA1 => DPRT_512X9_SRAM_19_VCC, 
        WIDTHB0 => DPRT_512X9_SRAM_19_VCC, WIDTHB1 => 
        DPRT_512X9_SRAM_19_VCC, PIPEA => DPRT_512X9_SRAM_19_VCC, 
        PIPEB => DPRT_512X9_SRAM_19_VCC, WMODEA => 
        DPRT_512X9_SRAM_19_GND, WMODEB => DPRT_512X9_SRAM_19_GND, 
        BLKA => ELINK_BLKA_0, BLKB => ELKS_RAM_BLKB_EN, WENA => 
        ELINK_RWA_0, WENB => ELKS_RWB, CLKA => CLK60MHZ, CLKB => 
        CLK_40M_GL, RESET => P_USB_MASTER_EN_c_0, DOUTA8 => 
        \DOUTA_1[8]\, DOUTA7 => ELINK_DOUTA_19(7), DOUTA6 => 
        ELINK_DOUTA_19(6), DOUTA5 => ELINK_DOUTA_19(5), DOUTA4
         => ELINK_DOUTA_19(4), DOUTA3 => ELINK_DOUTA_19(3), 
        DOUTA2 => ELINK_DOUTA_19(2), DOUTA1 => ELINK_DOUTA_19(1), 
        DOUTA0 => ELINK_DOUTA_19(0), DOUTB8 => \DOUTB_1[8]\, 
        DOUTB7 => PATT_ELK_DAT_19(7), DOUTB6 => 
        PATT_ELK_DAT_19(6), DOUTB5 => PATT_ELK_DAT_19(5), DOUTB4
         => PATT_ELK_DAT_19(4), DOUTB3 => PATT_ELK_DAT_19(3), 
        DOUTB2 => PATT_ELK_DAT_19(2), DOUTB1 => 
        PATT_ELK_DAT_19(1), DOUTB0 => PATT_ELK_DAT_19(0));
    
    VCC_i : VCC
      port map(Y => DPRT_512X9_SRAM_19_VCC);
    
    GND_i : GND
      port map(Y => DPRT_512X9_SRAM_19_GND);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity DPRT_512X9_SRAM_7 is

    port( ELINK_RWA_0         : in    std_logic;
          ELK_RX_SER_WORD_7   : in    std_logic_vector(7 downto 0);
          ELINK_DINA_7        : in    std_logic_vector(7 downto 0);
          ELINK_BLKA_0        : in    std_logic;
          ELKS_ADDRB_0_d0     : in    std_logic;
          ELKS_ADDRB_1        : in    std_logic;
          ELKS_ADDRB_3        : in    std_logic;
          ELKS_ADDRB_5        : in    std_logic;
          ELKS_ADDRB_7        : in    std_logic;
          ELKS_ADDRB_0_0      : in    std_logic;
          ELKS_ADDRB_0_2      : in    std_logic;
          ELKS_ADDRB_0_4      : in    std_logic;
          ELINK_ADDRA_7       : in    std_logic_vector(7 downto 0);
          PATT_ELK_DAT_7      : out   std_logic_vector(7 downto 0);
          ELINK_DOUTA_7       : out   std_logic_vector(7 downto 0);
          ELKS_RWB            : in    std_logic;
          P_USB_MASTER_EN_c_0 : in    std_logic;
          CLK_40M_GL          : in    std_logic;
          CLK60MHZ            : in    std_logic;
          ELKS_RAM_BLKB_EN    : in    std_logic
        );

end DPRT_512X9_SRAM_7;

architecture DEF_ARCH of DPRT_512X9_SRAM_7 is 

  component RAM4K9
    generic (MEMORYFILE:string := "");

    port( ADDRA11 : in    std_logic := 'U';
          ADDRA10 : in    std_logic := 'U';
          ADDRA9  : in    std_logic := 'U';
          ADDRA8  : in    std_logic := 'U';
          ADDRA7  : in    std_logic := 'U';
          ADDRA6  : in    std_logic := 'U';
          ADDRA5  : in    std_logic := 'U';
          ADDRA4  : in    std_logic := 'U';
          ADDRA3  : in    std_logic := 'U';
          ADDRA2  : in    std_logic := 'U';
          ADDRA1  : in    std_logic := 'U';
          ADDRA0  : in    std_logic := 'U';
          ADDRB11 : in    std_logic := 'U';
          ADDRB10 : in    std_logic := 'U';
          ADDRB9  : in    std_logic := 'U';
          ADDRB8  : in    std_logic := 'U';
          ADDRB7  : in    std_logic := 'U';
          ADDRB6  : in    std_logic := 'U';
          ADDRB5  : in    std_logic := 'U';
          ADDRB4  : in    std_logic := 'U';
          ADDRB3  : in    std_logic := 'U';
          ADDRB2  : in    std_logic := 'U';
          ADDRB1  : in    std_logic := 'U';
          ADDRB0  : in    std_logic := 'U';
          DINA8   : in    std_logic := 'U';
          DINA7   : in    std_logic := 'U';
          DINA6   : in    std_logic := 'U';
          DINA5   : in    std_logic := 'U';
          DINA4   : in    std_logic := 'U';
          DINA3   : in    std_logic := 'U';
          DINA2   : in    std_logic := 'U';
          DINA1   : in    std_logic := 'U';
          DINA0   : in    std_logic := 'U';
          DINB8   : in    std_logic := 'U';
          DINB7   : in    std_logic := 'U';
          DINB6   : in    std_logic := 'U';
          DINB5   : in    std_logic := 'U';
          DINB4   : in    std_logic := 'U';
          DINB3   : in    std_logic := 'U';
          DINB2   : in    std_logic := 'U';
          DINB1   : in    std_logic := 'U';
          DINB0   : in    std_logic := 'U';
          WIDTHA0 : in    std_logic := 'U';
          WIDTHA1 : in    std_logic := 'U';
          WIDTHB0 : in    std_logic := 'U';
          WIDTHB1 : in    std_logic := 'U';
          PIPEA   : in    std_logic := 'U';
          PIPEB   : in    std_logic := 'U';
          WMODEA  : in    std_logic := 'U';
          WMODEB  : in    std_logic := 'U';
          BLKA    : in    std_logic := 'U';
          BLKB    : in    std_logic := 'U';
          WENA    : in    std_logic := 'U';
          WENB    : in    std_logic := 'U';
          CLKA    : in    std_logic := 'U';
          CLKB    : in    std_logic := 'U';
          RESET   : in    std_logic := 'U';
          DOUTA8  : out   std_logic;
          DOUTA7  : out   std_logic;
          DOUTA6  : out   std_logic;
          DOUTA5  : out   std_logic;
          DOUTA4  : out   std_logic;
          DOUTA3  : out   std_logic;
          DOUTA2  : out   std_logic;
          DOUTA1  : out   std_logic;
          DOUTA0  : out   std_logic;
          DOUTB8  : out   std_logic;
          DOUTB7  : out   std_logic;
          DOUTB6  : out   std_logic;
          DOUTB5  : out   std_logic;
          DOUTB4  : out   std_logic;
          DOUTB3  : out   std_logic;
          DOUTB2  : out   std_logic;
          DOUTB1  : out   std_logic;
          DOUTB0  : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \DOUTA_1[8]\, \DOUTB_1[8]\, DPRT_512X9_SRAM_7_GND, 
        DPRT_512X9_SRAM_7_VCC : std_logic;

begin 


    DPRT_512X9_SRAM_R0C0 : RAM4K9
      generic map(MEMORYFILE => "DPRT_512X9_SRAM_R0C0.mem")

      port map(ADDRA11 => DPRT_512X9_SRAM_7_GND, ADDRA10 => 
        DPRT_512X9_SRAM_7_GND, ADDRA9 => DPRT_512X9_SRAM_7_GND, 
        ADDRA8 => DPRT_512X9_SRAM_7_GND, ADDRA7 => 
        ELINK_ADDRA_7(7), ADDRA6 => ELINK_ADDRA_7(6), ADDRA5 => 
        ELINK_ADDRA_7(5), ADDRA4 => ELINK_ADDRA_7(4), ADDRA3 => 
        ELINK_ADDRA_7(3), ADDRA2 => ELINK_ADDRA_7(2), ADDRA1 => 
        ELINK_ADDRA_7(1), ADDRA0 => ELINK_ADDRA_7(0), ADDRB11 => 
        DPRT_512X9_SRAM_7_GND, ADDRB10 => DPRT_512X9_SRAM_7_GND, 
        ADDRB9 => DPRT_512X9_SRAM_7_GND, ADDRB8 => 
        DPRT_512X9_SRAM_7_GND, ADDRB7 => ELKS_ADDRB_7, ADDRB6 => 
        ELKS_ADDRB_0_4, ADDRB5 => ELKS_ADDRB_5, ADDRB4 => 
        ELKS_ADDRB_0_2, ADDRB3 => ELKS_ADDRB_3, ADDRB2 => 
        ELKS_ADDRB_0_0, ADDRB1 => ELKS_ADDRB_1, ADDRB0 => 
        ELKS_ADDRB_0_d0, DINA8 => DPRT_512X9_SRAM_7_GND, DINA7
         => ELINK_DINA_7(7), DINA6 => ELINK_DINA_7(6), DINA5 => 
        ELINK_DINA_7(5), DINA4 => ELINK_DINA_7(4), DINA3 => 
        ELINK_DINA_7(3), DINA2 => ELINK_DINA_7(2), DINA1 => 
        ELINK_DINA_7(1), DINA0 => ELINK_DINA_7(0), DINB8 => 
        DPRT_512X9_SRAM_7_GND, DINB7 => ELK_RX_SER_WORD_7(7), 
        DINB6 => ELK_RX_SER_WORD_7(6), DINB5 => 
        ELK_RX_SER_WORD_7(5), DINB4 => ELK_RX_SER_WORD_7(4), 
        DINB3 => ELK_RX_SER_WORD_7(3), DINB2 => 
        ELK_RX_SER_WORD_7(2), DINB1 => ELK_RX_SER_WORD_7(1), 
        DINB0 => ELK_RX_SER_WORD_7(0), WIDTHA0 => 
        DPRT_512X9_SRAM_7_VCC, WIDTHA1 => DPRT_512X9_SRAM_7_VCC, 
        WIDTHB0 => DPRT_512X9_SRAM_7_VCC, WIDTHB1 => 
        DPRT_512X9_SRAM_7_VCC, PIPEA => DPRT_512X9_SRAM_7_VCC, 
        PIPEB => DPRT_512X9_SRAM_7_VCC, WMODEA => 
        DPRT_512X9_SRAM_7_GND, WMODEB => DPRT_512X9_SRAM_7_GND, 
        BLKA => ELINK_BLKA_0, BLKB => ELKS_RAM_BLKB_EN, WENA => 
        ELINK_RWA_0, WENB => ELKS_RWB, CLKA => CLK60MHZ, CLKB => 
        CLK_40M_GL, RESET => P_USB_MASTER_EN_c_0, DOUTA8 => 
        \DOUTA_1[8]\, DOUTA7 => ELINK_DOUTA_7(7), DOUTA6 => 
        ELINK_DOUTA_7(6), DOUTA5 => ELINK_DOUTA_7(5), DOUTA4 => 
        ELINK_DOUTA_7(4), DOUTA3 => ELINK_DOUTA_7(3), DOUTA2 => 
        ELINK_DOUTA_7(2), DOUTA1 => ELINK_DOUTA_7(1), DOUTA0 => 
        ELINK_DOUTA_7(0), DOUTB8 => \DOUTB_1[8]\, DOUTB7 => 
        PATT_ELK_DAT_7(7), DOUTB6 => PATT_ELK_DAT_7(6), DOUTB5
         => PATT_ELK_DAT_7(5), DOUTB4 => PATT_ELK_DAT_7(4), 
        DOUTB3 => PATT_ELK_DAT_7(3), DOUTB2 => PATT_ELK_DAT_7(2), 
        DOUTB1 => PATT_ELK_DAT_7(1), DOUTB0 => PATT_ELK_DAT_7(0));
    
    VCC_i : VCC
      port map(Y => DPRT_512X9_SRAM_7_VCC);
    
    GND_i : GND
      port map(Y => DPRT_512X9_SRAM_7_GND);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity CLK60M_TO_40M_4 is

    port( TFC_STRT_ADDR_0       : in    std_logic_vector(7 downto 0);
          TFC_STRT_ADDR         : out   std_logic_vector(7 downto 0);
          P_MASTER_POR_B_c_22   : in    std_logic;
          P_MASTER_POR_B_c_21   : in    std_logic;
          P_MASTER_POR_B_c_32_0 : in    std_logic;
          P_MASTER_POR_B_c_32   : in    std_logic;
          P_MASTER_POR_B_c_17   : in    std_logic;
          P_MASTER_POR_B_c_27   : in    std_logic;
          CLK_40M_GL            : in    std_logic
        );

end CLK60M_TO_40M_4;

architecture DEF_ARCH of CLK60M_TO_40M_4 is 

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component XO1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component MX2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal un1_SAMP_TWO_NE_4, un1_SAMP_TWO_5, un1_SAMP_TWO_4, 
        un1_SAMP_TWO_NE_1, un1_SAMP_TWO_NE_3, \TFC_STRT_ADDR[3]\, 
        \SAMP_TWO[3]_net_1\, un1_SAMP_TWO_2, un1_SAMP_TWO_NE_2, 
        \TFC_STRT_ADDR[1]\, \SAMP_TWO[1]_net_1\, un1_SAMP_TWO_0, 
        \TFC_STRT_ADDR[6]\, \SAMP_TWO[6]_net_1\, un1_SAMP_TWO_7, 
        n_sync_sm3, SUM1_0, \DELCNT[1]_net_1\, \DELCNT[0]_net_1\, 
        \SAMP_TWO[0]_net_1\, \TFC_STRT_ADDR[0]\, 
        \SAMP_TWO[2]_net_1\, \TFC_STRT_ADDR[2]\, \N_DELCNT[0]\, 
        \SYNC_SM[0]_net_1\, un7_delcnt, \N_SYNC_SM[0]\, 
        \SAMP_TWO[7]_net_1\, \TFC_STRT_ADDR[7]\, 
        \SAMP_TWO[5]_net_1\, \TFC_STRT_ADDR[5]\, 
        \SAMP_TWO[4]_net_1\, \TFC_STRT_ADDR[4]\, 
        \SAMP_ONE[0]_net_1\, \SAMP_ONE[1]_net_1\, 
        \SAMP_ONE[2]_net_1\, \SAMP_ONE[3]_net_1\, 
        \SAMP_ONE[4]_net_1\, \SAMP_ONE[5]_net_1\, 
        \SAMP_ONE[6]_net_1\, \SAMP_ONE[7]_net_1\, \GND\, \VCC\
         : std_logic;

begin 

    TFC_STRT_ADDR(7) <= \TFC_STRT_ADDR[7]\;
    TFC_STRT_ADDR(6) <= \TFC_STRT_ADDR[6]\;
    TFC_STRT_ADDR(5) <= \TFC_STRT_ADDR[5]\;
    TFC_STRT_ADDR(4) <= \TFC_STRT_ADDR[4]\;
    TFC_STRT_ADDR(3) <= \TFC_STRT_ADDR[3]\;
    TFC_STRT_ADDR(2) <= \TFC_STRT_ADDR[2]\;
    TFC_STRT_ADDR(1) <= \TFC_STRT_ADDR[1]\;
    TFC_STRT_ADDR(0) <= \TFC_STRT_ADDR[0]\;

    \SAMP_ONE[2]\ : DFN1C0
      port map(D => TFC_STRT_ADDR_0(2), CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_32, Q => \SAMP_ONE[2]_net_1\);
    
    \SYNC_SM_RNO_6[0]\ : XOR2
      port map(A => \SAMP_TWO[5]_net_1\, B => \TFC_STRT_ADDR[5]\, 
        Y => un1_SAMP_TWO_5);
    
    \DELCNT_RNIJAHN[1]\ : NOR2B
      port map(A => \DELCNT[1]_net_1\, B => \DELCNT[0]_net_1\, Y
         => un7_delcnt);
    
    \LOCAL_REG_VAL[3]\ : DFN1E1C0
      port map(D => \SAMP_TWO[3]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_17, E => un7_delcnt, Q => 
        \TFC_STRT_ADDR[3]\);
    
    \SYNC_SM[0]\ : DFN1C0
      port map(D => \N_SYNC_SM[0]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_27, Q => \SYNC_SM[0]_net_1\);
    
    \SYNC_SM_RNO_5[0]\ : XOR2
      port map(A => \SAMP_TWO[0]_net_1\, B => \TFC_STRT_ADDR[0]\, 
        Y => un1_SAMP_TWO_0);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \DELCNT[1]\ : DFN1C0
      port map(D => SUM1_0, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_32, Q => \DELCNT[1]_net_1\);
    
    \LOCAL_REG_VAL[5]\ : DFN1E1C0
      port map(D => \SAMP_TWO[5]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_17, E => un7_delcnt, Q => 
        \TFC_STRT_ADDR[5]\);
    
    \SYNC_SM_RNO_1[0]\ : XO1
      port map(A => \TFC_STRT_ADDR[3]\, B => \SAMP_TWO[3]_net_1\, 
        C => un1_SAMP_TWO_2, Y => un1_SAMP_TWO_NE_3);
    
    \SAMP_TWO[0]\ : DFN1C0
      port map(D => \SAMP_ONE[0]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_21, Q => \SAMP_TWO[0]_net_1\);
    
    \SAMP_ONE[1]\ : DFN1C0
      port map(D => TFC_STRT_ADDR_0(1), CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_32, Q => \SAMP_ONE[1]_net_1\);
    
    \SAMP_TWO[1]\ : DFN1C0
      port map(D => \SAMP_ONE[1]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_22, Q => \SAMP_TWO[1]_net_1\);
    
    \SYNC_SM_RNO_3[0]\ : OR3
      port map(A => un1_SAMP_TWO_5, B => un1_SAMP_TWO_4, C => 
        un1_SAMP_TWO_NE_1, Y => un1_SAMP_TWO_NE_4);
    
    \SYNC_SM_RNO_9[0]\ : XOR2
      port map(A => \SAMP_TWO[7]_net_1\, B => \TFC_STRT_ADDR[7]\, 
        Y => un1_SAMP_TWO_7);
    
    un2_n_delcnt_1_1_SUM1 : XOR2
      port map(A => \DELCNT[1]_net_1\, B => \DELCNT[0]_net_1\, Y
         => SUM1_0);
    
    \SAMP_TWO[3]\ : DFN1C0
      port map(D => \SAMP_ONE[3]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_22, Q => \SAMP_TWO[3]_net_1\);
    
    \SYNC_SM_RNO_8[0]\ : XO1
      port map(A => \TFC_STRT_ADDR[6]\, B => \SAMP_TWO[6]_net_1\, 
        C => un1_SAMP_TWO_7, Y => un1_SAMP_TWO_NE_1);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \SYNC_SM_RNO_4[0]\ : XOR2
      port map(A => \SAMP_TWO[2]_net_1\, B => \TFC_STRT_ADDR[2]\, 
        Y => un1_SAMP_TWO_2);
    
    \SYNC_SM_RNO[0]\ : MX2B
      port map(A => n_sync_sm3, B => un7_delcnt, S => 
        \SYNC_SM[0]_net_1\, Y => \N_SYNC_SM[0]\);
    
    \SAMP_ONE[4]\ : DFN1C0
      port map(D => TFC_STRT_ADDR_0(4), CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_32_0, Q => \SAMP_ONE[4]_net_1\);
    
    \LOCAL_REG_VAL[2]\ : DFN1E1C0
      port map(D => \SAMP_TWO[2]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_17, E => un7_delcnt, Q => 
        \TFC_STRT_ADDR[2]\);
    
    \SAMP_TWO[5]\ : DFN1C0
      port map(D => \SAMP_ONE[5]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_22, Q => \SAMP_TWO[5]_net_1\);
    
    \SAMP_TWO[4]\ : DFN1C0
      port map(D => \SAMP_ONE[4]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_22, Q => \SAMP_TWO[4]_net_1\);
    
    \SAMP_TWO[2]\ : DFN1C0
      port map(D => \SAMP_ONE[2]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_22, Q => \SAMP_TWO[2]_net_1\);
    
    \DELCNT_RNO[0]\ : NOR2A
      port map(A => \SYNC_SM[0]_net_1\, B => \DELCNT[0]_net_1\, Y
         => \N_DELCNT[0]\);
    
    \LOCAL_REG_VAL[0]\ : DFN1E1C0
      port map(D => \SAMP_TWO[0]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_17, E => un7_delcnt, Q => 
        \TFC_STRT_ADDR[0]\);
    
    \LOCAL_REG_VAL[7]\ : DFN1E1C0
      port map(D => \SAMP_TWO[7]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_17, E => un7_delcnt, Q => 
        \TFC_STRT_ADDR[7]\);
    
    \SYNC_SM_RNO_0[0]\ : OR3
      port map(A => un1_SAMP_TWO_NE_3, B => un1_SAMP_TWO_NE_2, C
         => un1_SAMP_TWO_NE_4, Y => n_sync_sm3);
    
    \DELCNT[0]\ : DFN1C0
      port map(D => \N_DELCNT[0]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_32, Q => \DELCNT[0]_net_1\);
    
    \LOCAL_REG_VAL[4]\ : DFN1E1C0
      port map(D => \SAMP_TWO[4]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_17, E => un7_delcnt, Q => 
        \TFC_STRT_ADDR[4]\);
    
    \SAMP_ONE[7]\ : DFN1C0
      port map(D => TFC_STRT_ADDR_0(7), CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_32_0, Q => \SAMP_ONE[7]_net_1\);
    
    \SYNC_SM_RNO_2[0]\ : XO1
      port map(A => \TFC_STRT_ADDR[1]\, B => \SAMP_TWO[1]_net_1\, 
        C => un1_SAMP_TWO_0, Y => un1_SAMP_TWO_NE_2);
    
    \SAMP_TWO[7]\ : DFN1C0
      port map(D => \SAMP_ONE[7]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_22, Q => \SAMP_TWO[7]_net_1\);
    
    \SAMP_ONE[5]\ : DFN1C0
      port map(D => TFC_STRT_ADDR_0(5), CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_32_0, Q => \SAMP_ONE[5]_net_1\);
    
    \LOCAL_REG_VAL[6]\ : DFN1E1C0
      port map(D => \SAMP_TWO[6]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_17, E => un7_delcnt, Q => 
        \TFC_STRT_ADDR[6]\);
    
    \SYNC_SM_RNO_7[0]\ : XOR2
      port map(A => \SAMP_TWO[4]_net_1\, B => \TFC_STRT_ADDR[4]\, 
        Y => un1_SAMP_TWO_4);
    
    \SAMP_ONE[6]\ : DFN1C0
      port map(D => TFC_STRT_ADDR_0(6), CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_32_0, Q => \SAMP_ONE[6]_net_1\);
    
    \SAMP_ONE[0]\ : DFN1C0
      port map(D => TFC_STRT_ADDR_0(0), CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_32, Q => \SAMP_ONE[0]_net_1\);
    
    \LOCAL_REG_VAL[1]\ : DFN1E1C0
      port map(D => \SAMP_TWO[1]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_17, E => un7_delcnt, Q => 
        \TFC_STRT_ADDR[1]\);
    
    \SAMP_TWO[6]\ : DFN1C0
      port map(D => \SAMP_ONE[6]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_22, Q => \SAMP_TWO[6]_net_1\);
    
    \SAMP_ONE[3]\ : DFN1C0
      port map(D => TFC_STRT_ADDR_0(3), CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_32, Q => \SAMP_ONE[3]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity DPRT_512X9_SRAM_9 is

    port( ELINK_RWA_0         : in    std_logic;
          ELK_RX_SER_WORD_9   : in    std_logic_vector(7 downto 0);
          ELINK_DINA_9        : in    std_logic_vector(7 downto 0);
          ELINK_BLKA_0        : in    std_logic;
          ELKS_ADDRB          : in    std_logic_vector(7 downto 0);
          ELINK_ADDRA_9       : in    std_logic_vector(7 downto 0);
          PATT_ELK_DAT_9      : out   std_logic_vector(7 downto 0);
          ELINK_DOUTA_9       : out   std_logic_vector(7 downto 0);
          ELKS_RWB            : in    std_logic;
          P_USB_MASTER_EN_c_0 : in    std_logic;
          CLK_40M_GL          : in    std_logic;
          CLK60MHZ            : in    std_logic;
          ELKS_RAM_BLKB_EN    : in    std_logic
        );

end DPRT_512X9_SRAM_9;

architecture DEF_ARCH of DPRT_512X9_SRAM_9 is 

  component RAM4K9
    generic (MEMORYFILE:string := "");

    port( ADDRA11 : in    std_logic := 'U';
          ADDRA10 : in    std_logic := 'U';
          ADDRA9  : in    std_logic := 'U';
          ADDRA8  : in    std_logic := 'U';
          ADDRA7  : in    std_logic := 'U';
          ADDRA6  : in    std_logic := 'U';
          ADDRA5  : in    std_logic := 'U';
          ADDRA4  : in    std_logic := 'U';
          ADDRA3  : in    std_logic := 'U';
          ADDRA2  : in    std_logic := 'U';
          ADDRA1  : in    std_logic := 'U';
          ADDRA0  : in    std_logic := 'U';
          ADDRB11 : in    std_logic := 'U';
          ADDRB10 : in    std_logic := 'U';
          ADDRB9  : in    std_logic := 'U';
          ADDRB8  : in    std_logic := 'U';
          ADDRB7  : in    std_logic := 'U';
          ADDRB6  : in    std_logic := 'U';
          ADDRB5  : in    std_logic := 'U';
          ADDRB4  : in    std_logic := 'U';
          ADDRB3  : in    std_logic := 'U';
          ADDRB2  : in    std_logic := 'U';
          ADDRB1  : in    std_logic := 'U';
          ADDRB0  : in    std_logic := 'U';
          DINA8   : in    std_logic := 'U';
          DINA7   : in    std_logic := 'U';
          DINA6   : in    std_logic := 'U';
          DINA5   : in    std_logic := 'U';
          DINA4   : in    std_logic := 'U';
          DINA3   : in    std_logic := 'U';
          DINA2   : in    std_logic := 'U';
          DINA1   : in    std_logic := 'U';
          DINA0   : in    std_logic := 'U';
          DINB8   : in    std_logic := 'U';
          DINB7   : in    std_logic := 'U';
          DINB6   : in    std_logic := 'U';
          DINB5   : in    std_logic := 'U';
          DINB4   : in    std_logic := 'U';
          DINB3   : in    std_logic := 'U';
          DINB2   : in    std_logic := 'U';
          DINB1   : in    std_logic := 'U';
          DINB0   : in    std_logic := 'U';
          WIDTHA0 : in    std_logic := 'U';
          WIDTHA1 : in    std_logic := 'U';
          WIDTHB0 : in    std_logic := 'U';
          WIDTHB1 : in    std_logic := 'U';
          PIPEA   : in    std_logic := 'U';
          PIPEB   : in    std_logic := 'U';
          WMODEA  : in    std_logic := 'U';
          WMODEB  : in    std_logic := 'U';
          BLKA    : in    std_logic := 'U';
          BLKB    : in    std_logic := 'U';
          WENA    : in    std_logic := 'U';
          WENB    : in    std_logic := 'U';
          CLKA    : in    std_logic := 'U';
          CLKB    : in    std_logic := 'U';
          RESET   : in    std_logic := 'U';
          DOUTA8  : out   std_logic;
          DOUTA7  : out   std_logic;
          DOUTA6  : out   std_logic;
          DOUTA5  : out   std_logic;
          DOUTA4  : out   std_logic;
          DOUTA3  : out   std_logic;
          DOUTA2  : out   std_logic;
          DOUTA1  : out   std_logic;
          DOUTA0  : out   std_logic;
          DOUTB8  : out   std_logic;
          DOUTB7  : out   std_logic;
          DOUTB6  : out   std_logic;
          DOUTB5  : out   std_logic;
          DOUTB4  : out   std_logic;
          DOUTB3  : out   std_logic;
          DOUTB2  : out   std_logic;
          DOUTB1  : out   std_logic;
          DOUTB0  : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \DOUTA_1[8]\, \DOUTB_1[8]\, DPRT_512X9_SRAM_9_GND, 
        DPRT_512X9_SRAM_9_VCC : std_logic;

begin 


    DPRT_512X9_SRAM_R0C0 : RAM4K9
      generic map(MEMORYFILE => "DPRT_512X9_SRAM_R0C0.mem")

      port map(ADDRA11 => DPRT_512X9_SRAM_9_GND, ADDRA10 => 
        DPRT_512X9_SRAM_9_GND, ADDRA9 => DPRT_512X9_SRAM_9_GND, 
        ADDRA8 => DPRT_512X9_SRAM_9_GND, ADDRA7 => 
        ELINK_ADDRA_9(7), ADDRA6 => ELINK_ADDRA_9(6), ADDRA5 => 
        ELINK_ADDRA_9(5), ADDRA4 => ELINK_ADDRA_9(4), ADDRA3 => 
        ELINK_ADDRA_9(3), ADDRA2 => ELINK_ADDRA_9(2), ADDRA1 => 
        ELINK_ADDRA_9(1), ADDRA0 => ELINK_ADDRA_9(0), ADDRB11 => 
        DPRT_512X9_SRAM_9_GND, ADDRB10 => DPRT_512X9_SRAM_9_GND, 
        ADDRB9 => DPRT_512X9_SRAM_9_GND, ADDRB8 => 
        DPRT_512X9_SRAM_9_GND, ADDRB7 => ELKS_ADDRB(7), ADDRB6
         => ELKS_ADDRB(6), ADDRB5 => ELKS_ADDRB(5), ADDRB4 => 
        ELKS_ADDRB(4), ADDRB3 => ELKS_ADDRB(3), ADDRB2 => 
        ELKS_ADDRB(2), ADDRB1 => ELKS_ADDRB(1), ADDRB0 => 
        ELKS_ADDRB(0), DINA8 => DPRT_512X9_SRAM_9_GND, DINA7 => 
        ELINK_DINA_9(7), DINA6 => ELINK_DINA_9(6), DINA5 => 
        ELINK_DINA_9(5), DINA4 => ELINK_DINA_9(4), DINA3 => 
        ELINK_DINA_9(3), DINA2 => ELINK_DINA_9(2), DINA1 => 
        ELINK_DINA_9(1), DINA0 => ELINK_DINA_9(0), DINB8 => 
        DPRT_512X9_SRAM_9_GND, DINB7 => ELK_RX_SER_WORD_9(7), 
        DINB6 => ELK_RX_SER_WORD_9(6), DINB5 => 
        ELK_RX_SER_WORD_9(5), DINB4 => ELK_RX_SER_WORD_9(4), 
        DINB3 => ELK_RX_SER_WORD_9(3), DINB2 => 
        ELK_RX_SER_WORD_9(2), DINB1 => ELK_RX_SER_WORD_9(1), 
        DINB0 => ELK_RX_SER_WORD_9(0), WIDTHA0 => 
        DPRT_512X9_SRAM_9_VCC, WIDTHA1 => DPRT_512X9_SRAM_9_VCC, 
        WIDTHB0 => DPRT_512X9_SRAM_9_VCC, WIDTHB1 => 
        DPRT_512X9_SRAM_9_VCC, PIPEA => DPRT_512X9_SRAM_9_VCC, 
        PIPEB => DPRT_512X9_SRAM_9_VCC, WMODEA => 
        DPRT_512X9_SRAM_9_GND, WMODEB => DPRT_512X9_SRAM_9_GND, 
        BLKA => ELINK_BLKA_0, BLKB => ELKS_RAM_BLKB_EN, WENA => 
        ELINK_RWA_0, WENB => ELKS_RWB, CLKA => CLK60MHZ, CLKB => 
        CLK_40M_GL, RESET => P_USB_MASTER_EN_c_0, DOUTA8 => 
        \DOUTA_1[8]\, DOUTA7 => ELINK_DOUTA_9(7), DOUTA6 => 
        ELINK_DOUTA_9(6), DOUTA5 => ELINK_DOUTA_9(5), DOUTA4 => 
        ELINK_DOUTA_9(4), DOUTA3 => ELINK_DOUTA_9(3), DOUTA2 => 
        ELINK_DOUTA_9(2), DOUTA1 => ELINK_DOUTA_9(1), DOUTA0 => 
        ELINK_DOUTA_9(0), DOUTB8 => \DOUTB_1[8]\, DOUTB7 => 
        PATT_ELK_DAT_9(7), DOUTB6 => PATT_ELK_DAT_9(6), DOUTB5
         => PATT_ELK_DAT_9(5), DOUTB4 => PATT_ELK_DAT_9(4), 
        DOUTB3 => PATT_ELK_DAT_9(3), DOUTB2 => PATT_ELK_DAT_9(2), 
        DOUTB1 => PATT_ELK_DAT_9(1), DOUTB0 => PATT_ELK_DAT_9(0));
    
    VCC_i : VCC
      port map(Y => DPRT_512X9_SRAM_9_VCC);
    
    GND_i : GND
      port map(Y => DPRT_512X9_SRAM_9_GND);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity DPRT_512X9_SRAM_18 is

    port( ELINK_RWA_0         : in    std_logic;
          ELK_RX_SER_WORD_18  : in    std_logic_vector(7 downto 0);
          ELINK_DINA_18       : in    std_logic_vector(7 downto 0);
          ELINK_BLKA_0        : in    std_logic;
          ELKS_ADDRB_0_d0     : in    std_logic;
          ELKS_ADDRB_1        : in    std_logic;
          ELKS_ADDRB_3        : in    std_logic;
          ELKS_ADDRB_5        : in    std_logic;
          ELKS_ADDRB_7        : in    std_logic;
          ELKS_ADDRB_0_0      : in    std_logic;
          ELKS_ADDRB_0_2      : in    std_logic;
          ELKS_ADDRB_0_4      : in    std_logic;
          ELINK_ADDRA_18      : in    std_logic_vector(7 downto 0);
          PATT_ELK_DAT_18     : out   std_logic_vector(7 downto 0);
          ELINK_DOUTA_18      : out   std_logic_vector(7 downto 0);
          ELKS_RWB            : in    std_logic;
          P_USB_MASTER_EN_c_0 : in    std_logic;
          CLK_40M_GL          : in    std_logic;
          CLK60MHZ            : in    std_logic;
          ELKS_RAM_BLKB_EN    : in    std_logic
        );

end DPRT_512X9_SRAM_18;

architecture DEF_ARCH of DPRT_512X9_SRAM_18 is 

  component RAM4K9
    generic (MEMORYFILE:string := "");

    port( ADDRA11 : in    std_logic := 'U';
          ADDRA10 : in    std_logic := 'U';
          ADDRA9  : in    std_logic := 'U';
          ADDRA8  : in    std_logic := 'U';
          ADDRA7  : in    std_logic := 'U';
          ADDRA6  : in    std_logic := 'U';
          ADDRA5  : in    std_logic := 'U';
          ADDRA4  : in    std_logic := 'U';
          ADDRA3  : in    std_logic := 'U';
          ADDRA2  : in    std_logic := 'U';
          ADDRA1  : in    std_logic := 'U';
          ADDRA0  : in    std_logic := 'U';
          ADDRB11 : in    std_logic := 'U';
          ADDRB10 : in    std_logic := 'U';
          ADDRB9  : in    std_logic := 'U';
          ADDRB8  : in    std_logic := 'U';
          ADDRB7  : in    std_logic := 'U';
          ADDRB6  : in    std_logic := 'U';
          ADDRB5  : in    std_logic := 'U';
          ADDRB4  : in    std_logic := 'U';
          ADDRB3  : in    std_logic := 'U';
          ADDRB2  : in    std_logic := 'U';
          ADDRB1  : in    std_logic := 'U';
          ADDRB0  : in    std_logic := 'U';
          DINA8   : in    std_logic := 'U';
          DINA7   : in    std_logic := 'U';
          DINA6   : in    std_logic := 'U';
          DINA5   : in    std_logic := 'U';
          DINA4   : in    std_logic := 'U';
          DINA3   : in    std_logic := 'U';
          DINA2   : in    std_logic := 'U';
          DINA1   : in    std_logic := 'U';
          DINA0   : in    std_logic := 'U';
          DINB8   : in    std_logic := 'U';
          DINB7   : in    std_logic := 'U';
          DINB6   : in    std_logic := 'U';
          DINB5   : in    std_logic := 'U';
          DINB4   : in    std_logic := 'U';
          DINB3   : in    std_logic := 'U';
          DINB2   : in    std_logic := 'U';
          DINB1   : in    std_logic := 'U';
          DINB0   : in    std_logic := 'U';
          WIDTHA0 : in    std_logic := 'U';
          WIDTHA1 : in    std_logic := 'U';
          WIDTHB0 : in    std_logic := 'U';
          WIDTHB1 : in    std_logic := 'U';
          PIPEA   : in    std_logic := 'U';
          PIPEB   : in    std_logic := 'U';
          WMODEA  : in    std_logic := 'U';
          WMODEB  : in    std_logic := 'U';
          BLKA    : in    std_logic := 'U';
          BLKB    : in    std_logic := 'U';
          WENA    : in    std_logic := 'U';
          WENB    : in    std_logic := 'U';
          CLKA    : in    std_logic := 'U';
          CLKB    : in    std_logic := 'U';
          RESET   : in    std_logic := 'U';
          DOUTA8  : out   std_logic;
          DOUTA7  : out   std_logic;
          DOUTA6  : out   std_logic;
          DOUTA5  : out   std_logic;
          DOUTA4  : out   std_logic;
          DOUTA3  : out   std_logic;
          DOUTA2  : out   std_logic;
          DOUTA1  : out   std_logic;
          DOUTA0  : out   std_logic;
          DOUTB8  : out   std_logic;
          DOUTB7  : out   std_logic;
          DOUTB6  : out   std_logic;
          DOUTB5  : out   std_logic;
          DOUTB4  : out   std_logic;
          DOUTB3  : out   std_logic;
          DOUTB2  : out   std_logic;
          DOUTB1  : out   std_logic;
          DOUTB0  : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \DOUTA_1[8]\, \DOUTB_1[8]\, DPRT_512X9_SRAM_18_GND, 
        DPRT_512X9_SRAM_18_VCC : std_logic;

begin 


    DPRT_512X9_SRAM_R0C0 : RAM4K9
      generic map(MEMORYFILE => "DPRT_512X9_SRAM_R0C0.mem")

      port map(ADDRA11 => DPRT_512X9_SRAM_18_GND, ADDRA10 => 
        DPRT_512X9_SRAM_18_GND, ADDRA9 => DPRT_512X9_SRAM_18_GND, 
        ADDRA8 => DPRT_512X9_SRAM_18_GND, ADDRA7 => 
        ELINK_ADDRA_18(7), ADDRA6 => ELINK_ADDRA_18(6), ADDRA5
         => ELINK_ADDRA_18(5), ADDRA4 => ELINK_ADDRA_18(4), 
        ADDRA3 => ELINK_ADDRA_18(3), ADDRA2 => ELINK_ADDRA_18(2), 
        ADDRA1 => ELINK_ADDRA_18(1), ADDRA0 => ELINK_ADDRA_18(0), 
        ADDRB11 => DPRT_512X9_SRAM_18_GND, ADDRB10 => 
        DPRT_512X9_SRAM_18_GND, ADDRB9 => DPRT_512X9_SRAM_18_GND, 
        ADDRB8 => DPRT_512X9_SRAM_18_GND, ADDRB7 => ELKS_ADDRB_7, 
        ADDRB6 => ELKS_ADDRB_0_4, ADDRB5 => ELKS_ADDRB_5, ADDRB4
         => ELKS_ADDRB_0_2, ADDRB3 => ELKS_ADDRB_3, ADDRB2 => 
        ELKS_ADDRB_0_0, ADDRB1 => ELKS_ADDRB_1, ADDRB0 => 
        ELKS_ADDRB_0_d0, DINA8 => DPRT_512X9_SRAM_18_GND, DINA7
         => ELINK_DINA_18(7), DINA6 => ELINK_DINA_18(6), DINA5
         => ELINK_DINA_18(5), DINA4 => ELINK_DINA_18(4), DINA3
         => ELINK_DINA_18(3), DINA2 => ELINK_DINA_18(2), DINA1
         => ELINK_DINA_18(1), DINA0 => ELINK_DINA_18(0), DINB8
         => DPRT_512X9_SRAM_18_GND, DINB7 => 
        ELK_RX_SER_WORD_18(7), DINB6 => ELK_RX_SER_WORD_18(6), 
        DINB5 => ELK_RX_SER_WORD_18(5), DINB4 => 
        ELK_RX_SER_WORD_18(4), DINB3 => ELK_RX_SER_WORD_18(3), 
        DINB2 => ELK_RX_SER_WORD_18(2), DINB1 => 
        ELK_RX_SER_WORD_18(1), DINB0 => ELK_RX_SER_WORD_18(0), 
        WIDTHA0 => DPRT_512X9_SRAM_18_VCC, WIDTHA1 => 
        DPRT_512X9_SRAM_18_VCC, WIDTHB0 => DPRT_512X9_SRAM_18_VCC, 
        WIDTHB1 => DPRT_512X9_SRAM_18_VCC, PIPEA => 
        DPRT_512X9_SRAM_18_VCC, PIPEB => DPRT_512X9_SRAM_18_VCC, 
        WMODEA => DPRT_512X9_SRAM_18_GND, WMODEB => 
        DPRT_512X9_SRAM_18_GND, BLKA => ELINK_BLKA_0, BLKB => 
        ELKS_RAM_BLKB_EN, WENA => ELINK_RWA_0, WENB => ELKS_RWB, 
        CLKA => CLK60MHZ, CLKB => CLK_40M_GL, RESET => 
        P_USB_MASTER_EN_c_0, DOUTA8 => \DOUTA_1[8]\, DOUTA7 => 
        ELINK_DOUTA_18(7), DOUTA6 => ELINK_DOUTA_18(6), DOUTA5
         => ELINK_DOUTA_18(5), DOUTA4 => ELINK_DOUTA_18(4), 
        DOUTA3 => ELINK_DOUTA_18(3), DOUTA2 => ELINK_DOUTA_18(2), 
        DOUTA1 => ELINK_DOUTA_18(1), DOUTA0 => ELINK_DOUTA_18(0), 
        DOUTB8 => \DOUTB_1[8]\, DOUTB7 => PATT_ELK_DAT_18(7), 
        DOUTB6 => PATT_ELK_DAT_18(6), DOUTB5 => 
        PATT_ELK_DAT_18(5), DOUTB4 => PATT_ELK_DAT_18(4), DOUTB3
         => PATT_ELK_DAT_18(3), DOUTB2 => PATT_ELK_DAT_18(2), 
        DOUTB1 => PATT_ELK_DAT_18(1), DOUTB0 => 
        PATT_ELK_DAT_18(0));
    
    VCC_i : VCC
      port map(Y => DPRT_512X9_SRAM_18_VCC);
    
    GND_i : GND
      port map(Y => DPRT_512X9_SRAM_18_GND);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity DPRT_512X9_SRAM_15 is

    port( ELINK_RWA_0         : in    std_logic;
          ELK_RX_SER_WORD_15  : in    std_logic_vector(7 downto 0);
          ELINK_DINA_15       : in    std_logic_vector(7 downto 0);
          ELINK_BLKA_0        : in    std_logic;
          ELKS_ADDRB          : in    std_logic_vector(7 downto 0);
          ELINK_ADDRA_15      : in    std_logic_vector(7 downto 0);
          PATT_ELK_DAT_15     : out   std_logic_vector(7 downto 0);
          ELINK_DOUTA_15      : out   std_logic_vector(7 downto 0);
          ELKS_RWB            : in    std_logic;
          P_USB_MASTER_EN_c_0 : in    std_logic;
          CLK_40M_GL          : in    std_logic;
          CLK60MHZ            : in    std_logic;
          ELKS_RAM_BLKB_EN    : in    std_logic
        );

end DPRT_512X9_SRAM_15;

architecture DEF_ARCH of DPRT_512X9_SRAM_15 is 

  component RAM4K9
    generic (MEMORYFILE:string := "");

    port( ADDRA11 : in    std_logic := 'U';
          ADDRA10 : in    std_logic := 'U';
          ADDRA9  : in    std_logic := 'U';
          ADDRA8  : in    std_logic := 'U';
          ADDRA7  : in    std_logic := 'U';
          ADDRA6  : in    std_logic := 'U';
          ADDRA5  : in    std_logic := 'U';
          ADDRA4  : in    std_logic := 'U';
          ADDRA3  : in    std_logic := 'U';
          ADDRA2  : in    std_logic := 'U';
          ADDRA1  : in    std_logic := 'U';
          ADDRA0  : in    std_logic := 'U';
          ADDRB11 : in    std_logic := 'U';
          ADDRB10 : in    std_logic := 'U';
          ADDRB9  : in    std_logic := 'U';
          ADDRB8  : in    std_logic := 'U';
          ADDRB7  : in    std_logic := 'U';
          ADDRB6  : in    std_logic := 'U';
          ADDRB5  : in    std_logic := 'U';
          ADDRB4  : in    std_logic := 'U';
          ADDRB3  : in    std_logic := 'U';
          ADDRB2  : in    std_logic := 'U';
          ADDRB1  : in    std_logic := 'U';
          ADDRB0  : in    std_logic := 'U';
          DINA8   : in    std_logic := 'U';
          DINA7   : in    std_logic := 'U';
          DINA6   : in    std_logic := 'U';
          DINA5   : in    std_logic := 'U';
          DINA4   : in    std_logic := 'U';
          DINA3   : in    std_logic := 'U';
          DINA2   : in    std_logic := 'U';
          DINA1   : in    std_logic := 'U';
          DINA0   : in    std_logic := 'U';
          DINB8   : in    std_logic := 'U';
          DINB7   : in    std_logic := 'U';
          DINB6   : in    std_logic := 'U';
          DINB5   : in    std_logic := 'U';
          DINB4   : in    std_logic := 'U';
          DINB3   : in    std_logic := 'U';
          DINB2   : in    std_logic := 'U';
          DINB1   : in    std_logic := 'U';
          DINB0   : in    std_logic := 'U';
          WIDTHA0 : in    std_logic := 'U';
          WIDTHA1 : in    std_logic := 'U';
          WIDTHB0 : in    std_logic := 'U';
          WIDTHB1 : in    std_logic := 'U';
          PIPEA   : in    std_logic := 'U';
          PIPEB   : in    std_logic := 'U';
          WMODEA  : in    std_logic := 'U';
          WMODEB  : in    std_logic := 'U';
          BLKA    : in    std_logic := 'U';
          BLKB    : in    std_logic := 'U';
          WENA    : in    std_logic := 'U';
          WENB    : in    std_logic := 'U';
          CLKA    : in    std_logic := 'U';
          CLKB    : in    std_logic := 'U';
          RESET   : in    std_logic := 'U';
          DOUTA8  : out   std_logic;
          DOUTA7  : out   std_logic;
          DOUTA6  : out   std_logic;
          DOUTA5  : out   std_logic;
          DOUTA4  : out   std_logic;
          DOUTA3  : out   std_logic;
          DOUTA2  : out   std_logic;
          DOUTA1  : out   std_logic;
          DOUTA0  : out   std_logic;
          DOUTB8  : out   std_logic;
          DOUTB7  : out   std_logic;
          DOUTB6  : out   std_logic;
          DOUTB5  : out   std_logic;
          DOUTB4  : out   std_logic;
          DOUTB3  : out   std_logic;
          DOUTB2  : out   std_logic;
          DOUTB1  : out   std_logic;
          DOUTB0  : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \DOUTA_1[8]\, \DOUTB_1[8]\, DPRT_512X9_SRAM_15_GND, 
        DPRT_512X9_SRAM_15_VCC : std_logic;

begin 


    DPRT_512X9_SRAM_R0C0 : RAM4K9
      generic map(MEMORYFILE => "DPRT_512X9_SRAM_R0C0.mem")

      port map(ADDRA11 => DPRT_512X9_SRAM_15_GND, ADDRA10 => 
        DPRT_512X9_SRAM_15_GND, ADDRA9 => DPRT_512X9_SRAM_15_GND, 
        ADDRA8 => DPRT_512X9_SRAM_15_GND, ADDRA7 => 
        ELINK_ADDRA_15(7), ADDRA6 => ELINK_ADDRA_15(6), ADDRA5
         => ELINK_ADDRA_15(5), ADDRA4 => ELINK_ADDRA_15(4), 
        ADDRA3 => ELINK_ADDRA_15(3), ADDRA2 => ELINK_ADDRA_15(2), 
        ADDRA1 => ELINK_ADDRA_15(1), ADDRA0 => ELINK_ADDRA_15(0), 
        ADDRB11 => DPRT_512X9_SRAM_15_GND, ADDRB10 => 
        DPRT_512X9_SRAM_15_GND, ADDRB9 => DPRT_512X9_SRAM_15_GND, 
        ADDRB8 => DPRT_512X9_SRAM_15_GND, ADDRB7 => ELKS_ADDRB(7), 
        ADDRB6 => ELKS_ADDRB(6), ADDRB5 => ELKS_ADDRB(5), ADDRB4
         => ELKS_ADDRB(4), ADDRB3 => ELKS_ADDRB(3), ADDRB2 => 
        ELKS_ADDRB(2), ADDRB1 => ELKS_ADDRB(1), ADDRB0 => 
        ELKS_ADDRB(0), DINA8 => DPRT_512X9_SRAM_15_GND, DINA7 => 
        ELINK_DINA_15(7), DINA6 => ELINK_DINA_15(6), DINA5 => 
        ELINK_DINA_15(5), DINA4 => ELINK_DINA_15(4), DINA3 => 
        ELINK_DINA_15(3), DINA2 => ELINK_DINA_15(2), DINA1 => 
        ELINK_DINA_15(1), DINA0 => ELINK_DINA_15(0), DINB8 => 
        DPRT_512X9_SRAM_15_GND, DINB7 => ELK_RX_SER_WORD_15(7), 
        DINB6 => ELK_RX_SER_WORD_15(6), DINB5 => 
        ELK_RX_SER_WORD_15(5), DINB4 => ELK_RX_SER_WORD_15(4), 
        DINB3 => ELK_RX_SER_WORD_15(3), DINB2 => 
        ELK_RX_SER_WORD_15(2), DINB1 => ELK_RX_SER_WORD_15(1), 
        DINB0 => ELK_RX_SER_WORD_15(0), WIDTHA0 => 
        DPRT_512X9_SRAM_15_VCC, WIDTHA1 => DPRT_512X9_SRAM_15_VCC, 
        WIDTHB0 => DPRT_512X9_SRAM_15_VCC, WIDTHB1 => 
        DPRT_512X9_SRAM_15_VCC, PIPEA => DPRT_512X9_SRAM_15_VCC, 
        PIPEB => DPRT_512X9_SRAM_15_VCC, WMODEA => 
        DPRT_512X9_SRAM_15_GND, WMODEB => DPRT_512X9_SRAM_15_GND, 
        BLKA => ELINK_BLKA_0, BLKB => ELKS_RAM_BLKB_EN, WENA => 
        ELINK_RWA_0, WENB => ELKS_RWB, CLKA => CLK60MHZ, CLKB => 
        CLK_40M_GL, RESET => P_USB_MASTER_EN_c_0, DOUTA8 => 
        \DOUTA_1[8]\, DOUTA7 => ELINK_DOUTA_15(7), DOUTA6 => 
        ELINK_DOUTA_15(6), DOUTA5 => ELINK_DOUTA_15(5), DOUTA4
         => ELINK_DOUTA_15(4), DOUTA3 => ELINK_DOUTA_15(3), 
        DOUTA2 => ELINK_DOUTA_15(2), DOUTA1 => ELINK_DOUTA_15(1), 
        DOUTA0 => ELINK_DOUTA_15(0), DOUTB8 => \DOUTB_1[8]\, 
        DOUTB7 => PATT_ELK_DAT_15(7), DOUTB6 => 
        PATT_ELK_DAT_15(6), DOUTB5 => PATT_ELK_DAT_15(5), DOUTB4
         => PATT_ELK_DAT_15(4), DOUTB3 => PATT_ELK_DAT_15(3), 
        DOUTB2 => PATT_ELK_DAT_15(2), DOUTB1 => 
        PATT_ELK_DAT_15(1), DOUTB0 => PATT_ELK_DAT_15(0));
    
    VCC_i : VCC
      port map(Y => DPRT_512X9_SRAM_15_VCC);
    
    GND_i : GND
      port map(Y => DPRT_512X9_SRAM_15_GND);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity DPRT_512X9_SRAM is

    port( TFC_RX_SER_WORD     : in    std_logic_vector(7 downto 0);
          TFC_DINA            : in    std_logic_vector(7 downto 0);
          TFC_ADDRB           : in    std_logic_vector(7 downto 0);
          TFC_ADDRA           : in    std_logic_vector(7 downto 0);
          PATT_TFC_DAT        : out   std_logic_vector(7 downto 0);
          TFC_DOUTA           : out   std_logic_vector(7 downto 0);
          TFC_RWB             : in    std_logic;
          TFC_RWA             : in    std_logic;
          P_USB_MASTER_EN_c_0 : in    std_logic;
          CLK_40M_GL          : in    std_logic;
          CLK60MHZ            : in    std_logic;
          TFC_RAM_BLKB_EN     : in    std_logic;
          TFC_BLKA            : in    std_logic
        );

end DPRT_512X9_SRAM;

architecture DEF_ARCH of DPRT_512X9_SRAM is 

  component RAM4K9
    generic (MEMORYFILE:string := "");

    port( ADDRA11 : in    std_logic := 'U';
          ADDRA10 : in    std_logic := 'U';
          ADDRA9  : in    std_logic := 'U';
          ADDRA8  : in    std_logic := 'U';
          ADDRA7  : in    std_logic := 'U';
          ADDRA6  : in    std_logic := 'U';
          ADDRA5  : in    std_logic := 'U';
          ADDRA4  : in    std_logic := 'U';
          ADDRA3  : in    std_logic := 'U';
          ADDRA2  : in    std_logic := 'U';
          ADDRA1  : in    std_logic := 'U';
          ADDRA0  : in    std_logic := 'U';
          ADDRB11 : in    std_logic := 'U';
          ADDRB10 : in    std_logic := 'U';
          ADDRB9  : in    std_logic := 'U';
          ADDRB8  : in    std_logic := 'U';
          ADDRB7  : in    std_logic := 'U';
          ADDRB6  : in    std_logic := 'U';
          ADDRB5  : in    std_logic := 'U';
          ADDRB4  : in    std_logic := 'U';
          ADDRB3  : in    std_logic := 'U';
          ADDRB2  : in    std_logic := 'U';
          ADDRB1  : in    std_logic := 'U';
          ADDRB0  : in    std_logic := 'U';
          DINA8   : in    std_logic := 'U';
          DINA7   : in    std_logic := 'U';
          DINA6   : in    std_logic := 'U';
          DINA5   : in    std_logic := 'U';
          DINA4   : in    std_logic := 'U';
          DINA3   : in    std_logic := 'U';
          DINA2   : in    std_logic := 'U';
          DINA1   : in    std_logic := 'U';
          DINA0   : in    std_logic := 'U';
          DINB8   : in    std_logic := 'U';
          DINB7   : in    std_logic := 'U';
          DINB6   : in    std_logic := 'U';
          DINB5   : in    std_logic := 'U';
          DINB4   : in    std_logic := 'U';
          DINB3   : in    std_logic := 'U';
          DINB2   : in    std_logic := 'U';
          DINB1   : in    std_logic := 'U';
          DINB0   : in    std_logic := 'U';
          WIDTHA0 : in    std_logic := 'U';
          WIDTHA1 : in    std_logic := 'U';
          WIDTHB0 : in    std_logic := 'U';
          WIDTHB1 : in    std_logic := 'U';
          PIPEA   : in    std_logic := 'U';
          PIPEB   : in    std_logic := 'U';
          WMODEA  : in    std_logic := 'U';
          WMODEB  : in    std_logic := 'U';
          BLKA    : in    std_logic := 'U';
          BLKB    : in    std_logic := 'U';
          WENA    : in    std_logic := 'U';
          WENB    : in    std_logic := 'U';
          CLKA    : in    std_logic := 'U';
          CLKB    : in    std_logic := 'U';
          RESET   : in    std_logic := 'U';
          DOUTA8  : out   std_logic;
          DOUTA7  : out   std_logic;
          DOUTA6  : out   std_logic;
          DOUTA5  : out   std_logic;
          DOUTA4  : out   std_logic;
          DOUTA3  : out   std_logic;
          DOUTA2  : out   std_logic;
          DOUTA1  : out   std_logic;
          DOUTA0  : out   std_logic;
          DOUTB8  : out   std_logic;
          DOUTB7  : out   std_logic;
          DOUTB6  : out   std_logic;
          DOUTB5  : out   std_logic;
          DOUTB4  : out   std_logic;
          DOUTB3  : out   std_logic;
          DOUTB2  : out   std_logic;
          DOUTB1  : out   std_logic;
          DOUTB0  : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \DOUTA_1[8]\, \DOUTB_1[8]\, DPRT_512X9_SRAM_GND, 
        DPRT_512X9_SRAM_VCC : std_logic;

begin 


    DPRT_512X9_SRAM_R0C0 : RAM4K9
      generic map(MEMORYFILE => "DPRT_512X9_SRAM_R0C0.mem")

      port map(ADDRA11 => DPRT_512X9_SRAM_GND, ADDRA10 => 
        DPRT_512X9_SRAM_GND, ADDRA9 => DPRT_512X9_SRAM_GND, 
        ADDRA8 => DPRT_512X9_SRAM_GND, ADDRA7 => TFC_ADDRA(7), 
        ADDRA6 => TFC_ADDRA(6), ADDRA5 => TFC_ADDRA(5), ADDRA4
         => TFC_ADDRA(4), ADDRA3 => TFC_ADDRA(3), ADDRA2 => 
        TFC_ADDRA(2), ADDRA1 => TFC_ADDRA(1), ADDRA0 => 
        TFC_ADDRA(0), ADDRB11 => DPRT_512X9_SRAM_GND, ADDRB10 => 
        DPRT_512X9_SRAM_GND, ADDRB9 => DPRT_512X9_SRAM_GND, 
        ADDRB8 => DPRT_512X9_SRAM_GND, ADDRB7 => TFC_ADDRB(7), 
        ADDRB6 => TFC_ADDRB(6), ADDRB5 => TFC_ADDRB(5), ADDRB4
         => TFC_ADDRB(4), ADDRB3 => TFC_ADDRB(3), ADDRB2 => 
        TFC_ADDRB(2), ADDRB1 => TFC_ADDRB(1), ADDRB0 => 
        TFC_ADDRB(0), DINA8 => DPRT_512X9_SRAM_GND, DINA7 => 
        TFC_DINA(7), DINA6 => TFC_DINA(6), DINA5 => TFC_DINA(5), 
        DINA4 => TFC_DINA(4), DINA3 => TFC_DINA(3), DINA2 => 
        TFC_DINA(2), DINA1 => TFC_DINA(1), DINA0 => TFC_DINA(0), 
        DINB8 => DPRT_512X9_SRAM_GND, DINB7 => TFC_RX_SER_WORD(7), 
        DINB6 => TFC_RX_SER_WORD(6), DINB5 => TFC_RX_SER_WORD(5), 
        DINB4 => TFC_RX_SER_WORD(4), DINB3 => TFC_RX_SER_WORD(3), 
        DINB2 => TFC_RX_SER_WORD(2), DINB1 => TFC_RX_SER_WORD(1), 
        DINB0 => TFC_RX_SER_WORD(0), WIDTHA0 => 
        DPRT_512X9_SRAM_VCC, WIDTHA1 => DPRT_512X9_SRAM_VCC, 
        WIDTHB0 => DPRT_512X9_SRAM_VCC, WIDTHB1 => 
        DPRT_512X9_SRAM_VCC, PIPEA => DPRT_512X9_SRAM_VCC, PIPEB
         => DPRT_512X9_SRAM_VCC, WMODEA => DPRT_512X9_SRAM_GND, 
        WMODEB => DPRT_512X9_SRAM_GND, BLKA => TFC_BLKA, BLKB => 
        TFC_RAM_BLKB_EN, WENA => TFC_RWA, WENB => TFC_RWB, CLKA
         => CLK60MHZ, CLKB => CLK_40M_GL, RESET => 
        P_USB_MASTER_EN_c_0, DOUTA8 => \DOUTA_1[8]\, DOUTA7 => 
        TFC_DOUTA(7), DOUTA6 => TFC_DOUTA(6), DOUTA5 => 
        TFC_DOUTA(5), DOUTA4 => TFC_DOUTA(4), DOUTA3 => 
        TFC_DOUTA(3), DOUTA2 => TFC_DOUTA(2), DOUTA1 => 
        TFC_DOUTA(1), DOUTA0 => TFC_DOUTA(0), DOUTB8 => 
        \DOUTB_1[8]\, DOUTB7 => PATT_TFC_DAT(7), DOUTB6 => 
        PATT_TFC_DAT(6), DOUTB5 => PATT_TFC_DAT(5), DOUTB4 => 
        PATT_TFC_DAT(4), DOUTB3 => PATT_TFC_DAT(3), DOUTB2 => 
        PATT_TFC_DAT(2), DOUTB1 => PATT_TFC_DAT(1), DOUTB0 => 
        PATT_TFC_DAT(0));
    
    VCC_i : VCC
      port map(Y => DPRT_512X9_SRAM_VCC);
    
    GND_i : GND
      port map(Y => DPRT_512X9_SRAM_GND);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity DPRT_512X9_SRAM_10 is

    port( ELINK_RWA_0         : in    std_logic;
          ELK_RX_SER_WORD_10  : in    std_logic_vector(7 downto 0);
          ELINK_DINA_10       : in    std_logic_vector(7 downto 0);
          ELINK_BLKA_0        : in    std_logic;
          ELKS_ADDRB_0_d0     : in    std_logic;
          ELKS_ADDRB_1        : in    std_logic;
          ELKS_ADDRB_3        : in    std_logic;
          ELKS_ADDRB_5        : in    std_logic;
          ELKS_ADDRB_7        : in    std_logic;
          ELKS_ADDRB_0_0      : in    std_logic;
          ELKS_ADDRB_0_2      : in    std_logic;
          ELKS_ADDRB_0_4      : in    std_logic;
          ELINK_ADDRA_10      : in    std_logic_vector(7 downto 0);
          PATT_ELK_DAT_10     : out   std_logic_vector(7 downto 0);
          ELINK_DOUTA_10      : out   std_logic_vector(7 downto 0);
          ELKS_RWB            : in    std_logic;
          P_USB_MASTER_EN_c_0 : in    std_logic;
          CLK_40M_GL          : in    std_logic;
          CLK60MHZ            : in    std_logic;
          ELKS_RAM_BLKB_EN    : in    std_logic
        );

end DPRT_512X9_SRAM_10;

architecture DEF_ARCH of DPRT_512X9_SRAM_10 is 

  component RAM4K9
    generic (MEMORYFILE:string := "");

    port( ADDRA11 : in    std_logic := 'U';
          ADDRA10 : in    std_logic := 'U';
          ADDRA9  : in    std_logic := 'U';
          ADDRA8  : in    std_logic := 'U';
          ADDRA7  : in    std_logic := 'U';
          ADDRA6  : in    std_logic := 'U';
          ADDRA5  : in    std_logic := 'U';
          ADDRA4  : in    std_logic := 'U';
          ADDRA3  : in    std_logic := 'U';
          ADDRA2  : in    std_logic := 'U';
          ADDRA1  : in    std_logic := 'U';
          ADDRA0  : in    std_logic := 'U';
          ADDRB11 : in    std_logic := 'U';
          ADDRB10 : in    std_logic := 'U';
          ADDRB9  : in    std_logic := 'U';
          ADDRB8  : in    std_logic := 'U';
          ADDRB7  : in    std_logic := 'U';
          ADDRB6  : in    std_logic := 'U';
          ADDRB5  : in    std_logic := 'U';
          ADDRB4  : in    std_logic := 'U';
          ADDRB3  : in    std_logic := 'U';
          ADDRB2  : in    std_logic := 'U';
          ADDRB1  : in    std_logic := 'U';
          ADDRB0  : in    std_logic := 'U';
          DINA8   : in    std_logic := 'U';
          DINA7   : in    std_logic := 'U';
          DINA6   : in    std_logic := 'U';
          DINA5   : in    std_logic := 'U';
          DINA4   : in    std_logic := 'U';
          DINA3   : in    std_logic := 'U';
          DINA2   : in    std_logic := 'U';
          DINA1   : in    std_logic := 'U';
          DINA0   : in    std_logic := 'U';
          DINB8   : in    std_logic := 'U';
          DINB7   : in    std_logic := 'U';
          DINB6   : in    std_logic := 'U';
          DINB5   : in    std_logic := 'U';
          DINB4   : in    std_logic := 'U';
          DINB3   : in    std_logic := 'U';
          DINB2   : in    std_logic := 'U';
          DINB1   : in    std_logic := 'U';
          DINB0   : in    std_logic := 'U';
          WIDTHA0 : in    std_logic := 'U';
          WIDTHA1 : in    std_logic := 'U';
          WIDTHB0 : in    std_logic := 'U';
          WIDTHB1 : in    std_logic := 'U';
          PIPEA   : in    std_logic := 'U';
          PIPEB   : in    std_logic := 'U';
          WMODEA  : in    std_logic := 'U';
          WMODEB  : in    std_logic := 'U';
          BLKA    : in    std_logic := 'U';
          BLKB    : in    std_logic := 'U';
          WENA    : in    std_logic := 'U';
          WENB    : in    std_logic := 'U';
          CLKA    : in    std_logic := 'U';
          CLKB    : in    std_logic := 'U';
          RESET   : in    std_logic := 'U';
          DOUTA8  : out   std_logic;
          DOUTA7  : out   std_logic;
          DOUTA6  : out   std_logic;
          DOUTA5  : out   std_logic;
          DOUTA4  : out   std_logic;
          DOUTA3  : out   std_logic;
          DOUTA2  : out   std_logic;
          DOUTA1  : out   std_logic;
          DOUTA0  : out   std_logic;
          DOUTB8  : out   std_logic;
          DOUTB7  : out   std_logic;
          DOUTB6  : out   std_logic;
          DOUTB5  : out   std_logic;
          DOUTB4  : out   std_logic;
          DOUTB3  : out   std_logic;
          DOUTB2  : out   std_logic;
          DOUTB1  : out   std_logic;
          DOUTB0  : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \DOUTA_1[8]\, \DOUTB_1[8]\, DPRT_512X9_SRAM_10_GND, 
        DPRT_512X9_SRAM_10_VCC : std_logic;

begin 


    DPRT_512X9_SRAM_R0C0 : RAM4K9
      generic map(MEMORYFILE => "DPRT_512X9_SRAM_R0C0.mem")

      port map(ADDRA11 => DPRT_512X9_SRAM_10_GND, ADDRA10 => 
        DPRT_512X9_SRAM_10_GND, ADDRA9 => DPRT_512X9_SRAM_10_GND, 
        ADDRA8 => DPRT_512X9_SRAM_10_GND, ADDRA7 => 
        ELINK_ADDRA_10(7), ADDRA6 => ELINK_ADDRA_10(6), ADDRA5
         => ELINK_ADDRA_10(5), ADDRA4 => ELINK_ADDRA_10(4), 
        ADDRA3 => ELINK_ADDRA_10(3), ADDRA2 => ELINK_ADDRA_10(2), 
        ADDRA1 => ELINK_ADDRA_10(1), ADDRA0 => ELINK_ADDRA_10(0), 
        ADDRB11 => DPRT_512X9_SRAM_10_GND, ADDRB10 => 
        DPRT_512X9_SRAM_10_GND, ADDRB9 => DPRT_512X9_SRAM_10_GND, 
        ADDRB8 => DPRT_512X9_SRAM_10_GND, ADDRB7 => ELKS_ADDRB_7, 
        ADDRB6 => ELKS_ADDRB_0_4, ADDRB5 => ELKS_ADDRB_5, ADDRB4
         => ELKS_ADDRB_0_2, ADDRB3 => ELKS_ADDRB_3, ADDRB2 => 
        ELKS_ADDRB_0_0, ADDRB1 => ELKS_ADDRB_1, ADDRB0 => 
        ELKS_ADDRB_0_d0, DINA8 => DPRT_512X9_SRAM_10_GND, DINA7
         => ELINK_DINA_10(7), DINA6 => ELINK_DINA_10(6), DINA5
         => ELINK_DINA_10(5), DINA4 => ELINK_DINA_10(4), DINA3
         => ELINK_DINA_10(3), DINA2 => ELINK_DINA_10(2), DINA1
         => ELINK_DINA_10(1), DINA0 => ELINK_DINA_10(0), DINB8
         => DPRT_512X9_SRAM_10_GND, DINB7 => 
        ELK_RX_SER_WORD_10(7), DINB6 => ELK_RX_SER_WORD_10(6), 
        DINB5 => ELK_RX_SER_WORD_10(5), DINB4 => 
        ELK_RX_SER_WORD_10(4), DINB3 => ELK_RX_SER_WORD_10(3), 
        DINB2 => ELK_RX_SER_WORD_10(2), DINB1 => 
        ELK_RX_SER_WORD_10(1), DINB0 => ELK_RX_SER_WORD_10(0), 
        WIDTHA0 => DPRT_512X9_SRAM_10_VCC, WIDTHA1 => 
        DPRT_512X9_SRAM_10_VCC, WIDTHB0 => DPRT_512X9_SRAM_10_VCC, 
        WIDTHB1 => DPRT_512X9_SRAM_10_VCC, PIPEA => 
        DPRT_512X9_SRAM_10_VCC, PIPEB => DPRT_512X9_SRAM_10_VCC, 
        WMODEA => DPRT_512X9_SRAM_10_GND, WMODEB => 
        DPRT_512X9_SRAM_10_GND, BLKA => ELINK_BLKA_0, BLKB => 
        ELKS_RAM_BLKB_EN, WENA => ELINK_RWA_0, WENB => ELKS_RWB, 
        CLKA => CLK60MHZ, CLKB => CLK_40M_GL, RESET => 
        P_USB_MASTER_EN_c_0, DOUTA8 => \DOUTA_1[8]\, DOUTA7 => 
        ELINK_DOUTA_10(7), DOUTA6 => ELINK_DOUTA_10(6), DOUTA5
         => ELINK_DOUTA_10(5), DOUTA4 => ELINK_DOUTA_10(4), 
        DOUTA3 => ELINK_DOUTA_10(3), DOUTA2 => ELINK_DOUTA_10(2), 
        DOUTA1 => ELINK_DOUTA_10(1), DOUTA0 => ELINK_DOUTA_10(0), 
        DOUTB8 => \DOUTB_1[8]\, DOUTB7 => PATT_ELK_DAT_10(7), 
        DOUTB6 => PATT_ELK_DAT_10(6), DOUTB5 => 
        PATT_ELK_DAT_10(5), DOUTB4 => PATT_ELK_DAT_10(4), DOUTB3
         => PATT_ELK_DAT_10(3), DOUTB2 => PATT_ELK_DAT_10(2), 
        DOUTB1 => PATT_ELK_DAT_10(1), DOUTB0 => 
        PATT_ELK_DAT_10(0));
    
    VCC_i : VCC
      port map(Y => DPRT_512X9_SRAM_10_VCC);
    
    GND_i : GND
      port map(Y => DPRT_512X9_SRAM_10_GND);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity DPRT_512X9_SRAM_8 is

    port( ELINK_RWA_0         : in    std_logic;
          ELK_RX_SER_WORD_8   : in    std_logic_vector(7 downto 0);
          ELINK_DINA_8        : in    std_logic_vector(7 downto 0);
          ELINK_BLKA_0        : in    std_logic;
          ELKS_ADDRB_0_d0     : in    std_logic;
          ELKS_ADDRB_1        : in    std_logic;
          ELKS_ADDRB_3        : in    std_logic;
          ELKS_ADDRB_5        : in    std_logic;
          ELKS_ADDRB_7        : in    std_logic;
          ELKS_ADDRB_0_0      : in    std_logic;
          ELKS_ADDRB_0_2      : in    std_logic;
          ELKS_ADDRB_0_4      : in    std_logic;
          ELINK_ADDRA_8       : in    std_logic_vector(7 downto 0);
          PATT_ELK_DAT_8      : out   std_logic_vector(7 downto 0);
          ELINK_DOUTA_8       : out   std_logic_vector(7 downto 0);
          ELKS_RWB            : in    std_logic;
          P_USB_MASTER_EN_c_0 : in    std_logic;
          CLK_40M_GL          : in    std_logic;
          CLK60MHZ            : in    std_logic;
          ELKS_RAM_BLKB_EN    : in    std_logic
        );

end DPRT_512X9_SRAM_8;

architecture DEF_ARCH of DPRT_512X9_SRAM_8 is 

  component RAM4K9
    generic (MEMORYFILE:string := "");

    port( ADDRA11 : in    std_logic := 'U';
          ADDRA10 : in    std_logic := 'U';
          ADDRA9  : in    std_logic := 'U';
          ADDRA8  : in    std_logic := 'U';
          ADDRA7  : in    std_logic := 'U';
          ADDRA6  : in    std_logic := 'U';
          ADDRA5  : in    std_logic := 'U';
          ADDRA4  : in    std_logic := 'U';
          ADDRA3  : in    std_logic := 'U';
          ADDRA2  : in    std_logic := 'U';
          ADDRA1  : in    std_logic := 'U';
          ADDRA0  : in    std_logic := 'U';
          ADDRB11 : in    std_logic := 'U';
          ADDRB10 : in    std_logic := 'U';
          ADDRB9  : in    std_logic := 'U';
          ADDRB8  : in    std_logic := 'U';
          ADDRB7  : in    std_logic := 'U';
          ADDRB6  : in    std_logic := 'U';
          ADDRB5  : in    std_logic := 'U';
          ADDRB4  : in    std_logic := 'U';
          ADDRB3  : in    std_logic := 'U';
          ADDRB2  : in    std_logic := 'U';
          ADDRB1  : in    std_logic := 'U';
          ADDRB0  : in    std_logic := 'U';
          DINA8   : in    std_logic := 'U';
          DINA7   : in    std_logic := 'U';
          DINA6   : in    std_logic := 'U';
          DINA5   : in    std_logic := 'U';
          DINA4   : in    std_logic := 'U';
          DINA3   : in    std_logic := 'U';
          DINA2   : in    std_logic := 'U';
          DINA1   : in    std_logic := 'U';
          DINA0   : in    std_logic := 'U';
          DINB8   : in    std_logic := 'U';
          DINB7   : in    std_logic := 'U';
          DINB6   : in    std_logic := 'U';
          DINB5   : in    std_logic := 'U';
          DINB4   : in    std_logic := 'U';
          DINB3   : in    std_logic := 'U';
          DINB2   : in    std_logic := 'U';
          DINB1   : in    std_logic := 'U';
          DINB0   : in    std_logic := 'U';
          WIDTHA0 : in    std_logic := 'U';
          WIDTHA1 : in    std_logic := 'U';
          WIDTHB0 : in    std_logic := 'U';
          WIDTHB1 : in    std_logic := 'U';
          PIPEA   : in    std_logic := 'U';
          PIPEB   : in    std_logic := 'U';
          WMODEA  : in    std_logic := 'U';
          WMODEB  : in    std_logic := 'U';
          BLKA    : in    std_logic := 'U';
          BLKB    : in    std_logic := 'U';
          WENA    : in    std_logic := 'U';
          WENB    : in    std_logic := 'U';
          CLKA    : in    std_logic := 'U';
          CLKB    : in    std_logic := 'U';
          RESET   : in    std_logic := 'U';
          DOUTA8  : out   std_logic;
          DOUTA7  : out   std_logic;
          DOUTA6  : out   std_logic;
          DOUTA5  : out   std_logic;
          DOUTA4  : out   std_logic;
          DOUTA3  : out   std_logic;
          DOUTA2  : out   std_logic;
          DOUTA1  : out   std_logic;
          DOUTA0  : out   std_logic;
          DOUTB8  : out   std_logic;
          DOUTB7  : out   std_logic;
          DOUTB6  : out   std_logic;
          DOUTB5  : out   std_logic;
          DOUTB4  : out   std_logic;
          DOUTB3  : out   std_logic;
          DOUTB2  : out   std_logic;
          DOUTB1  : out   std_logic;
          DOUTB0  : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \DOUTA_1[8]\, \DOUTB_1[8]\, DPRT_512X9_SRAM_8_GND, 
        DPRT_512X9_SRAM_8_VCC : std_logic;

begin 


    DPRT_512X9_SRAM_R0C0 : RAM4K9
      generic map(MEMORYFILE => "DPRT_512X9_SRAM_R0C0.mem")

      port map(ADDRA11 => DPRT_512X9_SRAM_8_GND, ADDRA10 => 
        DPRT_512X9_SRAM_8_GND, ADDRA9 => DPRT_512X9_SRAM_8_GND, 
        ADDRA8 => DPRT_512X9_SRAM_8_GND, ADDRA7 => 
        ELINK_ADDRA_8(7), ADDRA6 => ELINK_ADDRA_8(6), ADDRA5 => 
        ELINK_ADDRA_8(5), ADDRA4 => ELINK_ADDRA_8(4), ADDRA3 => 
        ELINK_ADDRA_8(3), ADDRA2 => ELINK_ADDRA_8(2), ADDRA1 => 
        ELINK_ADDRA_8(1), ADDRA0 => ELINK_ADDRA_8(0), ADDRB11 => 
        DPRT_512X9_SRAM_8_GND, ADDRB10 => DPRT_512X9_SRAM_8_GND, 
        ADDRB9 => DPRT_512X9_SRAM_8_GND, ADDRB8 => 
        DPRT_512X9_SRAM_8_GND, ADDRB7 => ELKS_ADDRB_7, ADDRB6 => 
        ELKS_ADDRB_0_4, ADDRB5 => ELKS_ADDRB_5, ADDRB4 => 
        ELKS_ADDRB_0_2, ADDRB3 => ELKS_ADDRB_3, ADDRB2 => 
        ELKS_ADDRB_0_0, ADDRB1 => ELKS_ADDRB_1, ADDRB0 => 
        ELKS_ADDRB_0_d0, DINA8 => DPRT_512X9_SRAM_8_GND, DINA7
         => ELINK_DINA_8(7), DINA6 => ELINK_DINA_8(6), DINA5 => 
        ELINK_DINA_8(5), DINA4 => ELINK_DINA_8(4), DINA3 => 
        ELINK_DINA_8(3), DINA2 => ELINK_DINA_8(2), DINA1 => 
        ELINK_DINA_8(1), DINA0 => ELINK_DINA_8(0), DINB8 => 
        DPRT_512X9_SRAM_8_GND, DINB7 => ELK_RX_SER_WORD_8(7), 
        DINB6 => ELK_RX_SER_WORD_8(6), DINB5 => 
        ELK_RX_SER_WORD_8(5), DINB4 => ELK_RX_SER_WORD_8(4), 
        DINB3 => ELK_RX_SER_WORD_8(3), DINB2 => 
        ELK_RX_SER_WORD_8(2), DINB1 => ELK_RX_SER_WORD_8(1), 
        DINB0 => ELK_RX_SER_WORD_8(0), WIDTHA0 => 
        DPRT_512X9_SRAM_8_VCC, WIDTHA1 => DPRT_512X9_SRAM_8_VCC, 
        WIDTHB0 => DPRT_512X9_SRAM_8_VCC, WIDTHB1 => 
        DPRT_512X9_SRAM_8_VCC, PIPEA => DPRT_512X9_SRAM_8_VCC, 
        PIPEB => DPRT_512X9_SRAM_8_VCC, WMODEA => 
        DPRT_512X9_SRAM_8_GND, WMODEB => DPRT_512X9_SRAM_8_GND, 
        BLKA => ELINK_BLKA_0, BLKB => ELKS_RAM_BLKB_EN, WENA => 
        ELINK_RWA_0, WENB => ELKS_RWB, CLKA => CLK60MHZ, CLKB => 
        CLK_40M_GL, RESET => P_USB_MASTER_EN_c_0, DOUTA8 => 
        \DOUTA_1[8]\, DOUTA7 => ELINK_DOUTA_8(7), DOUTA6 => 
        ELINK_DOUTA_8(6), DOUTA5 => ELINK_DOUTA_8(5), DOUTA4 => 
        ELINK_DOUTA_8(4), DOUTA3 => ELINK_DOUTA_8(3), DOUTA2 => 
        ELINK_DOUTA_8(2), DOUTA1 => ELINK_DOUTA_8(1), DOUTA0 => 
        ELINK_DOUTA_8(0), DOUTB8 => \DOUTB_1[8]\, DOUTB7 => 
        PATT_ELK_DAT_8(7), DOUTB6 => PATT_ELK_DAT_8(6), DOUTB5
         => PATT_ELK_DAT_8(5), DOUTB4 => PATT_ELK_DAT_8(4), 
        DOUTB3 => PATT_ELK_DAT_8(3), DOUTB2 => PATT_ELK_DAT_8(2), 
        DOUTB1 => PATT_ELK_DAT_8(1), DOUTB0 => PATT_ELK_DAT_8(0));
    
    VCC_i : VCC
      port map(Y => DPRT_512X9_SRAM_8_VCC);
    
    GND_i : GND
      port map(Y => DPRT_512X9_SRAM_8_GND);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity DPRT_512X9_SRAM_5 is

    port( ELINK_RWA_0         : in    std_logic;
          ELK_RX_SER_WORD_5   : in    std_logic_vector(7 downto 0);
          ELINK_DINA_5        : in    std_logic_vector(7 downto 0);
          ELINK_BLKA_0        : in    std_logic;
          ELKS_ADDRB_0_d0     : in    std_logic;
          ELKS_ADDRB_1        : in    std_logic;
          ELKS_ADDRB_3        : in    std_logic;
          ELKS_ADDRB_5        : in    std_logic;
          ELKS_ADDRB_7        : in    std_logic;
          ELKS_ADDRB_0_0      : in    std_logic;
          ELKS_ADDRB_0_2      : in    std_logic;
          ELKS_ADDRB_0_4      : in    std_logic;
          ELINK_ADDRA_5       : in    std_logic_vector(7 downto 0);
          PATT_ELK_DAT_5      : out   std_logic_vector(7 downto 0);
          ELINK_DOUTA_5       : out   std_logic_vector(7 downto 0);
          ELKS_RWB            : in    std_logic;
          P_USB_MASTER_EN_c_0 : in    std_logic;
          CLK_40M_GL          : in    std_logic;
          CLK60MHZ            : in    std_logic;
          ELKS_RAM_BLKB_EN    : in    std_logic
        );

end DPRT_512X9_SRAM_5;

architecture DEF_ARCH of DPRT_512X9_SRAM_5 is 

  component RAM4K9
    generic (MEMORYFILE:string := "");

    port( ADDRA11 : in    std_logic := 'U';
          ADDRA10 : in    std_logic := 'U';
          ADDRA9  : in    std_logic := 'U';
          ADDRA8  : in    std_logic := 'U';
          ADDRA7  : in    std_logic := 'U';
          ADDRA6  : in    std_logic := 'U';
          ADDRA5  : in    std_logic := 'U';
          ADDRA4  : in    std_logic := 'U';
          ADDRA3  : in    std_logic := 'U';
          ADDRA2  : in    std_logic := 'U';
          ADDRA1  : in    std_logic := 'U';
          ADDRA0  : in    std_logic := 'U';
          ADDRB11 : in    std_logic := 'U';
          ADDRB10 : in    std_logic := 'U';
          ADDRB9  : in    std_logic := 'U';
          ADDRB8  : in    std_logic := 'U';
          ADDRB7  : in    std_logic := 'U';
          ADDRB6  : in    std_logic := 'U';
          ADDRB5  : in    std_logic := 'U';
          ADDRB4  : in    std_logic := 'U';
          ADDRB3  : in    std_logic := 'U';
          ADDRB2  : in    std_logic := 'U';
          ADDRB1  : in    std_logic := 'U';
          ADDRB0  : in    std_logic := 'U';
          DINA8   : in    std_logic := 'U';
          DINA7   : in    std_logic := 'U';
          DINA6   : in    std_logic := 'U';
          DINA5   : in    std_logic := 'U';
          DINA4   : in    std_logic := 'U';
          DINA3   : in    std_logic := 'U';
          DINA2   : in    std_logic := 'U';
          DINA1   : in    std_logic := 'U';
          DINA0   : in    std_logic := 'U';
          DINB8   : in    std_logic := 'U';
          DINB7   : in    std_logic := 'U';
          DINB6   : in    std_logic := 'U';
          DINB5   : in    std_logic := 'U';
          DINB4   : in    std_logic := 'U';
          DINB3   : in    std_logic := 'U';
          DINB2   : in    std_logic := 'U';
          DINB1   : in    std_logic := 'U';
          DINB0   : in    std_logic := 'U';
          WIDTHA0 : in    std_logic := 'U';
          WIDTHA1 : in    std_logic := 'U';
          WIDTHB0 : in    std_logic := 'U';
          WIDTHB1 : in    std_logic := 'U';
          PIPEA   : in    std_logic := 'U';
          PIPEB   : in    std_logic := 'U';
          WMODEA  : in    std_logic := 'U';
          WMODEB  : in    std_logic := 'U';
          BLKA    : in    std_logic := 'U';
          BLKB    : in    std_logic := 'U';
          WENA    : in    std_logic := 'U';
          WENB    : in    std_logic := 'U';
          CLKA    : in    std_logic := 'U';
          CLKB    : in    std_logic := 'U';
          RESET   : in    std_logic := 'U';
          DOUTA8  : out   std_logic;
          DOUTA7  : out   std_logic;
          DOUTA6  : out   std_logic;
          DOUTA5  : out   std_logic;
          DOUTA4  : out   std_logic;
          DOUTA3  : out   std_logic;
          DOUTA2  : out   std_logic;
          DOUTA1  : out   std_logic;
          DOUTA0  : out   std_logic;
          DOUTB8  : out   std_logic;
          DOUTB7  : out   std_logic;
          DOUTB6  : out   std_logic;
          DOUTB5  : out   std_logic;
          DOUTB4  : out   std_logic;
          DOUTB3  : out   std_logic;
          DOUTB2  : out   std_logic;
          DOUTB1  : out   std_logic;
          DOUTB0  : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \DOUTA_1[8]\, \DOUTB_1[8]\, DPRT_512X9_SRAM_5_GND, 
        DPRT_512X9_SRAM_5_VCC : std_logic;

begin 


    DPRT_512X9_SRAM_R0C0 : RAM4K9
      generic map(MEMORYFILE => "DPRT_512X9_SRAM_R0C0.mem")

      port map(ADDRA11 => DPRT_512X9_SRAM_5_GND, ADDRA10 => 
        DPRT_512X9_SRAM_5_GND, ADDRA9 => DPRT_512X9_SRAM_5_GND, 
        ADDRA8 => DPRT_512X9_SRAM_5_GND, ADDRA7 => 
        ELINK_ADDRA_5(7), ADDRA6 => ELINK_ADDRA_5(6), ADDRA5 => 
        ELINK_ADDRA_5(5), ADDRA4 => ELINK_ADDRA_5(4), ADDRA3 => 
        ELINK_ADDRA_5(3), ADDRA2 => ELINK_ADDRA_5(2), ADDRA1 => 
        ELINK_ADDRA_5(1), ADDRA0 => ELINK_ADDRA_5(0), ADDRB11 => 
        DPRT_512X9_SRAM_5_GND, ADDRB10 => DPRT_512X9_SRAM_5_GND, 
        ADDRB9 => DPRT_512X9_SRAM_5_GND, ADDRB8 => 
        DPRT_512X9_SRAM_5_GND, ADDRB7 => ELKS_ADDRB_7, ADDRB6 => 
        ELKS_ADDRB_0_4, ADDRB5 => ELKS_ADDRB_5, ADDRB4 => 
        ELKS_ADDRB_0_2, ADDRB3 => ELKS_ADDRB_3, ADDRB2 => 
        ELKS_ADDRB_0_0, ADDRB1 => ELKS_ADDRB_1, ADDRB0 => 
        ELKS_ADDRB_0_d0, DINA8 => DPRT_512X9_SRAM_5_GND, DINA7
         => ELINK_DINA_5(7), DINA6 => ELINK_DINA_5(6), DINA5 => 
        ELINK_DINA_5(5), DINA4 => ELINK_DINA_5(4), DINA3 => 
        ELINK_DINA_5(3), DINA2 => ELINK_DINA_5(2), DINA1 => 
        ELINK_DINA_5(1), DINA0 => ELINK_DINA_5(0), DINB8 => 
        DPRT_512X9_SRAM_5_GND, DINB7 => ELK_RX_SER_WORD_5(7), 
        DINB6 => ELK_RX_SER_WORD_5(6), DINB5 => 
        ELK_RX_SER_WORD_5(5), DINB4 => ELK_RX_SER_WORD_5(4), 
        DINB3 => ELK_RX_SER_WORD_5(3), DINB2 => 
        ELK_RX_SER_WORD_5(2), DINB1 => ELK_RX_SER_WORD_5(1), 
        DINB0 => ELK_RX_SER_WORD_5(0), WIDTHA0 => 
        DPRT_512X9_SRAM_5_VCC, WIDTHA1 => DPRT_512X9_SRAM_5_VCC, 
        WIDTHB0 => DPRT_512X9_SRAM_5_VCC, WIDTHB1 => 
        DPRT_512X9_SRAM_5_VCC, PIPEA => DPRT_512X9_SRAM_5_VCC, 
        PIPEB => DPRT_512X9_SRAM_5_VCC, WMODEA => 
        DPRT_512X9_SRAM_5_GND, WMODEB => DPRT_512X9_SRAM_5_GND, 
        BLKA => ELINK_BLKA_0, BLKB => ELKS_RAM_BLKB_EN, WENA => 
        ELINK_RWA_0, WENB => ELKS_RWB, CLKA => CLK60MHZ, CLKB => 
        CLK_40M_GL, RESET => P_USB_MASTER_EN_c_0, DOUTA8 => 
        \DOUTA_1[8]\, DOUTA7 => ELINK_DOUTA_5(7), DOUTA6 => 
        ELINK_DOUTA_5(6), DOUTA5 => ELINK_DOUTA_5(5), DOUTA4 => 
        ELINK_DOUTA_5(4), DOUTA3 => ELINK_DOUTA_5(3), DOUTA2 => 
        ELINK_DOUTA_5(2), DOUTA1 => ELINK_DOUTA_5(1), DOUTA0 => 
        ELINK_DOUTA_5(0), DOUTB8 => \DOUTB_1[8]\, DOUTB7 => 
        PATT_ELK_DAT_5(7), DOUTB6 => PATT_ELK_DAT_5(6), DOUTB5
         => PATT_ELK_DAT_5(5), DOUTB4 => PATT_ELK_DAT_5(4), 
        DOUTB3 => PATT_ELK_DAT_5(3), DOUTB2 => PATT_ELK_DAT_5(2), 
        DOUTB1 => PATT_ELK_DAT_5(1), DOUTB0 => PATT_ELK_DAT_5(0));
    
    VCC_i : VCC
      port map(Y => DPRT_512X9_SRAM_5_VCC);
    
    GND_i : GND
      port map(Y => DPRT_512X9_SRAM_5_GND);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity USB_INTERFACE is

    port( OP_MODE_c_6_0          : out   std_logic;
          OP_MODE_c_5_0          : out   std_logic;
          OP_MODE_c_4_0          : out   std_logic;
          OP_MODE_c_3_0          : out   std_logic;
          OP_MODE_c_2_0          : out   std_logic;
          OP_MODE_c_1_0          : out   std_logic;
          OP_MODE_c_0_0          : out   std_logic;
          OP_MODE_c_1_d0         : out   std_logic;
          OP_MODE_c_5_d0         : out   std_logic;
          OP_MODE_c_4_d0         : out   std_logic;
          OP_MODE_c_0_d0         : out   std_logic;
          OP_MODE_0_0            : out   std_logic;
          OP_MODE_0_4            : out   std_logic;
          ELKS_STOP_ADDR         : out   std_logic_vector(7 downto 0);
          ELKS_STRT_ADDR         : out   std_logic_vector(7 downto 0);
          TFC_STOP_ADDR_0        : out   std_logic_vector(7 downto 0);
          TFC_STRT_ADDR_0        : out   std_logic_vector(7 downto 0);
          BIDIR_USB_ADBUS        : inout std_logic_vector(7 downto 0) := (others => 'Z');
          PATT_ELK_DAT_19        : out   std_logic_vector(7 downto 0);
          ELK_RX_SER_WORD_19     : in    std_logic_vector(7 downto 0);
          PATT_ELK_DAT_18        : out   std_logic_vector(7 downto 0);
          ELK_RX_SER_WORD_18     : in    std_logic_vector(7 downto 0);
          PATT_ELK_DAT_17        : out   std_logic_vector(7 downto 0);
          ELK_RX_SER_WORD_17     : in    std_logic_vector(7 downto 0);
          PATT_ELK_DAT_16        : out   std_logic_vector(7 downto 0);
          ELK_RX_SER_WORD_16     : in    std_logic_vector(7 downto 0);
          PATT_ELK_DAT_15        : out   std_logic_vector(7 downto 0);
          ELK_RX_SER_WORD_15     : in    std_logic_vector(7 downto 0);
          PATT_ELK_DAT_14        : out   std_logic_vector(7 downto 0);
          ELK_RX_SER_WORD_14     : in    std_logic_vector(7 downto 0);
          PATT_ELK_DAT_13        : out   std_logic_vector(7 downto 0);
          ELK_RX_SER_WORD_13     : in    std_logic_vector(7 downto 0);
          PATT_ELK_DAT_12        : out   std_logic_vector(7 downto 0);
          ELK_RX_SER_WORD_12     : in    std_logic_vector(7 downto 0);
          PATT_ELK_DAT_11        : out   std_logic_vector(7 downto 0);
          ELK_RX_SER_WORD_11     : in    std_logic_vector(7 downto 0);
          PATT_ELK_DAT_10        : out   std_logic_vector(7 downto 0);
          ELK_RX_SER_WORD_10     : in    std_logic_vector(7 downto 0);
          PATT_ELK_DAT_9         : out   std_logic_vector(7 downto 0);
          ELK_RX_SER_WORD_9      : in    std_logic_vector(7 downto 0);
          PATT_ELK_DAT_8         : out   std_logic_vector(7 downto 0);
          ELK_RX_SER_WORD_8      : in    std_logic_vector(7 downto 0);
          PATT_ELK_DAT_7         : out   std_logic_vector(7 downto 0);
          ELK_RX_SER_WORD_7      : in    std_logic_vector(7 downto 0);
          PATT_ELK_DAT_6         : out   std_logic_vector(7 downto 0);
          ELK_RX_SER_WORD_6      : in    std_logic_vector(7 downto 0);
          PATT_ELK_DAT_5         : out   std_logic_vector(7 downto 0);
          ELK_RX_SER_WORD_5      : in    std_logic_vector(7 downto 0);
          PATT_ELK_DAT_4         : out   std_logic_vector(7 downto 0);
          ELK_RX_SER_WORD_4      : in    std_logic_vector(7 downto 0);
          PATT_ELK_DAT_3         : out   std_logic_vector(7 downto 0);
          ELK_RX_SER_WORD_3      : in    std_logic_vector(7 downto 0);
          PATT_ELK_DAT_2         : out   std_logic_vector(7 downto 0);
          ELK_RX_SER_WORD_2      : in    std_logic_vector(7 downto 0);
          PATT_ELK_DAT_1         : out   std_logic_vector(7 downto 0);
          ELKS_ADDRB_0_0         : in    std_logic;
          ELKS_ADDRB_0_2         : in    std_logic;
          ELKS_ADDRB_0_4         : in    std_logic;
          ELK_RX_SER_WORD_1      : in    std_logic_vector(7 downto 0);
          PATT_ELK_DAT_0         : out   std_logic_vector(7 downto 0);
          ELKS_ADDRB             : in    std_logic_vector(7 downto 0);
          ELK_RX_SER_WORD_0      : in    std_logic_vector(7 downto 0);
          PATT_TFC_DAT           : out   std_logic_vector(7 downto 0);
          TFC_ADDRB              : in    std_logic_vector(7 downto 0);
          TFC_RX_SER_WORD        : in    std_logic_vector(7 downto 0);
          P_MASTER_POR_B_c_0_0   : in    std_logic;
          P_MASTER_POR_B_c_1     : in    std_logic;
          P_MASTER_POR_B_c       : in    std_logic;
          P_MASTER_POR_B_c_6     : in    std_logic;
          P_MASTER_POR_B_c_24    : in    std_logic;
          P_MASTER_POR_B_c_3     : in    std_logic;
          P_MASTER_POR_B_c_26    : in    std_logic;
          P_MASTER_POR_B_c_33    : in    std_logic;
          P_MASTER_POR_B_c_22_0  : in    std_logic;
          P_MASTER_POR_B_c_28    : in    std_logic;
          P_MASTER_POR_B_c_23    : in    std_logic;
          P_MASTER_POR_B_c_19    : in    std_logic;
          P_MASTER_POR_B_c_24_0  : in    std_logic;
          P_MASTER_POR_B_c_25    : in    std_logic;
          P_MASTER_POR_B_c_29    : in    std_logic;
          P_MASTER_POR_B_c_30    : in    std_logic;
          P_MASTER_POR_B_c_27    : in    std_logic;
          P_MASTER_POR_B_c_17    : in    std_logic;
          P_MASTER_POR_B_c_32    : in    std_logic;
          P_MASTER_POR_B_c_32_0  : in    std_logic;
          P_MASTER_POR_B_c_21    : in    std_logic;
          P_MASTER_POR_B_c_22    : in    std_logic;
          ELKS_RAM_BLKB_EN       : in    std_logic;
          ELKS_RWB               : in    std_logic;
          TFC_RAM_BLKB_EN        : in    std_logic;
          CLK_40M_GL             : in    std_logic;
          TFC_RWB                : in    std_logic;
          P_USB_MASTER_EN_c_1    : in    std_logic;
          P_USB_MASTER_EN_c_0    : in    std_logic;
          P_USB_MASTER_EN_c_2    : in    std_logic;
          P_USB_MASTER_EN_c_20   : in    std_logic;
          P_USB_MASTER_EN_c_6    : in    std_logic;
          P_USB_MASTER_EN_c_9    : in    std_logic;
          P_USB_MASTER_EN_c_11   : in    std_logic;
          P_USB_MASTER_EN_c_12   : in    std_logic;
          P_USB_MASTER_EN_c_14   : in    std_logic;
          P_USB_MASTER_EN_c_18   : in    std_logic;
          P_USB_MASTER_EN_c_7    : in    std_logic;
          P_USB_MASTER_EN_c_21   : in    std_logic;
          P_USB_MASTER_EN_c_17   : in    std_logic;
          P_USB_MASTER_EN_c_15   : in    std_logic;
          P_USB_MASTER_EN_c_4    : in    std_logic;
          USB_WR_BI              : out   std_logic;
          P_USB_MASTER_EN_c_3    : in    std_logic;
          P_USB_MASTER_EN_c_8    : in    std_logic;
          USB_SIWU_BI            : out   std_logic;
          P_USB_MASTER_EN_c_19   : in    std_logic;
          USB_OE_BI              : out   std_logic;
          USB_RD_BI              : out   std_logic;
          P_USB_MASTER_EN_c_13   : in    std_logic;
          P_USB_MASTER_EN_c_5    : in    std_logic;
          P_USB_MASTER_EN_c_10   : in    std_logic;
          P_USB_MASTER_EN_c_22   : in    std_logic;
          P_USB_TXE_B_c          : in    std_logic;
          P_USB_MASTER_EN_c_16   : in    std_logic;
          P_USB_MASTER_EN_c_22_0 : in    std_logic;
          P_USB_MASTER_EN_c_2_0  : in    std_logic;
          P_USB_MASTER_EN_c_1_0  : in    std_logic;
          P_USB_MASTER_EN_c      : in    std_logic;
          P_USB_RXF_B_c          : in    std_logic;
          CLK60MHZ               : in    std_logic
        );

end USB_INTERFACE;

architecture DEF_ARCH of USB_INTERFACE is 

  component DFN1E0C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component AO1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E0P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XO1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DPRT_512X9_SRAM_0
    port( ELINK_RWA_0         : in    std_logic := 'U';
          ELK_RX_SER_WORD_0   : in    std_logic_vector(7 downto 0) := (others => 'U');
          ELINK_DINA_0        : in    std_logic_vector(7 downto 0) := (others => 'U');
          ELINK_BLKA_0        : in    std_logic := 'U';
          ELKS_ADDRB          : in    std_logic_vector(7 downto 0) := (others => 'U');
          ELINK_ADDRA_0       : in    std_logic_vector(7 downto 0) := (others => 'U');
          PATT_ELK_DAT_0      : out   std_logic_vector(7 downto 0);
          ELINK_DOUTA_0       : out   std_logic_vector(7 downto 0);
          ELKS_RWB            : in    std_logic := 'U';
          P_USB_MASTER_EN_c_0 : in    std_logic := 'U';
          CLK_40M_GL          : in    std_logic := 'U';
          CLK60MHZ            : in    std_logic := 'U';
          ELKS_RAM_BLKB_EN    : in    std_logic := 'U'
        );
  end component;

  component AO1D
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DPRT_512X9_SRAM_13
    port( ELINK_RWA_0         : in    std_logic := 'U';
          ELK_RX_SER_WORD_13  : in    std_logic_vector(7 downto 0) := (others => 'U');
          ELINK_DINA_13       : in    std_logic_vector(7 downto 0) := (others => 'U');
          ELINK_BLKA_0        : in    std_logic := 'U';
          ELKS_ADDRB_0_d0     : in    std_logic := 'U';
          ELKS_ADDRB_1        : in    std_logic := 'U';
          ELKS_ADDRB_3        : in    std_logic := 'U';
          ELKS_ADDRB_5        : in    std_logic := 'U';
          ELKS_ADDRB_7        : in    std_logic := 'U';
          ELKS_ADDRB_0_0      : in    std_logic := 'U';
          ELKS_ADDRB_0_2      : in    std_logic := 'U';
          ELKS_ADDRB_0_4      : in    std_logic := 'U';
          ELINK_ADDRA_13      : in    std_logic_vector(7 downto 0) := (others => 'U');
          PATT_ELK_DAT_13     : out   std_logic_vector(7 downto 0);
          ELINK_DOUTA_13      : out   std_logic_vector(7 downto 0);
          ELKS_RWB            : in    std_logic := 'U';
          P_USB_MASTER_EN_c_0 : in    std_logic := 'U';
          CLK_40M_GL          : in    std_logic := 'U';
          CLK60MHZ            : in    std_logic := 'U';
          ELKS_RAM_BLKB_EN    : in    std_logic := 'U'
        );
  end component;

  component MX2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1E
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component DPRT_512X9_SRAM_12
    port( ELINK_RWA_0         : in    std_logic := 'U';
          ELK_RX_SER_WORD_12  : in    std_logic_vector(7 downto 0) := (others => 'U');
          ELINK_DINA_12       : in    std_logic_vector(7 downto 0) := (others => 'U');
          ELINK_BLKA_0        : in    std_logic := 'U';
          ELKS_ADDRB_0_d0     : in    std_logic := 'U';
          ELKS_ADDRB_1        : in    std_logic := 'U';
          ELKS_ADDRB_3        : in    std_logic := 'U';
          ELKS_ADDRB_5        : in    std_logic := 'U';
          ELKS_ADDRB_7        : in    std_logic := 'U';
          ELKS_ADDRB_0_0      : in    std_logic := 'U';
          ELKS_ADDRB_0_2      : in    std_logic := 'U';
          ELKS_ADDRB_0_4      : in    std_logic := 'U';
          ELINK_ADDRA_12      : in    std_logic_vector(7 downto 0) := (others => 'U');
          PATT_ELK_DAT_12     : out   std_logic_vector(7 downto 0);
          ELINK_DOUTA_12      : out   std_logic_vector(7 downto 0);
          ELKS_RWB            : in    std_logic := 'U';
          P_USB_MASTER_EN_c_0 : in    std_logic := 'U';
          CLK_40M_GL          : in    std_logic := 'U';
          CLK60MHZ            : in    std_logic := 'U';
          ELKS_RAM_BLKB_EN    : in    std_logic := 'U'
        );
  end component;

  component OA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFI1E1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          QN  : out   std_logic
        );
  end component;

  component DPRT_512X9_SRAM_11
    port( ELINK_RWA_0         : in    std_logic := 'U';
          ELK_RX_SER_WORD_11  : in    std_logic_vector(7 downto 0) := (others => 'U');
          ELINK_DINA_11       : in    std_logic_vector(7 downto 0) := (others => 'U');
          ELINK_BLKA_0        : in    std_logic := 'U';
          ELKS_ADDRB_0_d0     : in    std_logic := 'U';
          ELKS_ADDRB_1        : in    std_logic := 'U';
          ELKS_ADDRB_3        : in    std_logic := 'U';
          ELKS_ADDRB_5        : in    std_logic := 'U';
          ELKS_ADDRB_7        : in    std_logic := 'U';
          ELKS_ADDRB_0_0      : in    std_logic := 'U';
          ELKS_ADDRB_0_2      : in    std_logic := 'U';
          ELKS_ADDRB_0_4      : in    std_logic := 'U';
          ELINK_ADDRA_11      : in    std_logic_vector(7 downto 0) := (others => 'U');
          PATT_ELK_DAT_11     : out   std_logic_vector(7 downto 0);
          ELINK_DOUTA_11      : out   std_logic_vector(7 downto 0);
          ELKS_RWB            : in    std_logic := 'U';
          P_USB_MASTER_EN_c_0 : in    std_logic := 'U';
          CLK_40M_GL          : in    std_logic := 'U';
          CLK60MHZ            : in    std_logic := 'U';
          ELKS_RAM_BLKB_EN    : in    std_logic := 'U'
        );
  end component;

  component DPRT_512X9_SRAM_16
    port( ELINK_RWA_0         : in    std_logic := 'U';
          ELK_RX_SER_WORD_16  : in    std_logic_vector(7 downto 0) := (others => 'U');
          ELINK_DINA_16       : in    std_logic_vector(7 downto 0) := (others => 'U');
          ELINK_BLKA_0        : in    std_logic := 'U';
          ELKS_ADDRB_0_d0     : in    std_logic := 'U';
          ELKS_ADDRB_1        : in    std_logic := 'U';
          ELKS_ADDRB_3        : in    std_logic := 'U';
          ELKS_ADDRB_5        : in    std_logic := 'U';
          ELKS_ADDRB_7        : in    std_logic := 'U';
          ELKS_ADDRB_0_0      : in    std_logic := 'U';
          ELKS_ADDRB_0_2      : in    std_logic := 'U';
          ELKS_ADDRB_0_4      : in    std_logic := 'U';
          ELINK_ADDRA_16      : in    std_logic_vector(7 downto 0) := (others => 'U');
          PATT_ELK_DAT_16     : out   std_logic_vector(7 downto 0);
          ELINK_DOUTA_16      : out   std_logic_vector(7 downto 0);
          ELKS_RWB            : in    std_logic := 'U';
          P_USB_MASTER_EN_c_0 : in    std_logic := 'U';
          CLK_40M_GL          : in    std_logic := 'U';
          CLK60MHZ            : in    std_logic := 'U';
          ELKS_RAM_BLKB_EN    : in    std_logic := 'U'
        );
  end component;

  component CLK60M_TO_40M_4_1
    port( ELINKS_STRT_ADDR      : in    std_logic_vector(7 downto 0) := (others => 'U');
          ELKS_STRT_ADDR        : out   std_logic_vector(7 downto 0);
          P_MASTER_POR_B_c_28   : in    std_logic := 'U';
          P_MASTER_POR_B_c_22_0 : in    std_logic := 'U';
          P_MASTER_POR_B_c_33   : in    std_logic := 'U';
          P_MASTER_POR_B_c_21   : in    std_logic := 'U';
          P_MASTER_POR_B_c_32   : in    std_logic := 'U';
          CLK_40M_GL            : in    std_logic := 'U'
        );
  end component;

  component DFN1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component DPRT_512X9_SRAM_3
    port( ELINK_RWA_0         : in    std_logic := 'U';
          ELK_RX_SER_WORD_3   : in    std_logic_vector(7 downto 0) := (others => 'U');
          ELINK_DINA_3        : in    std_logic_vector(7 downto 0) := (others => 'U');
          ELINK_BLKA_0        : in    std_logic := 'U';
          ELKS_ADDRB_0_d0     : in    std_logic := 'U';
          ELKS_ADDRB_1        : in    std_logic := 'U';
          ELKS_ADDRB_3        : in    std_logic := 'U';
          ELKS_ADDRB_5        : in    std_logic := 'U';
          ELKS_ADDRB_7        : in    std_logic := 'U';
          ELKS_ADDRB_0_0      : in    std_logic := 'U';
          ELKS_ADDRB_0_2      : in    std_logic := 'U';
          ELKS_ADDRB_0_4      : in    std_logic := 'U';
          ELINK_ADDRA_3       : in    std_logic_vector(7 downto 0) := (others => 'U');
          PATT_ELK_DAT_3      : out   std_logic_vector(7 downto 0);
          ELINK_DOUTA_3       : out   std_logic_vector(7 downto 0);
          ELKS_RWB            : in    std_logic := 'U';
          P_USB_MASTER_EN_c_0 : in    std_logic := 'U';
          CLK_40M_GL          : in    std_logic := 'U';
          CLK60MHZ            : in    std_logic := 'U';
          ELKS_RAM_BLKB_EN    : in    std_logic := 'U'
        );
  end component;

  component DPRT_512X9_SRAM_2
    port( ELINK_RWA_0         : in    std_logic := 'U';
          ELK_RX_SER_WORD_2   : in    std_logic_vector(7 downto 0) := (others => 'U');
          ELINK_DINA_2        : in    std_logic_vector(7 downto 0) := (others => 'U');
          ELINK_BLKA_0        : in    std_logic := 'U';
          ELKS_ADDRB          : in    std_logic_vector(7 downto 0) := (others => 'U');
          ELINK_ADDRA_2       : in    std_logic_vector(7 downto 0) := (others => 'U');
          PATT_ELK_DAT_2      : out   std_logic_vector(7 downto 0);
          ELINK_DOUTA_2       : out   std_logic_vector(7 downto 0);
          ELKS_RWB            : in    std_logic := 'U';
          P_USB_MASTER_EN_c_0 : in    std_logic := 'U';
          CLK_40M_GL          : in    std_logic := 'U';
          CLK60MHZ            : in    std_logic := 'U';
          ELKS_RAM_BLKB_EN    : in    std_logic := 'U'
        );
  end component;

  component OAI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component DPRT_512X9_SRAM_1
    port( ELINK_RWA_0         : in    std_logic := 'U';
          ELK_RX_SER_WORD_1   : in    std_logic_vector(7 downto 0) := (others => 'U');
          ELINK_DINA_1        : in    std_logic_vector(7 downto 0) := (others => 'U');
          ELINK_BLKA_0        : in    std_logic := 'U';
          ELKS_ADDRB_0_d0     : in    std_logic := 'U';
          ELKS_ADDRB_1        : in    std_logic := 'U';
          ELKS_ADDRB_3        : in    std_logic := 'U';
          ELKS_ADDRB_5        : in    std_logic := 'U';
          ELKS_ADDRB_7        : in    std_logic := 'U';
          ELKS_ADDRB_0_0      : in    std_logic := 'U';
          ELKS_ADDRB_0_2      : in    std_logic := 'U';
          ELKS_ADDRB_0_4      : in    std_logic := 'U';
          ELINK_ADDRA_1       : in    std_logic_vector(7 downto 0) := (others => 'U');
          PATT_ELK_DAT_1      : out   std_logic_vector(7 downto 0);
          ELINK_DOUTA_1       : out   std_logic_vector(7 downto 0);
          ELKS_RWB            : in    std_logic := 'U';
          P_USB_MASTER_EN_c_0 : in    std_logic := 'U';
          CLK_40M_GL          : in    std_logic := 'U';
          CLK60MHZ            : in    std_logic := 'U';
          ELKS_RAM_BLKB_EN    : in    std_logic := 'U'
        );
  end component;

  component DPRT_512X9_SRAM_6
    port( ELINK_RWA_0         : in    std_logic := 'U';
          ELK_RX_SER_WORD_6   : in    std_logic_vector(7 downto 0) := (others => 'U');
          ELINK_DINA_6        : in    std_logic_vector(7 downto 0) := (others => 'U');
          ELINK_BLKA_0        : in    std_logic := 'U';
          ELKS_ADDRB_0_d0     : in    std_logic := 'U';
          ELKS_ADDRB_1        : in    std_logic := 'U';
          ELKS_ADDRB_3        : in    std_logic := 'U';
          ELKS_ADDRB_5        : in    std_logic := 'U';
          ELKS_ADDRB_7        : in    std_logic := 'U';
          ELKS_ADDRB_0_0      : in    std_logic := 'U';
          ELKS_ADDRB_0_2      : in    std_logic := 'U';
          ELKS_ADDRB_0_4      : in    std_logic := 'U';
          ELINK_ADDRA_6       : in    std_logic_vector(7 downto 0) := (others => 'U');
          PATT_ELK_DAT_6      : out   std_logic_vector(7 downto 0);
          ELINK_DOUTA_6       : out   std_logic_vector(7 downto 0);
          ELKS_RWB            : in    std_logic := 'U';
          P_USB_MASTER_EN_c_0 : in    std_logic := 'U';
          CLK_40M_GL          : in    std_logic := 'U';
          CLK60MHZ            : in    std_logic := 'U';
          ELKS_RAM_BLKB_EN    : in    std_logic := 'U'
        );
  end component;

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CLK60M_TO_40M_0
    port( OP_MODE              : inout   std_logic_vector(7 downto 0);
          OP_MODE_0_0          : in    std_logic := 'U';
          OP_MODE_0_4          : in    std_logic := 'U';
          OP_MODE_c_1_d0       : out   std_logic;
          OP_MODE_c_5_d0       : out   std_logic;
          OP_MODE_c_4_d0       : out   std_logic;
          OP_MODE_c_0_d0       : out   std_logic;
          OP_MODE_c_0_0        : out   std_logic;
          OP_MODE_c_1_0        : out   std_logic;
          OP_MODE_c_2_0        : out   std_logic;
          OP_MODE_c_3_0        : out   std_logic;
          OP_MODE_c_4_0        : out   std_logic;
          OP_MODE_c_5_0        : out   std_logic;
          OP_MODE_c_6_0        : out   std_logic;
          P_MASTER_POR_B_c_25  : in    std_logic := 'U';
          P_MASTER_POR_B_c_24  : in    std_logic := 'U';
          P_MASTER_POR_B_c_23  : in    std_logic := 'U';
          P_MASTER_POR_B_c_6   : in    std_logic := 'U';
          P_MASTER_POR_B_c     : in    std_logic := 'U';
          P_MASTER_POR_B_c_1   : in    std_logic := 'U';
          P_MASTER_POR_B_c_0_0 : in    std_logic := 'U';
          CLK_40M_GL           : in    std_logic := 'U'
        );
  end component;

  component BIDIR_LVTTL
    port( WR_USB_ADBUS    : in    std_logic_vector(7 downto 0) := (others => 'U');
          N_RD_USB_ADBUS  : out   std_logic_vector(7 downto 0);
          BIDIR_USB_ADBUS : inout   std_logic_vector(7 downto 0);
          TrienAux        : in    std_logic := 'U'
        );
  end component;

  component DPRT_512X9_SRAM_14
    port( ELINK_RWA_0         : in    std_logic := 'U';
          ELK_RX_SER_WORD_14  : in    std_logic_vector(7 downto 0) := (others => 'U');
          ELINK_DINA_14       : in    std_logic_vector(7 downto 0) := (others => 'U');
          ELINK_BLKA_0        : in    std_logic := 'U';
          ELKS_ADDRB_0_d0     : in    std_logic := 'U';
          ELKS_ADDRB_1        : in    std_logic := 'U';
          ELKS_ADDRB_3        : in    std_logic := 'U';
          ELKS_ADDRB_5        : in    std_logic := 'U';
          ELKS_ADDRB_7        : in    std_logic := 'U';
          ELKS_ADDRB_0_0      : in    std_logic := 'U';
          ELKS_ADDRB_0_2      : in    std_logic := 'U';
          ELKS_ADDRB_0_4      : in    std_logic := 'U';
          ELINK_ADDRA_14      : in    std_logic_vector(7 downto 0) := (others => 'U');
          PATT_ELK_DAT_14     : out   std_logic_vector(7 downto 0);
          ELINK_DOUTA_14      : out   std_logic_vector(7 downto 0);
          ELKS_RWB            : in    std_logic := 'U';
          P_USB_MASTER_EN_c_0 : in    std_logic := 'U';
          CLK_40M_GL          : in    std_logic := 'U';
          CLK60MHZ            : in    std_logic := 'U';
          ELKS_RAM_BLKB_EN    : in    std_logic := 'U'
        );
  end component;

  component DPRT_512X9_SRAM_17
    port( ELINK_RWA_0         : in    std_logic := 'U';
          ELK_RX_SER_WORD_17  : in    std_logic_vector(7 downto 0) := (others => 'U');
          ELINK_DINA_17       : in    std_logic_vector(7 downto 0) := (others => 'U');
          ELINK_BLKA_0        : in    std_logic := 'U';
          ELKS_ADDRB          : in    std_logic_vector(7 downto 0) := (others => 'U');
          ELINK_ADDRA_17      : in    std_logic_vector(7 downto 0) := (others => 'U');
          PATT_ELK_DAT_17     : out   std_logic_vector(7 downto 0);
          ELINK_DOUTA_17      : out   std_logic_vector(7 downto 0);
          ELKS_RWB            : in    std_logic := 'U';
          P_USB_MASTER_EN_c_0 : in    std_logic := 'U';
          CLK_40M_GL          : in    std_logic := 'U';
          CLK60MHZ            : in    std_logic := 'U';
          ELKS_RAM_BLKB_EN    : in    std_logic := 'U'
        );
  end component;

  component CLK60M_TO_40M_4_2
    port( ELINKS_STOP_ADDR    : in    std_logic_vector(7 downto 0) := (others => 'U');
          ELKS_STOP_ADDR      : out   std_logic_vector(7 downto 0);
          P_MASTER_POR_B_c_26 : in    std_logic := 'U';
          P_MASTER_POR_B_c_30 : in    std_logic := 'U';
          P_MASTER_POR_B_c_3  : in    std_logic := 'U';
          P_MASTER_POR_B_c_25 : in    std_logic := 'U';
          CLK_40M_GL          : in    std_logic := 'U'
        );
  end component;

  component CLK60M_TO_40M_4_0
    port( TFC_STOP_ADDR_0       : in    std_logic_vector(7 downto 0) := (others => 'U');
          TFC_STOP_ADDR         : out   std_logic_vector(7 downto 0);
          P_MASTER_POR_B_c_30   : in    std_logic := 'U';
          P_MASTER_POR_B_c_29   : in    std_logic := 'U';
          P_MASTER_POR_B_c_25   : in    std_logic := 'U';
          P_MASTER_POR_B_c_24_0 : in    std_logic := 'U';
          P_MASTER_POR_B_c_19   : in    std_logic := 'U';
          P_MASTER_POR_B_c_23   : in    std_logic := 'U';
          CLK_40M_GL            : in    std_logic := 'U'
        );
  end component;

  component DPRT_512X9_SRAM_4
    port( ELINK_RWA_0         : in    std_logic := 'U';
          ELK_RX_SER_WORD_4   : in    std_logic_vector(7 downto 0) := (others => 'U');
          ELINK_DINA_4        : in    std_logic_vector(7 downto 0) := (others => 'U');
          ELINK_BLKA_0        : in    std_logic := 'U';
          ELKS_ADDRB          : in    std_logic_vector(7 downto 0) := (others => 'U');
          ELINK_ADDRA_4       : in    std_logic_vector(7 downto 0) := (others => 'U');
          PATT_ELK_DAT_4      : out   std_logic_vector(7 downto 0);
          ELINK_DOUTA_4       : out   std_logic_vector(7 downto 0);
          ELKS_RWB            : in    std_logic := 'U';
          P_USB_MASTER_EN_c_0 : in    std_logic := 'U';
          CLK_40M_GL          : in    std_logic := 'U';
          CLK60MHZ            : in    std_logic := 'U';
          ELKS_RAM_BLKB_EN    : in    std_logic := 'U'
        );
  end component;

  component DPRT_512X9_SRAM_19
    port( ELINK_RWA_0         : in    std_logic := 'U';
          ELK_RX_SER_WORD_19  : in    std_logic_vector(7 downto 0) := (others => 'U');
          ELINK_DINA_19       : in    std_logic_vector(7 downto 0) := (others => 'U');
          ELINK_BLKA_0        : in    std_logic := 'U';
          ELKS_ADDRB          : in    std_logic_vector(7 downto 0) := (others => 'U');
          ELINK_ADDRA_19      : in    std_logic_vector(7 downto 0) := (others => 'U');
          PATT_ELK_DAT_19     : out   std_logic_vector(7 downto 0);
          ELINK_DOUTA_19      : out   std_logic_vector(7 downto 0);
          ELKS_RWB            : in    std_logic := 'U';
          P_USB_MASTER_EN_c_0 : in    std_logic := 'U';
          CLK_40M_GL          : in    std_logic := 'U';
          CLK60MHZ            : in    std_logic := 'U';
          ELKS_RAM_BLKB_EN    : in    std_logic := 'U'
        );
  end component;

  component DPRT_512X9_SRAM_7
    port( ELINK_RWA_0         : in    std_logic := 'U';
          ELK_RX_SER_WORD_7   : in    std_logic_vector(7 downto 0) := (others => 'U');
          ELINK_DINA_7        : in    std_logic_vector(7 downto 0) := (others => 'U');
          ELINK_BLKA_0        : in    std_logic := 'U';
          ELKS_ADDRB_0_d0     : in    std_logic := 'U';
          ELKS_ADDRB_1        : in    std_logic := 'U';
          ELKS_ADDRB_3        : in    std_logic := 'U';
          ELKS_ADDRB_5        : in    std_logic := 'U';
          ELKS_ADDRB_7        : in    std_logic := 'U';
          ELKS_ADDRB_0_0      : in    std_logic := 'U';
          ELKS_ADDRB_0_2      : in    std_logic := 'U';
          ELKS_ADDRB_0_4      : in    std_logic := 'U';
          ELINK_ADDRA_7       : in    std_logic_vector(7 downto 0) := (others => 'U');
          PATT_ELK_DAT_7      : out   std_logic_vector(7 downto 0);
          ELINK_DOUTA_7       : out   std_logic_vector(7 downto 0);
          ELKS_RWB            : in    std_logic := 'U';
          P_USB_MASTER_EN_c_0 : in    std_logic := 'U';
          CLK_40M_GL          : in    std_logic := 'U';
          CLK60MHZ            : in    std_logic := 'U';
          ELKS_RAM_BLKB_EN    : in    std_logic := 'U'
        );
  end component;

  component CLK60M_TO_40M_4
    port( TFC_STRT_ADDR_0       : in    std_logic_vector(7 downto 0) := (others => 'U');
          TFC_STRT_ADDR         : out   std_logic_vector(7 downto 0);
          P_MASTER_POR_B_c_22   : in    std_logic := 'U';
          P_MASTER_POR_B_c_21   : in    std_logic := 'U';
          P_MASTER_POR_B_c_32_0 : in    std_logic := 'U';
          P_MASTER_POR_B_c_32   : in    std_logic := 'U';
          P_MASTER_POR_B_c_17   : in    std_logic := 'U';
          P_MASTER_POR_B_c_27   : in    std_logic := 'U';
          CLK_40M_GL            : in    std_logic := 'U'
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DPRT_512X9_SRAM_9
    port( ELINK_RWA_0         : in    std_logic := 'U';
          ELK_RX_SER_WORD_9   : in    std_logic_vector(7 downto 0) := (others => 'U');
          ELINK_DINA_9        : in    std_logic_vector(7 downto 0) := (others => 'U');
          ELINK_BLKA_0        : in    std_logic := 'U';
          ELKS_ADDRB          : in    std_logic_vector(7 downto 0) := (others => 'U');
          ELINK_ADDRA_9       : in    std_logic_vector(7 downto 0) := (others => 'U');
          PATT_ELK_DAT_9      : out   std_logic_vector(7 downto 0);
          ELINK_DOUTA_9       : out   std_logic_vector(7 downto 0);
          ELKS_RWB            : in    std_logic := 'U';
          P_USB_MASTER_EN_c_0 : in    std_logic := 'U';
          CLK_40M_GL          : in    std_logic := 'U';
          CLK60MHZ            : in    std_logic := 'U';
          ELKS_RAM_BLKB_EN    : in    std_logic := 'U'
        );
  end component;

  component DPRT_512X9_SRAM_18
    port( ELINK_RWA_0         : in    std_logic := 'U';
          ELK_RX_SER_WORD_18  : in    std_logic_vector(7 downto 0) := (others => 'U');
          ELINK_DINA_18       : in    std_logic_vector(7 downto 0) := (others => 'U');
          ELINK_BLKA_0        : in    std_logic := 'U';
          ELKS_ADDRB_0_d0     : in    std_logic := 'U';
          ELKS_ADDRB_1        : in    std_logic := 'U';
          ELKS_ADDRB_3        : in    std_logic := 'U';
          ELKS_ADDRB_5        : in    std_logic := 'U';
          ELKS_ADDRB_7        : in    std_logic := 'U';
          ELKS_ADDRB_0_0      : in    std_logic := 'U';
          ELKS_ADDRB_0_2      : in    std_logic := 'U';
          ELKS_ADDRB_0_4      : in    std_logic := 'U';
          ELINK_ADDRA_18      : in    std_logic_vector(7 downto 0) := (others => 'U');
          PATT_ELK_DAT_18     : out   std_logic_vector(7 downto 0);
          ELINK_DOUTA_18      : out   std_logic_vector(7 downto 0);
          ELKS_RWB            : in    std_logic := 'U';
          P_USB_MASTER_EN_c_0 : in    std_logic := 'U';
          CLK_40M_GL          : in    std_logic := 'U';
          CLK60MHZ            : in    std_logic := 'U';
          ELKS_RAM_BLKB_EN    : in    std_logic := 'U'
        );
  end component;

  component DPRT_512X9_SRAM_15
    port( ELINK_RWA_0         : in    std_logic := 'U';
          ELK_RX_SER_WORD_15  : in    std_logic_vector(7 downto 0) := (others => 'U');
          ELINK_DINA_15       : in    std_logic_vector(7 downto 0) := (others => 'U');
          ELINK_BLKA_0        : in    std_logic := 'U';
          ELKS_ADDRB          : in    std_logic_vector(7 downto 0) := (others => 'U');
          ELINK_ADDRA_15      : in    std_logic_vector(7 downto 0) := (others => 'U');
          PATT_ELK_DAT_15     : out   std_logic_vector(7 downto 0);
          ELINK_DOUTA_15      : out   std_logic_vector(7 downto 0);
          ELKS_RWB            : in    std_logic := 'U';
          P_USB_MASTER_EN_c_0 : in    std_logic := 'U';
          CLK_40M_GL          : in    std_logic := 'U';
          CLK60MHZ            : in    std_logic := 'U';
          ELKS_RAM_BLKB_EN    : in    std_logic := 'U'
        );
  end component;

  component XNOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component DPRT_512X9_SRAM
    port( TFC_RX_SER_WORD     : in    std_logic_vector(7 downto 0) := (others => 'U');
          TFC_DINA            : in    std_logic_vector(7 downto 0) := (others => 'U');
          TFC_ADDRB           : in    std_logic_vector(7 downto 0) := (others => 'U');
          TFC_ADDRA           : in    std_logic_vector(7 downto 0) := (others => 'U');
          PATT_TFC_DAT        : out   std_logic_vector(7 downto 0);
          TFC_DOUTA           : out   std_logic_vector(7 downto 0);
          TFC_RWB             : in    std_logic := 'U';
          TFC_RWA             : in    std_logic := 'U';
          P_USB_MASTER_EN_c_0 : in    std_logic := 'U';
          CLK_40M_GL          : in    std_logic := 'U';
          CLK60MHZ            : in    std_logic := 'U';
          TFC_RAM_BLKB_EN     : in    std_logic := 'U';
          TFC_BLKA            : in    std_logic := 'U'
        );
  end component;

  component DPRT_512X9_SRAM_10
    port( ELINK_RWA_0         : in    std_logic := 'U';
          ELK_RX_SER_WORD_10  : in    std_logic_vector(7 downto 0) := (others => 'U');
          ELINK_DINA_10       : in    std_logic_vector(7 downto 0) := (others => 'U');
          ELINK_BLKA_0        : in    std_logic := 'U';
          ELKS_ADDRB_0_d0     : in    std_logic := 'U';
          ELKS_ADDRB_1        : in    std_logic := 'U';
          ELKS_ADDRB_3        : in    std_logic := 'U';
          ELKS_ADDRB_5        : in    std_logic := 'U';
          ELKS_ADDRB_7        : in    std_logic := 'U';
          ELKS_ADDRB_0_0      : in    std_logic := 'U';
          ELKS_ADDRB_0_2      : in    std_logic := 'U';
          ELKS_ADDRB_0_4      : in    std_logic := 'U';
          ELINK_ADDRA_10      : in    std_logic_vector(7 downto 0) := (others => 'U');
          PATT_ELK_DAT_10     : out   std_logic_vector(7 downto 0);
          ELINK_DOUTA_10      : out   std_logic_vector(7 downto 0);
          ELKS_RWB            : in    std_logic := 'U';
          P_USB_MASTER_EN_c_0 : in    std_logic := 'U';
          CLK_40M_GL          : in    std_logic := 'U';
          CLK60MHZ            : in    std_logic := 'U';
          ELKS_RAM_BLKB_EN    : in    std_logic := 'U'
        );
  end component;

  component DPRT_512X9_SRAM_8
    port( ELINK_RWA_0         : in    std_logic := 'U';
          ELK_RX_SER_WORD_8   : in    std_logic_vector(7 downto 0) := (others => 'U');
          ELINK_DINA_8        : in    std_logic_vector(7 downto 0) := (others => 'U');
          ELINK_BLKA_0        : in    std_logic := 'U';
          ELKS_ADDRB_0_d0     : in    std_logic := 'U';
          ELKS_ADDRB_1        : in    std_logic := 'U';
          ELKS_ADDRB_3        : in    std_logic := 'U';
          ELKS_ADDRB_5        : in    std_logic := 'U';
          ELKS_ADDRB_7        : in    std_logic := 'U';
          ELKS_ADDRB_0_0      : in    std_logic := 'U';
          ELKS_ADDRB_0_2      : in    std_logic := 'U';
          ELKS_ADDRB_0_4      : in    std_logic := 'U';
          ELINK_ADDRA_8       : in    std_logic_vector(7 downto 0) := (others => 'U');
          PATT_ELK_DAT_8      : out   std_logic_vector(7 downto 0);
          ELINK_DOUTA_8       : out   std_logic_vector(7 downto 0);
          ELKS_RWB            : in    std_logic := 'U';
          P_USB_MASTER_EN_c_0 : in    std_logic := 'U';
          CLK_40M_GL          : in    std_logic := 'U';
          CLK60MHZ            : in    std_logic := 'U';
          ELKS_RAM_BLKB_EN    : in    std_logic := 'U'
        );
  end component;

  component DPRT_512X9_SRAM_5
    port( ELINK_RWA_0         : in    std_logic := 'U';
          ELK_RX_SER_WORD_5   : in    std_logic_vector(7 downto 0) := (others => 'U');
          ELINK_DINA_5        : in    std_logic_vector(7 downto 0) := (others => 'U');
          ELINK_BLKA_0        : in    std_logic := 'U';
          ELKS_ADDRB_0_d0     : in    std_logic := 'U';
          ELKS_ADDRB_1        : in    std_logic := 'U';
          ELKS_ADDRB_3        : in    std_logic := 'U';
          ELKS_ADDRB_5        : in    std_logic := 'U';
          ELKS_ADDRB_7        : in    std_logic := 'U';
          ELKS_ADDRB_0_0      : in    std_logic := 'U';
          ELKS_ADDRB_0_2      : in    std_logic := 'U';
          ELKS_ADDRB_0_4      : in    std_logic := 'U';
          ELINK_ADDRA_5       : in    std_logic_vector(7 downto 0) := (others => 'U');
          PATT_ELK_DAT_5      : out   std_logic_vector(7 downto 0);
          ELINK_DOUTA_5       : out   std_logic_vector(7 downto 0);
          ELKS_RWB            : in    std_logic := 'U';
          P_USB_MASTER_EN_c_0 : in    std_logic := 'U';
          CLK_40M_GL          : in    std_logic := 'U';
          CLK60MHZ            : in    std_logic := 'U';
          ELKS_RAM_BLKB_EN    : in    std_logic := 'U'
        );
  end component;

  component XA1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \USB_RXF_B_0\, \SM_BANK_SEL_0[20]_net_1\, 
        un1_N_ELK_N_ACTIVE_2_sqmuxa, un1_REG_STATE_30, 
        \SM_BANK_SEL_0[21]_net_1\, N_1671, \REG_STATE_0[0]_net_1\, 
        \REG_STATE_ns_i_i_a2_0_RNIN0TJ41[0]_net_1\, 
        \REG_STATE_0[1]_net_1\, \USB_TXE_B_RNI75TNL2\, 
        \REG_STATE_0[2]_net_1\, \REG_STATE_RNIVPG2K2[2]_net_1\, 
        \REG_STATE_0[3]_net_1\, \REG_STATE_0_RNIGPV6T1[0]_net_1\, 
        \REG_STATE_0[4]_net_1\, \REG_STATE_RNIMO53U3[2]_net_1\, 
        \REG_STATE_0[5]_net_1\, \USB_TXE_B_RNIV2O4Q\, N_675_0, 
        N_1710_i_0, N_1691, N_312_0, \REG_STATE_d_0[30]\, 
        N_1359_2, N_1352_1, N_1763, N_290, 
        \RD_USB_ADBUS[4]_net_1\, N_1717, 
        \WR_XFER_TYPE_RNO[2]_net_1\, N_1824, N_1823, N_1822, 
        \WR_XFER_TYPE_RNO[3]_net_1\, N_1826, N_1825, 
        \WR_XFER_TYPE_RNO[4]_net_1\, N_1716, N_1827, N_1892, 
        N_1882, \RD_USB_ADBUS[3]_net_1\, N_1846, N_1902, 
        \RD_USB_ADBUS[2]_net_1\, N_1839, N_1351_4, N_1837, N_1836, 
        \RD_USB_ADBUS[5]_net_1\, \WR_XFER_TYPE[4]_net_1\, 
        \WR_XFER_TYPE[3]_net_1\, N_1881, \WR_XFER_TYPE[2]_net_1\, 
        N_1832, N_1842, N_1697, N_293, N_1702, 
        \RD_USB_ADBUS[7]_net_1\, N_1690_i, \REG_STATE[4]_net_1\, 
        \REG_STATE[1]_net_1\, \REG_STATE[3]_net_1\, N_2497, 
        \REG_STATE[0]_net_1\, \REG_STATE[2]_net_1\, N_1694, 
        N_1695, \WR_XFER_TYPE_RNO[5]_net_1\, 
        \WR_XFER_TYPE[5]_net_1\, N_1829, N_1700, N_1845, N_1352_4, 
        N_1847, TrienAux, un1_REG_STATE_23, N_251, 
        \SM_BANK_SEL[20]_net_1\, \ELK_N_ACTIVE\, N_1705, N_275, 
        N_444, N_443, N_1782, N_1782_1, N_1726, un1_REG_STATE_4, 
        N_1781, N_421, \REG_STATE_ns_i_i_a2_0_2[0]_net_1\, 
        N_244_1, \REG_STATE_ns_i_i_o2_6_1[0]_net_1\, N_78, N_312, 
        N_1566_i_i_0, N_1562_i, un1_REG_STATE_2_i_0, 
        un1_REG_STATE_4_0_a2_1, \REG_STATE_ns_i_a4_1_0[4]_net_1\, 
        N_2606, N_379, \TFC_STOP_ADDR_m[6]\, 
        \TFC_STOP_ADDR[6]_net_1\, N_1501, \TFC_STOP_ADDR_m[4]\, 
        \TFC_STOP_ADDR[4]_net_1\, \TFC_STOP_ADDR_m[2]\, 
        \TFC_STOP_ADDR[2]_net_1\, \TFC_STOP_ADDR_m[0]\, 
        \TFC_STOP_ADDR[0]_net_1\, N_429, N_1704, 
        \N_WR_USB_ADBUS_0_iv_0[0]_net_1\, 
        \N_WR_USB_ADBUS_0_iv_0[6]_net_1\, 
        \N_WR_USB_ADBUS_0_iv_0[2]_net_1\, 
        \N_WR_USB_ADBUS_0_iv_0[4]_net_1\, N_414_i, 
        \REG_STATE_ns_i_i_a2_0_1[0]\, N_487, 
        \REG_STATE_ns_i_i_o2_6_0[0]\, 
        \un1_N_WR_USB_ADBUS_0_sqmuxa_i_0\, \USB_TXE_B\, 
        \REG_STATE_ns_i_8_tz_1[4]_net_1\, 
        \REG_STATE_ns_i_8_tz_0[4]_net_1\, 
        \REG_STATE_ns_i_a4_2_0[4]\, \REG_STATE_ns_i_a4_5_1[4]\, 
        \REG_STATE_s23_i_2\, REG_STATE_s23_i_1, REG_STATE_s23_i_0, 
        N_243, N_261, \N_TFC_ADDRA_0_o2_0[7]\, 
        \REG_STATE_ns_i_i_2[0]\, N_358, N_357, 
        \REG_STATE_ns_i_i_0[0]\, N_2576, N_1374, 
        \REG_STATE_ns_i_4[4]\, \REG_STATE_ns_i_a4_0[4]\, 
        \REG_STATE_ns_i_a4_9_1[4]\, N_2597, \REG_STATE_ns_i_3[4]\, 
        N_264, \REG_STATE_ns_i_1[4]\, \REG_STATE_ns_i_8[4]\, 
        N_2570, N_1877_1, N_2566, \N_WR_USB_ADBUS_0_iv_25[7]\, 
        \N_WR_USB_ADBUS_0_iv_14[7]\, \N_WR_USB_ADBUS_0_iv_13[7]\, 
        \N_WR_USB_ADBUS_0_iv_22[7]\, \N_WR_USB_ADBUS_0_iv_24[7]\, 
        \N_WR_USB_ADBUS_0_iv_10[7]\, \N_WR_USB_ADBUS_0_iv_9[7]\, 
        \N_WR_USB_ADBUS_0_iv_20[7]\, \N_WR_USB_ADBUS_0_iv_23[7]\, 
        \N_WR_USB_ADBUS_0_iv_6[7]\, \ELINK_DOUTA_14_m[7]\, 
        \N_WR_USB_ADBUS_0_iv_18[7]\, \ELINK_DOUTA_11_m[7]\, 
        \ELINK_DOUTA_10_m[7]\, \N_WR_USB_ADBUS_0_iv_16[7]\, 
        \ELINK_DOUTA_3_m[7]\, \ELINK_DOUTA_18_m[7]\, 
        \N_WR_USB_ADBUS_0_iv_12[7]\, \TFC_DOUTA_m[7]\, 
        \ELINK_DOUTA_19_m[7]\, \N_WR_USB_ADBUS_0_iv_8[7]\, 
        \ELINK_DOUTA_12[7]\, un1_SM_BANK_SEL_33, 
        \ELINK_DOUTA_13_m[7]\, \ELINK_DOUTA_7[7]\, 
        un1_SM_BANK_SEL_37, \ELINK_DOUTA_9_m[7]\, 
        \ELINK_DOUTA_6[7]\, un1_SM_BANK_SEL_30, 
        \ELINK_DOUTA_8_m[7]\, \ELINK_DOUTA_4[7]\, 
        un1_SM_BANK_SEL_28, \ELINK_DOUTA_5_m[7]\, 
        \ELINK_DOUTA_17[7]\, un1_SM_BANK_SEL_40, 
        \ELINK_DOUTA_2_m[7]\, \ELINK_DOUTA_16[7]\, 
        un1_SM_BANK_SEL_39, \ELINK_DOUTA_1_m[7]\, 
        \ELINK_DOUTA_15[7]\, un1_SM_BANK_SEL_24, 
        \ELINK_DOUTA_0_m[7]\, \N_WR_USB_ADBUS_0_iv_3[7]\, 
        \N_WR_USB_ADBUS_0_iv_2[7]\, \N_WR_USB_ADBUS_0_iv_4[7]\, 
        \CHKSUM[7]_net_1\, \N_WR_USB_ADBUS_0_iv_1[7]\, N_1497, 
        \TFC_STRT_ADDR[7]_net_1\, \ELINKS_STOP_ADDR_m[7]\, 
        \WR_XFER_TYPE[7]_net_1\, N_398, 
        \N_WR_USB_ADBUS_0_iv_0[7]\, N_1499, 
        \ELINKS_STRT_ADDR[7]_net_1\, N_1569, 
        \TFC_STOP_ADDR[7]_net_1\, \OP_MODE_m[7]\, 
        \N_WR_USB_ADBUS_0_iv_25[5]\, \N_WR_USB_ADBUS_0_iv_14[5]\, 
        \N_WR_USB_ADBUS_0_iv_13[5]\, \N_WR_USB_ADBUS_0_iv_22[5]\, 
        \N_WR_USB_ADBUS_0_iv_24[5]\, \N_WR_USB_ADBUS_0_iv_10[5]\, 
        \N_WR_USB_ADBUS_0_iv_9[5]\, \N_WR_USB_ADBUS_0_iv_20[5]\, 
        \N_WR_USB_ADBUS_0_iv_23[5]\, \N_WR_USB_ADBUS_0_iv_6[5]\, 
        \ELINK_DOUTA_14_m[5]\, \N_WR_USB_ADBUS_0_iv_18[5]\, 
        \ELINK_DOUTA_11_m[5]\, \ELINK_DOUTA_10_m[5]\, 
        \N_WR_USB_ADBUS_0_iv_16[5]\, \ELINK_DOUTA_3_m[5]\, 
        \ELINK_DOUTA_18_m[5]\, \N_WR_USB_ADBUS_0_iv_12[5]\, 
        \TFC_DOUTA_m[5]\, \ELINK_DOUTA_19_m[5]\, 
        \N_WR_USB_ADBUS_0_iv_8[5]\, \ELINK_DOUTA_12[5]\, 
        \ELINK_DOUTA_13_m[5]\, \ELINK_DOUTA_7[5]\, 
        \ELINK_DOUTA_9_m[5]\, \ELINK_DOUTA_6_m[5]\, 
        \ELINK_DOUTA_8_m[5]\, \ELINK_DOUTA_4[5]\, 
        \ELINK_DOUTA_5_m[5]\, \ELINK_DOUTA_17[5]\, 
        \ELINK_DOUTA_2_m[5]\, \ELINK_DOUTA_16[5]\, 
        \ELINK_DOUTA_1_m[5]\, \ELINK_DOUTA_15[5]\, 
        \ELINK_DOUTA_0_m[5]\, \N_WR_USB_ADBUS_0_iv_3[5]\, 
        \N_WR_USB_ADBUS_0_iv_2[5]\, \N_WR_USB_ADBUS_0_iv_4[5]\, 
        \ELINKS_STRT_ADDR_m[5]\, \CHKSUM_m[5]\, 
        \TFC_STRT_ADDR[5]_net_1\, \ELINKS_STOP_ADDR_m[5]\, 
        \OP_MODE_m[5]\, \TFC_STOP_ADDR_m[5]\, \WR_XFER_TYPE_m[5]\, 
        \N_WR_USB_ADBUS_0_iv_25[0]\, \N_WR_USB_ADBUS_0_iv_14[0]\, 
        \N_WR_USB_ADBUS_0_iv_13[0]\, \N_WR_USB_ADBUS_0_iv_22[0]\, 
        \N_WR_USB_ADBUS_0_iv_24[0]\, \N_WR_USB_ADBUS_0_iv_10[0]\, 
        \N_WR_USB_ADBUS_0_iv_9[0]\, \N_WR_USB_ADBUS_0_iv_20[0]\, 
        \N_WR_USB_ADBUS_0_iv_23[0]\, \N_WR_USB_ADBUS_0_iv_8[0]\, 
        \N_WR_USB_ADBUS_0_iv_7[0]\, \N_WR_USB_ADBUS_0_iv_17[0]\, 
        \ELINK_DOUTA_17_m[0]\, \ELINK_DOUTA_1_m[0]\, 
        \N_WR_USB_ADBUS_0_iv_16[0]\, \ELINK_DOUTA_13_m[0]\, 
        \ELINK_DOUTA_12_m[0]\, \N_WR_USB_ADBUS_0_iv_12[0]\, 
        \N_WR_USB_ADBUS_0_iv_5[0]\, \N_WR_USB_ADBUS_0_iv_4[0]\, 
        \ELINK_DOUTA_3_m[0]\, \ELINK_DOUTA_2[0]\, 
        un1_SM_BANK_SEL_32, \ELINK_DOUTA_18_m[0]\, 
        \ELINK_DOUTA_0[0]\, un1_SM_BANK_SEL_31, 
        \ELINK_DOUTA_16_m[0]\, \TFC_DOUTA[0]\, 
        \ELINK_DOUTA_15_m[0]\, \ELINK_DOUTA_14[0]\, 
        un1_SM_BANK_SEL_23, \ELINK_DOUTA_19_m[0]\, 
        \ELINK_DOUTA_10[0]\, un1_SM_BANK_SEL_34, 
        \ELINK_DOUTA_11_m[0]\, \ELINK_DOUTA_8[0]\, 
        un1_SM_BANK_SEL_38, \ELINK_DOUTA_9_m[0]\, 
        \ELINK_DOUTA_6[0]\, \ELINK_DOUTA_7_m[0]\, 
        \ELINK_DOUTA_4[0]\, \ELINK_DOUTA_5_m[0]\, 
        \CHKSUM[0]_net_1\, \N_WR_USB_ADBUS_0_iv_3[0]\, 
        \TFC_STRT_ADDR[0]_net_1\, \N_WR_USB_ADBUS_0_iv_2[0]\, 
        \WR_XFER_TYPE[0]_net_1\, \ELINKS_STOP_ADDR_m[0]\, 
        \OP_MODE_m[0]\, \ELINKS_STRT_ADDR_m[0]\, 
        \N_WR_USB_ADBUS_0_iv_24[6]\, \N_WR_USB_ADBUS_0_iv_13[6]\, 
        \N_WR_USB_ADBUS_0_iv_12[6]\, \N_WR_USB_ADBUS_0_iv_21[6]\, 
        \N_WR_USB_ADBUS_0_iv_23[6]\, \N_WR_USB_ADBUS_0_iv_9[6]\, 
        \N_WR_USB_ADBUS_0_iv_8[6]\, \N_WR_USB_ADBUS_0_iv_19[6]\, 
        \N_WR_USB_ADBUS_0_iv_22[6]\, \N_WR_USB_ADBUS_0_iv_7[6]\, 
        \N_WR_USB_ADBUS_0_iv_6[6]\, \N_WR_USB_ADBUS_0_iv_16[6]\, 
        \ELINK_DOUTA_14_m[6]\, \ELINK_DOUTA_1_m[6]\, 
        \N_WR_USB_ADBUS_0_iv_15[6]\, \ELINK_DOUTA_8_m[6]\, 
        \ELINK_DOUTA_19_m[6]\, \N_WR_USB_ADBUS_0_iv_11[6]\, 
        \N_WR_USB_ADBUS_0_iv_4[6]\, \N_WR_USB_ADBUS_0_iv_3[6]\, 
        \ELINK_DOUTA_3_m[6]\, \ELINK_DOUTA_2[6]\, 
        \ELINK_DOUTA_15_m[6]\, \ELINK_DOUTA_0[6]\, 
        \ELINK_DOUTA_13_m[6]\, \ELINK_DOUTA_11[6]\, 
        un1_SM_BANK_SEL_26, \ELINK_DOUTA_12_m[6]\, 
        \ELINK_DOUTA_9[6]\, un1_SM_BANK_SEL_42, 
        \ELINK_DOUTA_10_m[6]\, \ELINK_DOUTA_17[6]\, 
        \ELINK_DOUTA_18_m[6]\, \ELINK_DOUTA_7[6]\, 
        \ELINK_DOUTA_16_m[6]\, \ELINK_DOUTA_5[6]\, 
        un1_SM_BANK_SEL_35, \ELINK_DOUTA_6_m[6]\, \TFC_DOUTA[6]\, 
        \ELINK_DOUTA_4_m[6]\, \CHKSUM[6]_net_1\, 
        \N_WR_USB_ADBUS_0_iv_2[6]\, \TFC_STRT_ADDR[6]_net_1\, 
        \ELINKS_STOP_ADDR_m[6]\, \OP_MODE_m[6]\, 
        \ELINKS_STRT_ADDR_m[6]\, \N_WR_USB_ADBUS_0_iv_25[1]\, 
        \N_WR_USB_ADBUS_0_iv_14[1]\, \N_WR_USB_ADBUS_0_iv_13[1]\, 
        \N_WR_USB_ADBUS_0_iv_22[1]\, \N_WR_USB_ADBUS_0_iv_24[1]\, 
        \N_WR_USB_ADBUS_0_iv_10[1]\, \N_WR_USB_ADBUS_0_iv_9[1]\, 
        \N_WR_USB_ADBUS_0_iv_20[1]\, \N_WR_USB_ADBUS_0_iv_23[1]\, 
        \N_WR_USB_ADBUS_0_iv_6[1]\, \ELINK_DOUTA_14_m[1]\, 
        \N_WR_USB_ADBUS_0_iv_18[1]\, \ELINK_DOUTA_11_m[1]\, 
        \ELINK_DOUTA_10_m[1]\, \N_WR_USB_ADBUS_0_iv_16[1]\, 
        \ELINK_DOUTA_3_m[1]\, \ELINK_DOUTA_18_m[1]\, 
        \N_WR_USB_ADBUS_0_iv_12[1]\, \TFC_DOUTA_m[1]\, 
        \ELINK_DOUTA_19_m[1]\, \N_WR_USB_ADBUS_0_iv_8[1]\, 
        \ELINK_DOUTA_12[1]\, \ELINK_DOUTA_13_m[1]\, 
        \ELINK_DOUTA_7[1]\, \ELINK_DOUTA_9_m[1]\, 
        \ELINK_DOUTA_6[1]\, \ELINK_DOUTA_8_m[1]\, 
        \ELINK_DOUTA_4[1]\, \ELINK_DOUTA_5_m[1]\, 
        \ELINK_DOUTA_17[1]\, \ELINK_DOUTA_2_m[1]\, 
        \ELINK_DOUTA_16[1]\, \ELINK_DOUTA_1_m[1]\, 
        \ELINK_DOUTA_15[1]\, \ELINK_DOUTA_0_m[1]\, 
        \N_WR_USB_ADBUS_0_iv_3[1]\, \N_WR_USB_ADBUS_0_iv_2[1]\, 
        \N_WR_USB_ADBUS_0_iv_4[1]\, \ELINKS_STRT_ADDR_m[1]\, 
        \CHKSUM_m[1]\, \TFC_STRT_ADDR[1]_net_1\, 
        \ELINKS_STOP_ADDR_m[1]\, \OP_MODE_m[1]\, 
        \TFC_STOP_ADDR_m[1]\, \WR_XFER_TYPE_m[1]\, 
        \N_WR_USB_ADBUS_0_iv_26[2]\, \N_WR_USB_ADBUS_0_iv_18[2]\, 
        \N_WR_USB_ADBUS_0_iv_17[2]\, \N_WR_USB_ADBUS_0_iv_24[2]\, 
        \N_WR_USB_ADBUS_0_iv_10[2]\, \N_WR_USB_ADBUS_0_iv_9[2]\, 
        \N_WR_USB_ADBUS_0_iv_20[2]\, \N_WR_USB_ADBUS_0_iv_22[2]\, 
        \ELINK_DOUTA_17_m[2]\, \ELINK_DOUTA_1_m[2]\, 
        \N_WR_USB_ADBUS_0_iv_16[2]\, \N_WR_USB_ADBUS_0_iv_21[2]\, 
        \ELINK_DOUTA_15_m[2]\, \TFC_DOUTA_m[2]\, 
        \N_WR_USB_ADBUS_0_iv_14[2]\, \ELINK_DOUTA_13_m[2]\, 
        \ELINK_DOUTA_12_m[2]\, \N_WR_USB_ADBUS_0_iv_12[2]\, 
        \ELINK_DOUTA_5_m[2]\, \ELINK_DOUTA_4_m[2]\, 
        \N_WR_USB_ADBUS_0_iv_8[2]\, \N_WR_USB_ADBUS_0_iv_5[2]\, 
        \N_WR_USB_ADBUS_0_iv_4[2]\, \ELINK_DOUTA_3_m[2]\, 
        \ELINK_DOUTA_2[2]\, \ELINK_DOUTA_18_m[2]\, 
        \ELINK_DOUTA_0[2]\, \ELINK_DOUTA_16_m[2]\, 
        \ELINK_DOUTA_14[2]\, \ELINK_DOUTA_19_m[2]\, 
        \ELINK_DOUTA_10[2]\, \ELINK_DOUTA_11_m[2]\, 
        \ELINK_DOUTA_8[2]\, \ELINK_DOUTA_9_m[2]\, 
        \ELINK_DOUTA_6[2]\, \ELINK_DOUTA_7_m[2]\, 
        \CHKSUM[2]_net_1\, \N_WR_USB_ADBUS_0_iv_3[2]\, 
        \TFC_STRT_ADDR[2]_net_1\, \N_WR_USB_ADBUS_0_iv_2[2]\, 
        \ELINKS_STOP_ADDR_m[2]\, \OP_MODE_m[2]\, 
        \ELINKS_STRT_ADDR_m[2]\, \N_WR_USB_ADBUS_0_iv_25[3]\, 
        \N_WR_USB_ADBUS_0_iv_14[3]\, \N_WR_USB_ADBUS_0_iv_13[3]\, 
        \N_WR_USB_ADBUS_0_iv_22[3]\, \N_WR_USB_ADBUS_0_iv_24[3]\, 
        \N_WR_USB_ADBUS_0_iv_10[3]\, \N_WR_USB_ADBUS_0_iv_9[3]\, 
        \N_WR_USB_ADBUS_0_iv_20[3]\, \N_WR_USB_ADBUS_0_iv_23[3]\, 
        \N_WR_USB_ADBUS_0_iv_6[3]\, \ELINK_DOUTA_14_m[3]\, 
        \N_WR_USB_ADBUS_0_iv_18[3]\, \ELINK_DOUTA_11_m[3]\, 
        \ELINK_DOUTA_10_m[3]\, \N_WR_USB_ADBUS_0_iv_16[3]\, 
        \ELINK_DOUTA_3_m[3]\, \ELINK_DOUTA_18_m[3]\, 
        \N_WR_USB_ADBUS_0_iv_12[3]\, \TFC_DOUTA_m[3]\, 
        \ELINK_DOUTA_19_m[3]\, \N_WR_USB_ADBUS_0_iv_8[3]\, 
        \ELINK_DOUTA_12[3]\, \ELINK_DOUTA_13_m[3]\, 
        \ELINK_DOUTA_7[3]\, \ELINK_DOUTA_9_m[3]\, 
        \ELINK_DOUTA_6[3]\, \ELINK_DOUTA_8_m[3]\, 
        \ELINK_DOUTA_4[3]\, \ELINK_DOUTA_5_m[3]\, 
        \ELINK_DOUTA_17[3]\, \ELINK_DOUTA_2_m[3]\, 
        \ELINK_DOUTA_16[3]\, \ELINK_DOUTA_1_m[3]\, 
        \ELINK_DOUTA_15[3]\, \ELINK_DOUTA_0_m[3]\, 
        \N_WR_USB_ADBUS_0_iv_3[3]\, \N_WR_USB_ADBUS_0_iv_2[3]\, 
        \N_WR_USB_ADBUS_0_iv_4[3]\, \ELINKS_STRT_ADDR_m[3]\, 
        \CHKSUM_m[3]\, \TFC_STRT_ADDR[3]_net_1\, 
        \ELINKS_STOP_ADDR_m[3]\, \OP_MODE_m[3]\, 
        \TFC_STOP_ADDR_m[3]\, \WR_XFER_TYPE_m[3]\, 
        \N_WR_USB_ADBUS_0_iv_25[4]\, \N_WR_USB_ADBUS_0_iv_14[4]\, 
        \N_WR_USB_ADBUS_0_iv_13[4]\, \N_WR_USB_ADBUS_0_iv_22[4]\, 
        \N_WR_USB_ADBUS_0_iv_24[4]\, \N_WR_USB_ADBUS_0_iv_10[4]\, 
        \N_WR_USB_ADBUS_0_iv_9[4]\, \N_WR_USB_ADBUS_0_iv_20[4]\, 
        \N_WR_USB_ADBUS_0_iv_23[4]\, \N_WR_USB_ADBUS_0_iv_8[4]\, 
        \N_WR_USB_ADBUS_0_iv_7[4]\, \N_WR_USB_ADBUS_0_iv_17[4]\, 
        \ELINK_DOUTA_17_m[4]\, \ELINK_DOUTA_1_m[4]\, 
        \N_WR_USB_ADBUS_0_iv_16[4]\, \ELINK_DOUTA_13_m[4]\, 
        \ELINK_DOUTA_12_m[4]\, \N_WR_USB_ADBUS_0_iv_12[4]\, 
        \N_WR_USB_ADBUS_0_iv_5[4]\, \N_WR_USB_ADBUS_0_iv_4[4]\, 
        \ELINK_DOUTA_3_m[4]\, \ELINK_DOUTA_2[4]\, 
        \ELINK_DOUTA_18_m[4]\, \ELINK_DOUTA_0[4]\, 
        \ELINK_DOUTA_16_m[4]\, \TFC_DOUTA[4]\, 
        \ELINK_DOUTA_15_m[4]\, \ELINK_DOUTA_14[4]\, 
        \ELINK_DOUTA_19_m[4]\, \ELINK_DOUTA_10[4]\, 
        \ELINK_DOUTA_11_m[4]\, \ELINK_DOUTA_8[4]\, 
        \ELINK_DOUTA_9_m[4]\, \ELINK_DOUTA_6[4]\, 
        \ELINK_DOUTA_7_m[4]\, \ELINK_DOUTA_4[4]\, 
        \ELINK_DOUTA_5_m[4]\, \CHKSUM[4]_net_1\, 
        \N_WR_USB_ADBUS_0_iv_3[4]\, \TFC_STRT_ADDR[4]_net_1\, 
        \N_WR_USB_ADBUS_0_iv_2[4]\, \ELINKS_STOP_ADDR_m[4]\, 
        \OP_MODE_m[4]\, \ELINKS_STRT_ADDR_m[4]\, 
        \REG_STATE_ns_i_4[1]\, \REG_STATE_ns_i_a4_0[1]\, 
        N_1282_tz, N_2587, \REG_STATE_ns_i_3[1]\, N_1278_tz, 
        \REG_STATE_ns_i_a4_8_0[1]\, \REG_STATE_ns_i_2[1]\, 
        N_1275_tz, \REG_STATE_ns_i_1[1]\, N_2539, N_2546, N_2537, 
        \REG_STATE_ns_i_i_0[2]\, \REG_STATE_ns_i_i_a5_1_3[0]\, 
        N_504, N_384, \REG_STATE_ns_i_i_a5_1_2[0]\, N_282, 
        N_USB_OE_BI_iv_0_i_a2_0_1, N_385_1, 
        \REG_STATE_ns_i_1_0[3]\, \REG_STATE_ns_i_a4_0_0[3]\, 
        N_1259_tz, N_2592, \REG_STATE_ns_i_0[3]\, 
        \REG_STATE_ns_i_1_tz[3]\, N_2561, N_2498, 
        \REG_STATE_ns_i_i_a2_0[0]_net_1\, N_1351_8, N_1398_i_0_0, 
        N_2616, N_2617, un1_N_ELK_N_ACTIVE_0_sqmuxa_15_0_a2_0_0, 
        \REG_STATE_ns_i_a2_1[4]\, N_285, \REG_STATE_ns_i_a2_0[4]\, 
        REG_STATE_tr67_5, N_1404_8, N_1387_i, N_287, N_413, N_412, 
        N_1359_1, \REG_STATE_ns_i_i_a2_5_0[0]\, N_452, 
        \REG_STATE_ns_i_a2_0[1]\, REG_STATE_tr74_1, 
        \N_ELINK_RWA_i_a2_0_a5_0[16]\, \SM_BANK_SEL[6]_net_1\, 
        \SM_BANK_SEL[5]_net_1\, \SM_BANK_SEL[4]_net_1\, 
        \N_ELINK_RWA_0_iv_0_o2_i_a5_0[15]\, 
        \SM_BANK_SEL[3]_net_1\, 
        \N_ELINK_RWA_0_iv_0_o2_i_a5_0[13]\, N_462, 
        un1_N_ELK_N_ACTIVE_2_sqmuxa_0_a2_0_0, N_1903, 
        \REG_STATE_ns_i_a2_0[3]\, N_480, un1_REG_STATE_40_i_o2_0, 
        N_1751, un1_REG_STATE_40_i_a2_0_0, N_1877, 
        un1_REG_STATE_26_0_1, N_2526_1, N_1745_i, 
        un1_REG_STATE_26_0_0, N_1749, 
        \REG_STATE_ns_i_i_o2_10_5[2]\, 
        \REG_STATE_ns_i_i_o2_10_3[2]\, 
        \REG_STATE_ns_i_i_o2_10_2[2]\, N_349, N_470, N_256, N_415, 
        N_418, \REG_STATE_ns_i_i_o2_10_0[2]\, N_417, N_433_1, 
        N_260, N_428, \N_ELINK_BLKA_0_iv_0_o2_i_a5_2[9]\, N_461, 
        \N_ELINK_BLKA_0_iv_0_o2_i_a5_0[9]\, N_477, 
        \SM_BANK_SEL[9]_net_1\, \SM_BANK_SEL[11]_net_1\, 
        \REG_STATE_ns_i_a2_0_0[5]\, \REG_STATE_ns_i_a2_0_0_2[5]\, 
        \REG_STATE_ns_i_a2_4_2[5]\, un1_REG_STATE_28_0_0, 
        N_1761_i, REG_ADDR_n2_i_0, \REG_ADDR[0]_net_1\, 
        \REG_ADDR[1]_net_1\, \REG_ADDR[2]_net_1\, N_USB_RD_BI_i_5, 
        N_1869, N_1868, N_USB_RD_BI_i_4, N_USB_RD_BI_i_1, N_1865, 
        N_1744_i, N_1864, \N_ELINK_BLKA_0_iv_0_o2_i_a5_1[11]\, 
        N_469, \SM_BANK_SEL[7]_net_1\, N_1351_i_i_a5_2, 
        N_1351_i_i_a5_0, N_465, N_1387_i_0_2, N_1387_i_0_1, N_459, 
        N_356, N_1368_i_i_a5_0, \RD_XFER_TYPE[1]_net_1\, 
        \RD_XFER_TYPE[0]_net_1\, N_1370_i_i_a5_0, N_1398_i_0_a2_3, 
        N_474, N_252, \REG_STATE_ns_i_tz_1[5]\, N_2577, 
        \REG_STATE_ns_i_tz_0[5]\, N_2515, un1_REG_STATE_35_i_a2_0, 
        \RD_USB_ADBUS[6]_net_1\, \REG_STATE_ns_i_i_a2_1_0[0]\, 
        N_TFC_STRT_ADDR_T_0_sqmuxa_0_a2_0, \USB_RXF_B\, 
        \N_ELINK_RWA_3[0]\, N_143, N_616_11, \N_ELINK_RWA_1[0]\, 
        \SM_BANK_SEL[17]_net_1\, \SM_BANK_SEL[18]_net_1\, N_616_2, 
        \N_ELINK_RWA_3[1]\, \N_ELINK_RWA_1[1]\, 
        \SM_BANK_SEL[19]_net_1\, \N_ELINK_RWA_1[2]\, N_618_1, 
        \N_ELINK_RWA_3[5]\, N_620_10, \N_ELINK_RWA_1[5]\, 
        \SM_BANK_SEL[15]_net_1\, \SM_BANK_SEL[13]_net_1\, N_616_4, 
        \N_ELINK_RWA_3[3]\, \N_ELINK_RWA_1[3]\, 
        \N_ELINK_RWA_1[6]\, N_622_3, \N_ELINK_RWA_3[7]\, 
        \N_ELINK_RWA_1[7]\, REG_STATE_tr67_3, N_1404_7, N_1404_6, 
        REG_STATE_tr67_0, REG_STATE_tr67_1, 
        \WR_XFER_TYPE[1]_net_1\, REG_STATE_tr72_6_5, 
        REG_STATE_tr72_6_3, REG_STATE_tr72_6_0, 
        REG_STATE_tr72_6_1, \REG_STATE_ns_i_i_a2_9_0[0]\, 
        \REG_STATE[5]_net_1\, REG_STATE_tr73_9, REG_STATE_tr73_7, 
        REG_STATE_tr73_6, N_1421_3, REG_STATE_tr73_2, 
        REG_STATE_tr73_1, REG_STATE_tr73_4, \REG_ADDR[6]_net_1\, 
        \REG_ADDR[7]_net_1\, \REG_ADDR[8]_net_1\, 
        \REG_ADDR[3]_net_1\, \REG_ADDR[4]_net_1\, 
        \REG_ADDR[5]_net_1\, REG_STATE_ns_i_245_tz_0, 
        \REG_STATE_ns_i_a4_1_1_0[1]\, N_1879_1, 
        \REG_STATE_ns_i_a4_10_0[1]\, \REG_STATE_ns_i_a2_0_0_0[5]\, 
        \REG_STATE_ns_i_a2_4_0[5]\, 
        \REG_STATE_ns_i_a2_4_tz_tz_tz_tz[5]\, \N_ELINK_RWA_0[8]\, 
        N_624_15, \N_ELINK_RWA_1[4]\, \N_ELINK_RWA_3[14]\, N_365, 
        \N_ELINK_RWA_1[14]\, \N_ELINK_RWA_2[10]\, 
        \N_ELINK_RWA_0[10]\, \SM_BANK_SEL[10]_net_1\, 
        REG_STATE_tr74_tz_tz_tz_5, REG_STATE_tr74_tz_tz_tz_6, 
        REG_STATE_tr74_0, REG_STATE_s22_i_0, N_1499_2_i_0, 
        REG_STATE_tr49_6, REG_STATE_tr49_3, REG_STATE_tr49_2, 
        REG_STATE_tr49_4, N_491, \N_ELINK_RWA_1[12]\, 
        \N_ELINK_RWA_0_iv_0_o2_0[18]\, N_463, N_394, 
        \REG_STATE_ns_i_i_a5_1_1_0[2]\, REG_STATE_s20_i_0, 
        N_1367_i_i_a2_3, N_1367_i_i_a2_2, N_1351_3, 
        N_1367_i_i_a2_0, N_1359_6, \N_ELINK_RWA_16_0[0]\, 
        un1_REG_STATE_40_i_a2_2_0, un1_REG_STATE_39_i_a2_0, 
        N_1862_1, \REG_STATE_ns_i_1_tz_1[3]\, N_339, 
        \REG_STATE_ns_i_1_tz_0[3]\, N_2600, \N_ELINK_RWA_15_1[8]\, 
        \SM_BANK_SEL[12]_net_1\, N_1778, N_1739, 
        \REG_STATE_ns_i_i_a5_0_1_0[2]\, N_USB_OE_BI_iv_0_i_a2_0_5, 
        N_USB_OE_BI_iv_0_i_a2_0_4, N_1352_5, 
        \REG_STATE_ns_i_a4_3_0[4]\, N_1398_i_0_a2_1, 
        N_1398_i_0_a2_0, N_USB_RD_BI_i_a2_4_3, 
        N_USB_RD_BI_i_a2_4_1, \N_TFC_ADDRA_0_a2_1_1[7]\, N_292, 
        \REG_STATE_ns_i_a4_7_0[4]\, N_2613, 
        \N_TFC_ADDRA_0_a2_6_0[7]\, un1_REG_STATE_40_i_a2_3_0, 
        \REG_STATE_ns_i_a4_3_1_0[1]\, N_2571_1, 
        un1_REG_STATE_40_i_a2_0, \N_ELINK_BLKA_10_0[10]\, 
        \SM_BANK_SEL[16]_net_1\, REG_STATE_tr74_tz_tz_tz_4, 
        REG_STATE_tr74_tz_tz_tz_2, \REG_STATE_ns_i_a2_2_0[4]\, 
        \SI_CNT[3]_net_1\, \SI_CNT[2]_net_1\, N_1367_i_i_o2_0_2, 
        \RD_XFER_TYPE[4]_net_1\, \RD_XFER_TYPE[5]_net_1\, 
        N_1367_i_i_o2_0_1, \RD_XFER_TYPE[7]_net_1\, 
        \RD_XFER_TYPE[6]_net_1\, N_1367_i_i_o2_0_0, 
        \RD_XFER_TYPE[3]_net_1\, \RD_XFER_TYPE[2]_net_1\, 
        \N_WR_USB_ADBUS[0]\, \N_WR_USB_ADBUS[1]\, 
        \N_WR_USB_ADBUS[2]\, \N_WR_USB_ADBUS[3]\, 
        \N_WR_USB_ADBUS[4]\, \N_WR_USB_ADBUS[5]\, 
        \N_WR_USB_ADBUS[6]\, \N_WR_USB_ADBUS[7]\, N_616_16, N_618, 
        N_1419, N_1879, N_2581, N_359, 
        \WR_XFER_TYPE_RNO[0]_net_1\, N_1816, N_1818, N_1817, 
        N_513, \RD_USB_ADBUS_RNIP4GES[4]_net_1\, N_393, N_464, 
        N_392, \REG_STATE_d[30]\, N_1736, \RD_USB_ADBUS[0]_net_1\, 
        \RD_USB_ADBUS[1]_net_1\, N_TFC_STRT_ADDR_T_0_sqmuxa, 
        N_2629, N_675, N_257, N_1756, N_1886, N_1887, N_1911, 
        N_1713, un1_REG_STATE_26, N_1784, N_454, 
        N_OP_MODE_T_0_sqmuxa, N_1765, N_396, REG_ADDRe, N_1673, 
        N_1867, N_1866, N_511_1, N_388, N_274, N_255, N_273, 
        N_277, N_1821, N_1819, \WR_XFER_TYPE_RNO[1]_net_1\, 
        N_1820, N_44, N_2607, N_678, N_1862, N_488, N_489, N_310, 
        N_510, N_457, N_456, N_268, \REG_STATE_ns_i_6[4]\, N_438, 
        N_2462, N_441, N_440, N_439, N_436, N_414_1, 
        un1_REG_STATE_28, N_1779, \SM_BANK_SEL[14]_net_1\, N_622, 
        \REG_STATE_ns_i_i_a5_1[2]\, \REG_STATE_ns_i_a4_6_1[4]\, 
        N_2467, \REG_STATE_ns_i_a4_3_0[3]\, 
        \REG_STATE_ns_i_8_tz[4]\, N_2454_tz, N_2520, 
        \REG_STATE_ns_i_a4_8_0_a5_0[4]\, N_1294_tz, N_311, N_2602, 
        \REG_STATE_ns_i_a4_7_0[1]\, N_2628, N_2477_i, N_2622, 
        \REG_STATE_ns_i_a4_1_0[3]\, N_63, \SM_BANK_SEL[1]_net_1\, 
        X_BLKA_i, N_63_tz, \ELINK_BLKA[18]_net_1\, N_65, N_65_tz, 
        N_503, \ELINK_BLKA[15]_net_1\, N_67, N_67_tz, 
        \ELINK_BLKA[13]_net_1\, REG_ADDR_n8, REG_ADDR_75_0, 
        REG_ADDR_n7, REG_ADDR_c6, REG_ADDR_n6, REG_ADDR_c5, 
        REG_ADDR_n4, REG_ADDR_c3, REG_ADDR_n3, REG_ADDR_n5, 
        REG_ADDR_c4, SI_CNT_n3, N_1630, \N_ELINK_BLKA_0_iv[17]\, 
        N_131, \ELINK_BLKA[17]_net_1\, X_BLKA_i_m_16, 
        \N_ELINK_BLKA_0_iv[19]\, N_130, \ELINK_BLKA[19]_net_1\, 
        X_BLKA_i_m_18, N_162, \SM_BANK_SEL[8]_net_1\, N_164, 
        N_165, \ELINK_BLKA[5]_net_1\, N_167, 
        \ELINK_BLKA[1]_net_1\, N_170, \SM_BANK_SEL[0]_net_1\, 
        un1_USB_RXF_B_m, N_174, \SM_BANK_SEL[2]_net_1\, N_175, 
        \ELINK_RWA[15]_net_1\, N_177, \ELINK_RWA[13]_net_1\, 
        N_180, N_182, N_183, \ELINK_RWA[5]_net_1\, N_185, 
        \ELINK_RWA[1]_net_1\, \N_ELINK_BLKA_0_iv[11]\, 
        \ELINK_BLKA[11]_net_1\, \N_ELINK_BLKA_0_iv[9]\, 
        \ELINK_BLKA[9]_net_1\, \N_ELINK_BLKA_0_iv[5]\, 
        \N_ELINK_BLKA_0_iv[1]\, \N_ELINK_RWA_0_iv[19]\, 
        \ELINK_RWA[19]_net_1\, \N_ELINK_RWA_0_iv[17]\, 
        \ELINK_RWA[17]_net_1\, \N_ELINK_RWA_0_iv[15]\, 
        \N_ELINK_RWA_0_iv[13]\, \N_ELINK_RWA_0_iv[11]\, 
        \ELINK_RWA[11]_net_1\, \N_ELINK_RWA_0_iv[9]\, 
        \ELINK_RWA[9]_net_1\, \N_ELINK_RWA_0_iv[5]\, 
        \N_ELINK_RWA_0_iv[1]\, N_1905, N_1703, N_1679, N_1871, 
        N_1669, \RD_XFER_TYPE_RNO[7]_net_1\, N_1808, 
        \RD_XFER_TYPE_RNO[6]_net_1\, N_1806, 
        \RD_XFER_TYPE_RNO[5]_net_1\, N_1804, 
        \RD_XFER_TYPE_RNO[2]_net_1\, N_1798, 
        \RD_XFER_TYPE_RNO[1]_net_1\, N_1796, 
        \RD_XFER_TYPE_RNO[0]_net_1\, N_1794, N_1891, N_1849, 
        N_1848, N_1843, N_1841, N_1840, N_1838, N_1835, 
        \N_ELINK_BLKA_0_iv[16]\, \ELINK_BLKA_i_m[16]\, 
        \ELINK_BLKA[16]_net_1\, \N_ELINK_BLKA_0_iv[14]\, 
        \ELINK_BLKA_i_m[14]\, \ELINK_BLKA[14]_net_1\, 
        \N_ELINK_BLKA_0_iv[12]\, \ELINK_BLKA_i_m[12]\, 
        \ELINK_BLKA[12]_net_1\, \N_ELINK_BLKA_0_iv[10]\, 
        \ELINK_BLKA_i_m[10]\, \ELINK_BLKA[10]_net_1\, 
        \N_ELINK_BLKA_0_iv[8]\, \ELINK_BLKA_i_m[8]\, 
        \ELINK_BLKA[8]_net_1\, \N_ELINK_BLKA_0_iv[6]\, 
        \ELINK_BLKA[6]_net_1\, X_BLKA_i_m_5, 
        \N_ELINK_BLKA_0_iv[3]\, \ELINK_BLKA_i_m[3]\, 
        \ELINK_BLKA[3]_net_1\, \N_ELINK_BLKA_0_iv[2]\, 
        \ELINK_BLKA[2]_net_1\, X_BLKA_i_m_1, 
        \N_ELINK_BLKA_0_iv[0]\, \ELINK_BLKA_i_m[0]\, 
        \ELINK_BLKA[0]_net_1\, \N_ELINK_RWA_0_iv[16]\, 
        \ELINK_RWA_i_m[16]\, \ELINK_RWA[16]_net_1\, 
        \N_ELINK_RWA_0_iv[14]\, \ELINK_RWA_i_m[14]\, 
        \ELINK_RWA[14]_net_1\, \N_ELINK_RWA_0_iv[12]\, 
        \ELINK_RWA_i_m[12]\, \ELINK_RWA[12]_net_1\, 
        \N_ELINK_RWA_0_iv[10]\, \ELINK_RWA_i_m[10]\, 
        \ELINK_RWA[10]_net_1\, \N_ELINK_RWA_0_iv[8]\, 
        \ELINK_RWA_i_m[8]\, \ELINK_RWA[8]_net_1\, 
        \N_ELINK_RWA_0_iv[6]\, \ELINK_RWA_i_m[6]\, 
        \ELINK_RWA[6]_net_1\, \N_ELINK_RWA_0_iv[3]\, 
        \ELINK_RWA_i_m[3]\, \ELINK_RWA[3]_net_1\, 
        \N_ELINK_RWA_0_iv[2]\, \ELINK_RWA_i_m[2]\, 
        \ELINK_RWA[2]_net_1\, \N_ELINK_RWA_0_iv[0]\, 
        \ELINK_RWA_i_m[0]\, \ELINK_RWA[0]_net_1\, 
        \ELINK_DOUTA_19[7]\, un1_SM_BANK_SEL_41, 
        \ELINK_DOUTA_18[7]\, un1_SM_BANK_SEL_25, 
        \ELINK_DOUTA_14[7]\, \ELINK_DOUTA_13[7]\, 
        un1_SM_BANK_SEL_29, \ELINK_DOUTA_11[7]\, 
        \ELINK_DOUTA_10[7]\, \ELINK_DOUTA_9[7]\, 
        \ELINK_DOUTA_8[7]\, \ELINK_DOUTA_5[7]\, 
        \ELINK_DOUTA_3[7]\, un1_SM_BANK_SEL_43, 
        \ELINK_DOUTA_2[7]\, \ELINK_DOUTA_1[7]\, 
        un1_SM_BANK_SEL_36, \ELINK_DOUTA_0[7]\, \TFC_DOUTA[7]\, 
        N_1730_i, \ELINKS_STOP_ADDR[7]_net_1\, \OP_MODE[7]_net_1\, 
        \ELINK_DOUTA_19[6]\, \ELINK_DOUTA_18[6]\, 
        \ELINK_DOUTA_16[6]\, \ELINK_DOUTA_15[6]\, 
        \ELINK_DOUTA_14[6]\, \ELINK_DOUTA_13[6]\, 
        \ELINK_DOUTA_12[6]\, \ELINK_DOUTA_10[6]\, 
        \ELINK_DOUTA_8[6]\, \ELINK_DOUTA_6[6]\, 
        \ELINK_DOUTA_4[6]\, \ELINK_DOUTA_3[6]\, 
        \ELINK_DOUTA_1[6]\, \ELINKS_STOP_ADDR[6]_net_1\, 
        \ELINKS_STRT_ADDR[6]_net_1\, \OP_MODE[6]_net_1\, 
        \ELINK_DOUTA_19[5]\, \ELINK_DOUTA_18[5]\, 
        \ELINK_DOUTA_14[5]\, \ELINK_DOUTA_13[5]\, 
        \ELINK_DOUTA_11[5]\, \ELINK_DOUTA_10[5]\, 
        \ELINK_DOUTA_9[5]\, \ELINK_DOUTA_8[5]\, 
        \ELINK_DOUTA_6[5]\, \ELINK_DOUTA_5[5]\, 
        \ELINK_DOUTA_3[5]\, \ELINK_DOUTA_2[5]\, 
        \ELINK_DOUTA_1[5]\, \ELINK_DOUTA_0[5]\, \TFC_DOUTA[5]\, 
        \CHKSUM[5]_net_1\, \ELINKS_STOP_ADDR[5]_net_1\, 
        \ELINKS_STRT_ADDR[5]_net_1\, \TFC_STOP_ADDR[5]_net_1\, 
        \OP_MODE[5]_net_1\, \ELINK_DOUTA_19[4]\, 
        \ELINK_DOUTA_18[4]\, \ELINK_DOUTA_17[4]\, 
        \ELINK_DOUTA_16[4]\, \ELINK_DOUTA_15[4]\, 
        \ELINK_DOUTA_13[4]\, \ELINK_DOUTA_12[4]\, 
        \ELINK_DOUTA_11[4]\, \ELINK_DOUTA_9[4]\, 
        \ELINK_DOUTA_7[4]\, \ELINK_DOUTA_5[4]\, 
        \ELINK_DOUTA_3[4]\, \ELINK_DOUTA_1[4]\, 
        \ELINKS_STOP_ADDR[4]_net_1\, \ELINKS_STRT_ADDR[4]_net_1\, 
        \OP_MODE[4]_net_1\, \ELINK_DOUTA_19[3]\, 
        \ELINK_DOUTA_18[3]\, \ELINK_DOUTA_14[3]\, 
        \ELINK_DOUTA_13[3]\, \ELINK_DOUTA_11[3]\, 
        \ELINK_DOUTA_10[3]\, \ELINK_DOUTA_9[3]\, 
        \ELINK_DOUTA_8[3]\, \ELINK_DOUTA_5[3]\, 
        \ELINK_DOUTA_3[3]\, \ELINK_DOUTA_2[3]\, 
        \ELINK_DOUTA_1[3]\, \ELINK_DOUTA_0[3]\, \TFC_DOUTA[3]\, 
        \CHKSUM[3]_net_1\, \ELINKS_STOP_ADDR[3]_net_1\, 
        \ELINKS_STRT_ADDR[3]_net_1\, \TFC_STOP_ADDR[3]_net_1\, 
        \OP_MODE[3]_net_1\, \ELINK_DOUTA_19[2]\, 
        \ELINK_DOUTA_18[2]\, \ELINK_DOUTA_17[2]\, 
        \ELINK_DOUTA_16[2]\, \ELINK_DOUTA_15[2]\, 
        \ELINK_DOUTA_13[2]\, \ELINK_DOUTA_12[2]\, 
        \ELINK_DOUTA_11[2]\, \ELINK_DOUTA_9[2]\, 
        \ELINK_DOUTA_7[2]\, \ELINK_DOUTA_5[2]\, 
        \ELINK_DOUTA_4[2]\, \ELINK_DOUTA_3[2]\, 
        \ELINK_DOUTA_1[2]\, \TFC_DOUTA[2]\, 
        \ELINKS_STOP_ADDR[2]_net_1\, \ELINKS_STRT_ADDR[2]_net_1\, 
        \OP_MODE[2]_net_1\, \ELINK_DOUTA_19[1]\, 
        \ELINK_DOUTA_18[1]\, \ELINK_DOUTA_14[1]\, 
        \ELINK_DOUTA_13[1]\, \ELINK_DOUTA_11[1]\, 
        \ELINK_DOUTA_10[1]\, \ELINK_DOUTA_9[1]\, 
        \ELINK_DOUTA_8[1]\, \ELINK_DOUTA_5[1]\, 
        \ELINK_DOUTA_3[1]\, \ELINK_DOUTA_2[1]\, 
        \ELINK_DOUTA_1[1]\, \ELINK_DOUTA_0[1]\, \TFC_DOUTA[1]\, 
        \CHKSUM[1]_net_1\, \ELINKS_STOP_ADDR[1]_net_1\, 
        \ELINKS_STRT_ADDR[1]_net_1\, \TFC_STOP_ADDR[1]_net_1\, 
        \OP_MODE[1]_net_1\, \ELINK_DOUTA_19[0]\, 
        \ELINK_DOUTA_18[0]\, \ELINK_DOUTA_17[0]\, 
        \ELINK_DOUTA_16[0]\, \ELINK_DOUTA_15[0]\, 
        \ELINK_DOUTA_13[0]\, \ELINK_DOUTA_12[0]\, 
        \ELINK_DOUTA_11[0]\, \ELINK_DOUTA_9[0]\, 
        \ELINK_DOUTA_7[0]\, \ELINK_DOUTA_5[0]\, 
        \ELINK_DOUTA_3[0]\, \ELINK_DOUTA_1[0]\, 
        \ELINKS_STOP_ADDR[0]_net_1\, \ELINKS_STRT_ADDR[0]_net_1\, 
        \OP_MODE[0]_net_1\, N_TFC_BLKA, \SM_BANK_SEL[21]_net_1\, 
        un1_SM_BANK_SEL_21, un1_SM_BANK_SEL_15, 
        un1_SM_BANK_SEL_12, un1_SM_BANK_SEL_11, 
        un1_SM_BANK_SEL_10, un1_SM_BANK_SEL_9, un1_SM_BANK_SEL_7, 
        un1_SM_BANK_SEL_5, \N_TFC_DINA[0]\, N_206, 
        \N_TFC_DINA[3]\, \N_TFC_ADDRA[7]\, \N_TFC_ADDRA[6]\, 
        \N_TFC_ADDRA[5]\, \N_TFC_ADDRA[3]\, \N_TFC_ADDRA[2]\, 
        N_486, N_198, N_197, \N_TFC_DINA[1]\, \N_TFC_DINA[2]\, 
        \N_TFC_DINA[5]\, \N_TFC_DINA[6]\, \N_TFC_DINA[7]\, N_142, 
        N_346, N_ELINKS_STOP_ADDR_T_0_sqmuxa, N_1907, N_1860, 
        N_1917, N_1833, N_1834, N_1873, N_1893, N_1772, N_1737, 
        \ELK_N_ACTIVE_RNO\, N_1698, N_1728, N_254, N_446, N_427, 
        \N_TFC_ADDRA[0]\, REG_ADDR_n1, N_2624, N_199, N_200, 
        \N_TFC_ADDRA[1]\, \N_TFC_ADDRA[4]\, un1_SM_BANK_SEL_1, 
        un1_SM_BANK_SEL_2, un1_SM_BANK_SEL_16, un1_SM_BANK_SEL_20, 
        N_424, N_432, N_259, N_253, N_2537_1, N_1729, SI_CNTe, 
        un1_REG_STATE_18, \ELINK_RWA_i_m[7]\, 
        \ELINK_RWA[7]_net_1\, \N_ELINK_RWA_0_iv[7]\, 
        \ELINK_BLKA_i_m[7]\, \ELINK_BLKA[7]_net_1\, 
        \N_ELINK_BLKA_0_iv[7]\, N_1675, \N_ELINK_RWA_0_iv[18]\, 
        N_171, \ELINK_RWA[18]_net_1\, N_449, N_450, N_262_i, 
        N_1800, N_1802, \RD_XFER_TYPE_RNO[3]_net_1\, 
        \RD_XFER_TYPE_RNO[4]_net_1\, \WR_XFER_TYPE_RNO[7]_net_1\, 
        SI_CNT_n1, \SI_CNT[1]_net_1\, \SI_CNT[0]_net_1\, N_2625, 
        N_350, \N_TFC_DINA[4]\, un1_SM_BANK_SEL_4, 
        un1_SM_BANK_SEL_6, un1_SM_BANK_SEL_8, un1_SM_BANK_SEL_19, 
        N_1844, N_1850, N_1851, N_471, N_1352_2, N_437, N_234, 
        un1_REG_STATE_22, N_226, N_228, 
        N_TFC_STOP_ADDR_T_0_sqmuxa, N_1587, N_1593, N_236, N_232, 
        N_230, \ELINK_RWA_i_m[4]\, \ELINK_RWA[4]_net_1\, 
        \N_ELINK_RWA_0_iv[4]\, \ELINK_BLKA_i_m[4]\, 
        \ELINK_BLKA[4]_net_1\, \N_ELINK_BLKA_0_iv[4]\, 
        N_ELINKS_STRT_ADDR_T_0_sqmuxa, \TFC_BLKA\, \TFC_RWA\, 
        \TFC_STRT_ADDR_T[0]_net_1\, \TFC_STRT_ADDR_T[1]_net_1\, 
        \TFC_STRT_ADDR_T[2]_net_1\, \TFC_STRT_ADDR_T[3]_net_1\, 
        \TFC_STRT_ADDR_T[4]_net_1\, \TFC_STRT_ADDR_T[5]_net_1\, 
        \TFC_STRT_ADDR_T[6]_net_1\, \TFC_STRT_ADDR_T[7]_net_1\, 
        \TFC_STOP_ADDR_T[0]_net_1\, \TFC_STOP_ADDR_T[1]_net_1\, 
        \TFC_STOP_ADDR_T[2]_net_1\, \TFC_STOP_ADDR_T[3]_net_1\, 
        \TFC_STOP_ADDR_T[4]_net_1\, \TFC_STOP_ADDR_T[5]_net_1\, 
        \TFC_STOP_ADDR_T[6]_net_1\, \TFC_STOP_ADDR_T[7]_net_1\, 
        \OP_MODE_T[0]_net_1\, \OP_MODE_T[1]_net_1\, 
        \OP_MODE_T[2]_net_1\, \OP_MODE_T[3]_net_1\, 
        \OP_MODE_T[4]_net_1\, \OP_MODE_T[5]_net_1\, 
        \OP_MODE_T[6]_net_1\, \OP_MODE_T[7]_net_1\, 
        \ELINKS_STRT_ADDR_T[0]_net_1\, 
        \ELINKS_STRT_ADDR_T[1]_net_1\, 
        \ELINKS_STRT_ADDR_T[2]_net_1\, 
        \ELINKS_STRT_ADDR_T[3]_net_1\, 
        \ELINKS_STRT_ADDR_T[4]_net_1\, 
        \ELINKS_STRT_ADDR_T[5]_net_1\, 
        \ELINKS_STRT_ADDR_T[6]_net_1\, 
        \ELINKS_STRT_ADDR_T[7]_net_1\, 
        \ELINKS_STOP_ADDR_T[0]_net_1\, 
        \ELINKS_STOP_ADDR_T[1]_net_1\, 
        \ELINKS_STOP_ADDR_T[2]_net_1\, 
        \ELINKS_STOP_ADDR_T[3]_net_1\, 
        \ELINKS_STOP_ADDR_T[4]_net_1\, 
        \ELINKS_STOP_ADDR_T[5]_net_1\, 
        \ELINKS_STOP_ADDR_T[6]_net_1\, 
        \ELINKS_STOP_ADDR_T[7]_net_1\, \ELINK_DINA_8[0]_net_1\, 
        \ELINK_DINA_8[1]_net_1\, \ELINK_DINA_8[2]_net_1\, 
        \ELINK_DINA_8[3]_net_1\, \ELINK_DINA_8[4]_net_1\, 
        \ELINK_DINA_8[5]_net_1\, \ELINK_DINA_8[6]_net_1\, 
        \ELINK_DINA_8[7]_net_1\, \ELINK_DINA_7[0]_net_1\, 
        \ELINK_DINA_7[1]_net_1\, \ELINK_DINA_7[2]_net_1\, 
        \ELINK_DINA_7[3]_net_1\, \ELINK_DINA_7[4]_net_1\, 
        \ELINK_DINA_7[5]_net_1\, \ELINK_DINA_7[6]_net_1\, 
        \ELINK_DINA_7[7]_net_1\, \ELINK_DINA_6[0]_net_1\, 
        \ELINK_DINA_6[1]_net_1\, \ELINK_DINA_6[2]_net_1\, 
        \ELINK_DINA_6[3]_net_1\, \ELINK_DINA_6[4]_net_1\, 
        \ELINK_DINA_6[5]_net_1\, \ELINK_DINA_6[6]_net_1\, 
        \ELINK_DINA_6[7]_net_1\, \ELINK_DINA_5[0]_net_1\, 
        \ELINK_DINA_5[1]_net_1\, \ELINK_DINA_5[2]_net_1\, 
        \ELINK_DINA_5[3]_net_1\, \ELINK_DINA_5[4]_net_1\, 
        \ELINK_DINA_5[5]_net_1\, \ELINK_DINA_5[6]_net_1\, 
        \ELINK_DINA_5[7]_net_1\, \ELINK_DINA_4[0]_net_1\, 
        \ELINK_DINA_4[1]_net_1\, \ELINK_DINA_4[2]_net_1\, 
        \ELINK_DINA_4[3]_net_1\, \ELINK_DINA_4[4]_net_1\, 
        \ELINK_DINA_4[5]_net_1\, \ELINK_DINA_4[6]_net_1\, 
        \ELINK_DINA_4[7]_net_1\, \ELINK_DINA_3[0]_net_1\, 
        \ELINK_DINA_3[1]_net_1\, \ELINK_DINA_3[2]_net_1\, 
        \ELINK_DINA_3[3]_net_1\, \ELINK_DINA_3[4]_net_1\, 
        \ELINK_DINA_3[5]_net_1\, \ELINK_DINA_3[6]_net_1\, 
        \ELINK_DINA_3[7]_net_1\, \ELINK_DINA_2[0]_net_1\, 
        \ELINK_DINA_2[1]_net_1\, \ELINK_DINA_2[2]_net_1\, 
        \ELINK_DINA_2[3]_net_1\, \ELINK_DINA_2[4]_net_1\, 
        \ELINK_DINA_2[5]_net_1\, \ELINK_DINA_2[6]_net_1\, 
        \ELINK_DINA_2[7]_net_1\, \ELINK_DINA_1[0]_net_1\, 
        \ELINK_DINA_1[1]_net_1\, \ELINK_DINA_1[2]_net_1\, 
        \ELINK_DINA_1[3]_net_1\, \ELINK_DINA_1[4]_net_1\, 
        \ELINK_DINA_1[5]_net_1\, \ELINK_DINA_1[6]_net_1\, 
        \ELINK_DINA_1[7]_net_1\, \ELINK_DINA_0[0]_net_1\, 
        \ELINK_DINA_0[1]_net_1\, \ELINK_DINA_0[2]_net_1\, 
        \ELINK_DINA_0[3]_net_1\, \ELINK_DINA_0[4]_net_1\, 
        \ELINK_DINA_0[5]_net_1\, \ELINK_DINA_0[6]_net_1\, 
        \ELINK_DINA_0[7]_net_1\, \WR_USB_ADBUS[0]_net_1\, 
        \WR_USB_ADBUS[1]_net_1\, \WR_USB_ADBUS[2]_net_1\, 
        \WR_USB_ADBUS[3]_net_1\, \WR_USB_ADBUS[4]_net_1\, 
        \WR_USB_ADBUS[5]_net_1\, \WR_USB_ADBUS[6]_net_1\, 
        \WR_USB_ADBUS[7]_net_1\, \ELINK_ADDRA_1[0]_net_1\, 
        \ELINK_ADDRA_1[1]_net_1\, \ELINK_ADDRA_1[2]_net_1\, 
        \ELINK_ADDRA_1[3]_net_1\, \ELINK_ADDRA_1[4]_net_1\, 
        \ELINK_ADDRA_1[5]_net_1\, \ELINK_ADDRA_1[6]_net_1\, 
        \ELINK_ADDRA_1[7]_net_1\, \ELINK_ADDRA_0[0]_net_1\, 
        \ELINK_ADDRA_0[1]_net_1\, \ELINK_ADDRA_0[2]_net_1\, 
        \ELINK_ADDRA_0[3]_net_1\, \ELINK_ADDRA_0[4]_net_1\, 
        \ELINK_ADDRA_0[5]_net_1\, \ELINK_ADDRA_0[6]_net_1\, 
        \ELINK_ADDRA_0[7]_net_1\, \TFC_DINA[0]_net_1\, 
        \TFC_DINA[1]_net_1\, \TFC_DINA[2]_net_1\, 
        \TFC_DINA[3]_net_1\, \TFC_DINA[4]_net_1\, 
        \TFC_DINA[5]_net_1\, \TFC_DINA[6]_net_1\, 
        \TFC_DINA[7]_net_1\, \ELINK_DINA_19[0]_net_1\, 
        \ELINK_DINA_19[1]_net_1\, \ELINK_DINA_19[2]_net_1\, 
        \ELINK_DINA_19[3]_net_1\, \ELINK_DINA_19[4]_net_1\, 
        \ELINK_DINA_19[5]_net_1\, \ELINK_DINA_19[6]_net_1\, 
        \ELINK_DINA_19[7]_net_1\, \ELINK_DINA_18[0]_net_1\, 
        \ELINK_DINA_18[1]_net_1\, \ELINK_DINA_18[2]_net_1\, 
        \ELINK_DINA_18[3]_net_1\, \ELINK_DINA_18[4]_net_1\, 
        \ELINK_DINA_18[5]_net_1\, \ELINK_DINA_18[6]_net_1\, 
        \ELINK_DINA_18[7]_net_1\, \ELINK_DINA_17[0]_net_1\, 
        \ELINK_DINA_17[1]_net_1\, \ELINK_DINA_17[2]_net_1\, 
        \ELINK_DINA_17[3]_net_1\, \ELINK_DINA_17[4]_net_1\, 
        \ELINK_DINA_17[5]_net_1\, \ELINK_DINA_17[6]_net_1\, 
        \ELINK_DINA_17[7]_net_1\, \ELINK_DINA_16[0]_net_1\, 
        \ELINK_DINA_16[1]_net_1\, \ELINK_DINA_16[2]_net_1\, 
        \ELINK_DINA_16[3]_net_1\, \ELINK_DINA_16[4]_net_1\, 
        \ELINK_DINA_16[5]_net_1\, \ELINK_DINA_16[6]_net_1\, 
        \ELINK_DINA_16[7]_net_1\, \ELINK_DINA_15[0]_net_1\, 
        \ELINK_DINA_15[1]_net_1\, \ELINK_DINA_15[2]_net_1\, 
        \ELINK_DINA_15[3]_net_1\, \ELINK_DINA_15[4]_net_1\, 
        \ELINK_DINA_15[5]_net_1\, \ELINK_DINA_15[6]_net_1\, 
        \ELINK_DINA_15[7]_net_1\, \ELINK_DINA_14[0]_net_1\, 
        \ELINK_DINA_14[1]_net_1\, \ELINK_DINA_14[2]_net_1\, 
        \ELINK_DINA_14[3]_net_1\, \ELINK_DINA_14[4]_net_1\, 
        \ELINK_DINA_14[5]_net_1\, \ELINK_DINA_14[6]_net_1\, 
        \ELINK_DINA_14[7]_net_1\, \ELINK_DINA_13[0]_net_1\, 
        \ELINK_DINA_13[1]_net_1\, \ELINK_DINA_13[2]_net_1\, 
        \ELINK_DINA_13[3]_net_1\, \ELINK_DINA_13[4]_net_1\, 
        \ELINK_DINA_13[5]_net_1\, \ELINK_DINA_13[6]_net_1\, 
        \ELINK_DINA_13[7]_net_1\, \ELINK_DINA_12[0]_net_1\, 
        \ELINK_DINA_12[1]_net_1\, \ELINK_DINA_12[2]_net_1\, 
        \ELINK_DINA_12[3]_net_1\, \ELINK_DINA_12[4]_net_1\, 
        \ELINK_DINA_12[5]_net_1\, \ELINK_DINA_12[6]_net_1\, 
        \ELINK_DINA_12[7]_net_1\, \ELINK_DINA_11[0]_net_1\, 
        \ELINK_DINA_11[1]_net_1\, \ELINK_DINA_11[2]_net_1\, 
        \ELINK_DINA_11[3]_net_1\, \ELINK_DINA_11[4]_net_1\, 
        \ELINK_DINA_11[5]_net_1\, \ELINK_DINA_11[6]_net_1\, 
        \ELINK_DINA_11[7]_net_1\, \ELINK_DINA_10[0]_net_1\, 
        \ELINK_DINA_10[1]_net_1\, \ELINK_DINA_10[2]_net_1\, 
        \ELINK_DINA_10[3]_net_1\, \ELINK_DINA_10[4]_net_1\, 
        \ELINK_DINA_10[5]_net_1\, \ELINK_DINA_10[6]_net_1\, 
        \ELINK_DINA_10[7]_net_1\, \ELINK_DINA_9[0]_net_1\, 
        \ELINK_DINA_9[1]_net_1\, \ELINK_DINA_9[2]_net_1\, 
        \ELINK_DINA_9[3]_net_1\, \ELINK_DINA_9[4]_net_1\, 
        \ELINK_DINA_9[5]_net_1\, \ELINK_DINA_9[6]_net_1\, 
        \ELINK_DINA_9[7]_net_1\, \ELINK_ADDRA_16[0]_net_1\, 
        \ELINK_ADDRA_16[1]_net_1\, \ELINK_ADDRA_16[2]_net_1\, 
        \ELINK_ADDRA_16[3]_net_1\, \ELINK_ADDRA_16[4]_net_1\, 
        \ELINK_ADDRA_16[5]_net_1\, \ELINK_ADDRA_16[6]_net_1\, 
        \ELINK_ADDRA_16[7]_net_1\, \ELINK_ADDRA_15[0]_net_1\, 
        \ELINK_ADDRA_15[1]_net_1\, \ELINK_ADDRA_15[2]_net_1\, 
        \ELINK_ADDRA_15[3]_net_1\, \ELINK_ADDRA_15[4]_net_1\, 
        \ELINK_ADDRA_15[5]_net_1\, \ELINK_ADDRA_15[6]_net_1\, 
        \ELINK_ADDRA_15[7]_net_1\, \ELINK_ADDRA_14[0]_net_1\, 
        \ELINK_ADDRA_14[1]_net_1\, \ELINK_ADDRA_14[2]_net_1\, 
        \ELINK_ADDRA_14[3]_net_1\, \ELINK_ADDRA_14[4]_net_1\, 
        \ELINK_ADDRA_14[5]_net_1\, \ELINK_ADDRA_14[6]_net_1\, 
        \ELINK_ADDRA_14[7]_net_1\, \ELINK_ADDRA_13[0]_net_1\, 
        \ELINK_ADDRA_13[1]_net_1\, \ELINK_ADDRA_13[2]_net_1\, 
        \ELINK_ADDRA_13[3]_net_1\, \ELINK_ADDRA_13[4]_net_1\, 
        \ELINK_ADDRA_13[5]_net_1\, \ELINK_ADDRA_13[6]_net_1\, 
        \ELINK_ADDRA_13[7]_net_1\, \ELINK_ADDRA_12[0]_net_1\, 
        \ELINK_ADDRA_12[1]_net_1\, \ELINK_ADDRA_12[2]_net_1\, 
        \ELINK_ADDRA_12[3]_net_1\, \ELINK_ADDRA_12[4]_net_1\, 
        \ELINK_ADDRA_12[5]_net_1\, \ELINK_ADDRA_12[6]_net_1\, 
        \ELINK_ADDRA_12[7]_net_1\, \ELINK_ADDRA_11[0]_net_1\, 
        \ELINK_ADDRA_11[1]_net_1\, \ELINK_ADDRA_11[2]_net_1\, 
        \ELINK_ADDRA_11[3]_net_1\, \ELINK_ADDRA_11[4]_net_1\, 
        \ELINK_ADDRA_11[5]_net_1\, \ELINK_ADDRA_11[6]_net_1\, 
        \ELINK_ADDRA_11[7]_net_1\, \ELINK_ADDRA_10[0]_net_1\, 
        \ELINK_ADDRA_10[1]_net_1\, \ELINK_ADDRA_10[2]_net_1\, 
        \ELINK_ADDRA_10[3]_net_1\, \ELINK_ADDRA_10[4]_net_1\, 
        \ELINK_ADDRA_10[5]_net_1\, \ELINK_ADDRA_10[6]_net_1\, 
        \ELINK_ADDRA_10[7]_net_1\, \ELINK_ADDRA_9[0]_net_1\, 
        \ELINK_ADDRA_9[1]_net_1\, \ELINK_ADDRA_9[2]_net_1\, 
        \ELINK_ADDRA_9[3]_net_1\, \ELINK_ADDRA_9[4]_net_1\, 
        \ELINK_ADDRA_9[5]_net_1\, \ELINK_ADDRA_9[6]_net_1\, 
        \ELINK_ADDRA_9[7]_net_1\, \ELINK_ADDRA_8[0]_net_1\, 
        \ELINK_ADDRA_8[1]_net_1\, \ELINK_ADDRA_8[2]_net_1\, 
        \ELINK_ADDRA_8[3]_net_1\, \ELINK_ADDRA_8[4]_net_1\, 
        \ELINK_ADDRA_8[5]_net_1\, \ELINK_ADDRA_8[6]_net_1\, 
        \ELINK_ADDRA_8[7]_net_1\, \ELINK_ADDRA_7[0]_net_1\, 
        \ELINK_ADDRA_7[1]_net_1\, \ELINK_ADDRA_7[2]_net_1\, 
        \ELINK_ADDRA_7[3]_net_1\, \ELINK_ADDRA_7[4]_net_1\, 
        \ELINK_ADDRA_7[5]_net_1\, \ELINK_ADDRA_7[6]_net_1\, 
        \ELINK_ADDRA_7[7]_net_1\, \ELINK_ADDRA_6[0]_net_1\, 
        \ELINK_ADDRA_6[1]_net_1\, \ELINK_ADDRA_6[2]_net_1\, 
        \ELINK_ADDRA_6[3]_net_1\, \ELINK_ADDRA_6[4]_net_1\, 
        \ELINK_ADDRA_6[5]_net_1\, \ELINK_ADDRA_6[6]_net_1\, 
        \ELINK_ADDRA_6[7]_net_1\, \ELINK_ADDRA_5[0]_net_1\, 
        \ELINK_ADDRA_5[1]_net_1\, \ELINK_ADDRA_5[2]_net_1\, 
        \ELINK_ADDRA_5[3]_net_1\, \ELINK_ADDRA_5[4]_net_1\, 
        \ELINK_ADDRA_5[5]_net_1\, \ELINK_ADDRA_5[6]_net_1\, 
        \ELINK_ADDRA_5[7]_net_1\, \ELINK_ADDRA_4[0]_net_1\, 
        \ELINK_ADDRA_4[1]_net_1\, \ELINK_ADDRA_4[2]_net_1\, 
        \ELINK_ADDRA_4[3]_net_1\, \ELINK_ADDRA_4[4]_net_1\, 
        \ELINK_ADDRA_4[5]_net_1\, \ELINK_ADDRA_4[6]_net_1\, 
        \ELINK_ADDRA_4[7]_net_1\, \ELINK_ADDRA_3[0]_net_1\, 
        \ELINK_ADDRA_3[1]_net_1\, \ELINK_ADDRA_3[2]_net_1\, 
        \ELINK_ADDRA_3[3]_net_1\, \ELINK_ADDRA_3[4]_net_1\, 
        \ELINK_ADDRA_3[5]_net_1\, \ELINK_ADDRA_3[6]_net_1\, 
        \ELINK_ADDRA_3[7]_net_1\, \ELINK_ADDRA_2[0]_net_1\, 
        \ELINK_ADDRA_2[1]_net_1\, \ELINK_ADDRA_2[2]_net_1\, 
        \ELINK_ADDRA_2[3]_net_1\, \ELINK_ADDRA_2[4]_net_1\, 
        \ELINK_ADDRA_2[5]_net_1\, \ELINK_ADDRA_2[6]_net_1\, 
        \ELINK_ADDRA_2[7]_net_1\, \TFC_ADDRA[0]_net_1\, 
        \TFC_ADDRA[1]_net_1\, \TFC_ADDRA[2]_net_1\, 
        \TFC_ADDRA[3]_net_1\, \TFC_ADDRA[4]_net_1\, 
        \TFC_ADDRA[5]_net_1\, \TFC_ADDRA[6]_net_1\, 
        \TFC_ADDRA[7]_net_1\, \ELINK_ADDRA_19[0]_net_1\, 
        \ELINK_ADDRA_19[1]_net_1\, \ELINK_ADDRA_19[2]_net_1\, 
        \ELINK_ADDRA_19[3]_net_1\, \ELINK_ADDRA_19[4]_net_1\, 
        \ELINK_ADDRA_19[5]_net_1\, \ELINK_ADDRA_19[6]_net_1\, 
        \ELINK_ADDRA_19[7]_net_1\, \ELINK_ADDRA_18[0]_net_1\, 
        \ELINK_ADDRA_18[1]_net_1\, \ELINK_ADDRA_18[2]_net_1\, 
        \ELINK_ADDRA_18[3]_net_1\, \ELINK_ADDRA_18[4]_net_1\, 
        \ELINK_ADDRA_18[5]_net_1\, \ELINK_ADDRA_18[6]_net_1\, 
        \ELINK_ADDRA_18[7]_net_1\, \ELINK_ADDRA_17[0]_net_1\, 
        \ELINK_ADDRA_17[1]_net_1\, \ELINK_ADDRA_17[2]_net_1\, 
        \ELINK_ADDRA_17[3]_net_1\, \ELINK_ADDRA_17[4]_net_1\, 
        \ELINK_ADDRA_17[5]_net_1\, \ELINK_ADDRA_17[6]_net_1\, 
        \ELINK_ADDRA_17[7]_net_1\, \N_RD_USB_ADBUS[0]\, 
        \N_RD_USB_ADBUS[1]\, \N_RD_USB_ADBUS[2]\, 
        \N_RD_USB_ADBUS[3]\, \N_RD_USB_ADBUS[4]\, 
        \N_RD_USB_ADBUS[5]\, \N_RD_USB_ADBUS[6]\, 
        \N_RD_USB_ADBUS[7]\, \OP_MODE_0[0]\, \OP_MODE_0[4]\, 
        \GND\, \VCC\ : std_logic;

    for all : DPRT_512X9_SRAM_0
	Use entity work.DPRT_512X9_SRAM_0(DEF_ARCH);
    for all : DPRT_512X9_SRAM_13
	Use entity work.DPRT_512X9_SRAM_13(DEF_ARCH);
    for all : DPRT_512X9_SRAM_12
	Use entity work.DPRT_512X9_SRAM_12(DEF_ARCH);
    for all : DPRT_512X9_SRAM_11
	Use entity work.DPRT_512X9_SRAM_11(DEF_ARCH);
    for all : DPRT_512X9_SRAM_16
	Use entity work.DPRT_512X9_SRAM_16(DEF_ARCH);
    for all : CLK60M_TO_40M_4_1
	Use entity work.CLK60M_TO_40M_4_1(DEF_ARCH);
    for all : DPRT_512X9_SRAM_3
	Use entity work.DPRT_512X9_SRAM_3(DEF_ARCH);
    for all : DPRT_512X9_SRAM_2
	Use entity work.DPRT_512X9_SRAM_2(DEF_ARCH);
    for all : DPRT_512X9_SRAM_1
	Use entity work.DPRT_512X9_SRAM_1(DEF_ARCH);
    for all : DPRT_512X9_SRAM_6
	Use entity work.DPRT_512X9_SRAM_6(DEF_ARCH);
    for all : CLK60M_TO_40M_0
	Use entity work.CLK60M_TO_40M_0(DEF_ARCH);
    for all : BIDIR_LVTTL
	Use entity work.BIDIR_LVTTL(DEF_ARCH);
    for all : DPRT_512X9_SRAM_14
	Use entity work.DPRT_512X9_SRAM_14(DEF_ARCH);
    for all : DPRT_512X9_SRAM_17
	Use entity work.DPRT_512X9_SRAM_17(DEF_ARCH);
    for all : CLK60M_TO_40M_4_2
	Use entity work.CLK60M_TO_40M_4_2(DEF_ARCH);
    for all : CLK60M_TO_40M_4_0
	Use entity work.CLK60M_TO_40M_4_0(DEF_ARCH);
    for all : DPRT_512X9_SRAM_4
	Use entity work.DPRT_512X9_SRAM_4(DEF_ARCH);
    for all : DPRT_512X9_SRAM_19
	Use entity work.DPRT_512X9_SRAM_19(DEF_ARCH);
    for all : DPRT_512X9_SRAM_7
	Use entity work.DPRT_512X9_SRAM_7(DEF_ARCH);
    for all : CLK60M_TO_40M_4
	Use entity work.CLK60M_TO_40M_4(DEF_ARCH);
    for all : DPRT_512X9_SRAM_9
	Use entity work.DPRT_512X9_SRAM_9(DEF_ARCH);
    for all : DPRT_512X9_SRAM_18
	Use entity work.DPRT_512X9_SRAM_18(DEF_ARCH);
    for all : DPRT_512X9_SRAM_15
	Use entity work.DPRT_512X9_SRAM_15(DEF_ARCH);
    for all : DPRT_512X9_SRAM
	Use entity work.DPRT_512X9_SRAM(DEF_ARCH);
    for all : DPRT_512X9_SRAM_10
	Use entity work.DPRT_512X9_SRAM_10(DEF_ARCH);
    for all : DPRT_512X9_SRAM_8
	Use entity work.DPRT_512X9_SRAM_8(DEF_ARCH);
    for all : DPRT_512X9_SRAM_5
	Use entity work.DPRT_512X9_SRAM_5(DEF_ARCH);
begin 

    OP_MODE_0_0 <= \OP_MODE_0[0]\;
    OP_MODE_0_4 <= \OP_MODE_0[4]\;

    \TFC_ADDRA[4]\ : DFN1E0C0
      port map(D => \N_TFC_ADDRA[4]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_9, E => N_142, Q => 
        \TFC_ADDRA[4]_net_1\);
    
    \SM_BANK_SEL_RNIJ57M1[8]\ : OR3C
      port map(A => N_477, B => N_365, C => N_143, Y => 
        \N_ELINK_RWA_1[12]\);
    
    \RD_USB_ADBUS_RNIFM0T[7]\ : NOR2A
      port map(A => N_1351_4, B => \RD_USB_ADBUS[7]_net_1\, Y => 
        N_465);
    
    \WR_USB_ADBUS_RNO_4[0]\ : AO1
      port map(A => \ELINK_DOUTA_8[0]\, B => un1_SM_BANK_SEL_38, 
        C => \ELINK_DOUTA_9_m[0]\, Y => 
        \N_WR_USB_ADBUS_0_iv_9[0]\);
    
    \TFC_ADDRA[7]\ : DFN1E0C0
      port map(D => \N_TFC_ADDRA[7]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_10, E => N_142, Q => 
        \TFC_ADDRA[7]_net_1\);
    
    \ELINK_RWA_RNO[18]\ : AOI1
      port map(A => \SM_BANK_SEL[1]_net_1\, B => un1_USB_RXF_B_m, 
        C => N_171, Y => \N_ELINK_RWA_0_iv[18]\);
    
    \WR_USB_ADBUS_RNO_16[2]\ : AO1
      port map(A => \ELINK_DOUTA_6[2]\, B => un1_SM_BANK_SEL_30, 
        C => \ELINK_DOUTA_7_m[2]\, Y => 
        \N_WR_USB_ADBUS_0_iv_8[2]\);
    
    \SI_CNT_RNI1PT8[1]\ : NOR2B
      port map(A => \SI_CNT[0]_net_1\, B => \SI_CNT[1]_net_1\, Y
         => N_2607);
    
    \ELINK_BLKA_RNO_0[17]\ : NOR2B
      port map(A => \SM_BANK_SEL[2]_net_1\, B => X_BLKA_i, Y => 
        X_BLKA_i_m_16);
    
    \WR_USB_ADBUS_RNO_6[4]\ : AO1
      port map(A => \ELINK_DOUTA_6[4]\, B => un1_SM_BANK_SEL_30, 
        C => \ELINK_DOUTA_7_m[4]\, Y => 
        \N_WR_USB_ADBUS_0_iv_8[4]\);
    
    \TFC_DINA[5]\ : DFN1E0C0
      port map(D => \N_TFC_DINA[5]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_4, E => N_142, Q => \TFC_DINA[5]_net_1\);
    
    \SM_BANK_SEL_RNIE4P72[2]\ : NOR3A
      port map(A => \SM_BANK_SEL[2]_net_1\, B => N_312, C => 
        N_1566_i_i_0, Y => un1_SM_BANK_SEL_40);
    
    \ELINK_DINA_0[1]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[1]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_5, E => un1_SM_BANK_SEL_6, Q => 
        \ELINK_DINA_0[1]_net_1\);
    
    \WR_USB_ADBUS_RNO_10[4]\ : AO1A
      port map(A => N_243, B => \TFC_DOUTA[4]\, C => 
        \ELINK_DOUTA_15_m[4]\, Y => \N_WR_USB_ADBUS_0_iv_13[4]\);
    
    \WR_USB_ADBUS_RNO_15[4]\ : NOR2B
      port map(A => \ELINK_DOUTA_12[4]\, B => un1_SM_BANK_SEL_33, 
        Y => \ELINK_DOUTA_12_m[4]\);
    
    \WR_USB_ADBUS_RNO_10[0]\ : AO1A
      port map(A => N_243, B => \TFC_DOUTA[0]\, C => 
        \ELINK_DOUTA_15_m[0]\, Y => \N_WR_USB_ADBUS_0_iv_13[0]\);
    
    \REG_STATE_RNIUON31[0]\ : NOR2B
      port map(A => N_1690_i, B => \REG_STATE[0]_net_1\, Y => 
        N_1891);
    
    \ELINK_DINA_18[3]\ : DFN1E0C0
      port map(D => \N_TFC_DINA[3]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_21, E => N_198, Q => 
        \ELINK_DINA_18[3]_net_1\);
    
    \REG_STATE_0_RNITRSJ1[0]\ : NOR3A
      port map(A => N_2477_i, B => \REG_STATE_0[1]_net_1\, C => 
        \REG_STATE_0[0]_net_1\, Y => N_2561);
    
    \ELINK_DINA_17[5]\ : DFN1E0C0
      port map(D => \N_TFC_DINA[5]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_19, E => N_197, Q => 
        \ELINK_DINA_17[5]_net_1\);
    
    \WR_USB_ADBUS_RNO_7[1]\ : NOR2B
      port map(A => \ELINK_DOUTA_14[1]\, B => un1_SM_BANK_SEL_23, 
        Y => \ELINK_DOUTA_14_m[1]\);
    
    \RD_USB_ADBUS[1]\ : DFN1C0
      port map(D => \N_RD_USB_ADBUS[1]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_22, Q => \RD_USB_ADBUS[1]_net_1\);
    
    \ELINK_BLKA_RNO_0[5]\ : OA1B
      port map(A => N_616_16, B => \N_ELINK_RWA_3[5]\, C => 
        \ELINK_BLKA[5]_net_1\, Y => N_165);
    
    \SM_BANK_SEL_RNO[2]\ : NOR3B
      port map(A => un1_N_ELK_N_ACTIVE_0_sqmuxa_15_0_a2_0_0, B
         => N_1351_4, C => N_1697, Y => N_1840);
    
    \ELINK_RWA_RNO[4]\ : AOI1
      port map(A => \SM_BANK_SEL[15]_net_1\, B => un1_USB_RXF_B_m, 
        C => \ELINK_RWA_i_m[4]\, Y => \N_ELINK_RWA_0_iv[4]\);
    
    \SM_BANK_SEL_RNIQ1VN[19]\ : OR3A
      port map(A => N_143, B => N_616_11, C => \N_ELINK_RWA_1[1]\, 
        Y => \N_ELINK_RWA_3[1]\);
    
    \WR_USB_ADBUS_RNO_31[4]\ : NOR3B
      port map(A => N_1730_i, B => \ELINKS_STOP_ADDR[4]_net_1\, C
         => N_1726, Y => \ELINKS_STOP_ADDR_m[4]\);
    
    \WR_USB_ADBUS_RNO_16[7]\ : AO1
      port map(A => \ELINK_DOUTA_4[7]\, B => un1_SM_BANK_SEL_28, 
        C => \ELINK_DOUTA_5_m[7]\, Y => 
        \N_WR_USB_ADBUS_0_iv_12[7]\);
    
    \RD_USB_ADBUS[5]\ : DFN1C0
      port map(D => \N_RD_USB_ADBUS[5]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_22, Q => \RD_USB_ADBUS[5]_net_1\);
    
    \RD_USB_ADBUS[2]\ : DFN1C0
      port map(D => \N_RD_USB_ADBUS[2]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_22, Q => \RD_USB_ADBUS[2]_net_1\);
    
    \ELINK_DINA_16[7]\ : DFN1E0C0
      port map(D => \N_TFC_DINA[7]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_18, E => N_200, Q => 
        \ELINK_DINA_16[7]_net_1\);
    
    \REG_ADDR_RNO[8]\ : XA1B
      port map(A => REG_ADDR_75_0, B => \REG_ADDR[8]_net_1\, C
         => N_675_0, Y => REG_ADDR_n8);
    
    \WR_USB_ADBUS_RNO_4[2]\ : NOR2B
      port map(A => \ELINK_DOUTA_1[2]\, B => un1_SM_BANK_SEL_36, 
        Y => \ELINK_DOUTA_1_m[2]\);
    
    \ELINK_ADDRA_17[4]\ : DFN1E0C0
      port map(D => \N_TFC_ADDRA[4]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_11, E => N_197, Q => 
        \ELINK_ADDRA_17[4]_net_1\);
    
    \REG_STATE_ns_i_i_o2_1_RNO_4[0]\ : NOR3B
      port map(A => \REG_STATE_0[3]_net_1\, B => N_1499_2_i_0, C
         => \USB_TXE_B\, Y => N_439);
    
    \ELINK_ADDRA_9[3]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[3]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_10, E => un1_SM_BANK_SEL_9, Q => 
        \ELINK_ADDRA_9[3]_net_1\);
    
    \REG_STATE_RNIMO53U3[2]\ : NOR3
      port map(A => \REG_STATE_ns_i_3[4]\, B => 
        \REG_STATE_ns_i_6[4]\, C => \REG_STATE_ns_i_4[4]\, Y => 
        \REG_STATE_RNIMO53U3[2]_net_1\);
    
    \REG_ADDR_RNI1O7P2[2]\ : AO1
      port map(A => N_1398_i_0_a2_3, B => N_474, C => N_252, Y
         => N_1398_i_0_0);
    
    \ELINK_DINA_10[0]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[0]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_9, E => un1_SM_BANK_SEL_20, Q => 
        \ELINK_DINA_10[0]_net_1\);
    
    \ELINK_DINA_9[4]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[4]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_20, E => un1_SM_BANK_SEL_9, Q => 
        \ELINK_DINA_9[4]_net_1\);
    
    \ELINK_RWA[4]\ : DFN1E0P0
      port map(D => \N_ELINK_RWA_0_iv[4]\, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_6, E => \SM_BANK_SEL_0[20]_net_1\, 
        Q => \ELINK_RWA[4]_net_1\);
    
    \ELINK_DINA_2[6]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[6]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_9, E => un1_SM_BANK_SEL_5, Q => 
        \ELINK_DINA_2[6]_net_1\);
    
    \WR_XFER_TYPE_RNI4KSS_0[7]\ : NOR2A
      port map(A => \WR_XFER_TYPE[7]_net_1\, B => 
        \WR_XFER_TYPE[1]_net_1\, Y => REG_STATE_tr67_1);
    
    \SM_BANK_SEL_RNI8BHH[3]\ : NOR3
      port map(A => \SM_BANK_SEL[6]_net_1\, B => 
        \SM_BANK_SEL[5]_net_1\, C => \SM_BANK_SEL[3]_net_1\, Y
         => \N_ELINK_RWA_0_iv_0_o2_i_a5_0[15]\);
    
    \ELINK_DINA_10[4]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[4]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_9, E => un1_SM_BANK_SEL_20, Q => 
        \ELINK_DINA_10[4]_net_1\);
    
    \REG_STATE_0_RNI1JQ94[4]\ : OR3A
      port map(A => \REG_STATE_0[4]_net_1\, B => N_2577, C => 
        \REG_STATE_ns_i_tz_0[5]\, Y => \REG_STATE_ns_i_tz_1[5]\);
    
    REG_STATE_s23_i_2 : OR2
      port map(A => REG_STATE_s23_i_1, B => REG_STATE_s23_i_0, Y
         => \REG_STATE_s23_i_2\);
    
    USB_RXF_B_0_RNI3CDL61 : OA1
      port map(A => \REG_STATE_ns_i_a4_8_0_a5_0[4]\, B => 
        \REG_STATE_ns_i_a4_6_1[4]\, C => N_2597, Y => 
        \REG_STATE_ns_i_6[4]\);
    
    \ELINK_RWA[11]\ : DFN1E0P0
      port map(D => \N_ELINK_RWA_0_iv[11]\, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_11, E => \SM_BANK_SEL_0[20]_net_1\, 
        Q => \ELINK_RWA[11]_net_1\);
    
    \ELINK_DINA_5[6]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[6]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_14, E => un1_SM_BANK_SEL_15, Q => 
        \ELINK_DINA_5[6]_net_1\);
    
    \REG_STATE_RNIU1LF1[2]\ : NOR2A
      port map(A => N_470, B => \REG_STATE[2]_net_1\, Y => N_504);
    
    \SM_BANK_SEL_RNO[7]\ : NOR3C
      port map(A => \RD_USB_ADBUS[2]_net_1\, B => N_1892, C => 
        N_1902, Y => N_1842);
    
    \WR_USB_ADBUS_RNO_31[7]\ : AO1C
      port map(A => N_1499, B => \ELINKS_STRT_ADDR[7]_net_1\, C
         => N_1569, Y => \N_WR_USB_ADBUS_0_iv_1[7]\);
    
    \WR_USB_ADBUS_RNO_6[1]\ : OR3
      port map(A => \N_WR_USB_ADBUS_0_iv_3[1]\, B => 
        \N_WR_USB_ADBUS_0_iv_2[1]\, C => 
        \N_WR_USB_ADBUS_0_iv_4[1]\, Y => 
        \N_WR_USB_ADBUS_0_iv_6[1]\);
    
    \SM_BANK_SEL_RNO[6]\ : NOR3C
      port map(A => \RD_USB_ADBUS[2]_net_1\, B => N_1892, C => 
        N_1351_4, Y => N_1837);
    
    \REG_STATE_RNI2KQN_0[4]\ : NOR2
      port map(A => \REG_STATE[4]_net_1\, B => 
        \REG_STATE[2]_net_1\, Y => N_1877_1);
    
    \ELINK_BLKA_RNO[3]\ : AOI1
      port map(A => \SM_BANK_SEL[16]_net_1\, B => X_BLKA_i, C => 
        \ELINK_BLKA_i_m[3]\, Y => \N_ELINK_BLKA_0_iv[3]\);
    
    USB_RXF_B_0_RNICKDL2 : NOR2B
      port map(A => N_1730_i, B => N_1907, Y => 
        N_ELINKS_STRT_ADDR_T_0_sqmuxa);
    
    \OP_MODE_T[1]\ : DFN1E1C0
      port map(D => \RD_USB_ADBUS[1]_net_1\, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_17, E => N_OP_MODE_T_0_sqmuxa, Q
         => \OP_MODE_T[1]_net_1\);
    
    \WR_USB_ADBUS_RNO_23[6]\ : NOR2B
      port map(A => \ELINK_DOUTA_12[6]\, B => un1_SM_BANK_SEL_33, 
        Y => \ELINK_DOUTA_12_m[6]\);
    
    \REG_STATE_RNITNN31[1]\ : NOR2A
      port map(A => N_1710_i_0, B => \REG_STATE[1]_net_1\, Y => 
        N_1745_i);
    
    \ELINK_DINA_14[4]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[4]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_16, E => un1_SM_BANK_SEL_1, Q => 
        \ELINK_DINA_14[4]_net_1\);
    
    \ELINK_DINA_13[0]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[0]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_14, E => un1_SM_BANK_SEL_2, Q => 
        \ELINK_DINA_13[0]_net_1\);
    
    \REG_ADDR_RNIOTCP[5]\ : NOR3B
      port map(A => N_261, B => \REG_ADDR[5]_net_1\, C => 
        \SM_BANK_SEL_0[21]_net_1\, Y => \N_TFC_ADDRA[5]\);
    
    \ELINK_ADDRA_12[6]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[6]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_2_0, E => un1_SM_BANK_SEL_7, Q => 
        \ELINK_ADDRA_12[6]_net_1\);
    
    \ELINK_ADDRA_17[5]\ : DFN1E0C0
      port map(D => \N_TFC_ADDRA[5]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_11, E => N_197, Q => 
        \ELINK_ADDRA_17[5]_net_1\);
    
    \SI_CNT_RNI6MRH[3]\ : NOR2B
      port map(A => \REG_STATE_ns_i_a2_2_0[4]\, B => N_2607, Y
         => N_2613);
    
    \ELINK_RWA_RNO[16]\ : AOI1
      port map(A => \SM_BANK_SEL[3]_net_1\, B => un1_USB_RXF_B_m, 
        C => \ELINK_RWA_i_m[16]\, Y => \N_ELINK_RWA_0_iv[16]\);
    
    \REG_STATE_RNI5NQN_1[5]\ : NOR2
      port map(A => \REG_STATE[5]_net_1\, B => 
        \REG_STATE[4]_net_1\, Y => N_1351_3);
    
    \REG_STATE_0_RNIU5QV1[0]\ : XO1
      port map(A => \REG_STATE_0[2]_net_1\, B => 
        \REG_STATE_0[0]_net_1\, C => N_1691, Y => N_1703);
    
    \WR_USB_ADBUS_RNO_14[1]\ : NOR2B
      port map(A => \ELINK_DOUTA_3[1]\, B => un1_SM_BANK_SEL_43, 
        Y => \ELINK_DOUTA_3_m[1]\);
    
    \ELINK_ADDRA_18[2]\ : DFN1E0C0
      port map(D => \N_TFC_ADDRA[2]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_12, E => N_198, Q => 
        \ELINK_ADDRA_18[2]_net_1\);
    
    \ELINK_ADDRA_19[1]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[1]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_13, E => un1_SM_BANK_SEL_11, Q => 
        \ELINK_ADDRA_19[1]_net_1\);
    
    \ELINK_ADDRA_17[3]\ : DFN1E0C0
      port map(D => \N_TFC_ADDRA[3]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_10, E => N_197, Q => 
        \ELINK_ADDRA_17[3]_net_1\);
    
    \REG_STATE[2]\ : DFN1C0
      port map(D => \REG_STATE_RNIVPG2K2[2]_net_1\, CLK => 
        CLK60MHZ, CLR => P_USB_MASTER_EN_c_22_0, Q => 
        \REG_STATE[2]_net_1\);
    
    \ELINK_ADDRA_4[5]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[5]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_2_0, E => un1_SM_BANK_SEL_8, Q => 
        \ELINK_ADDRA_4[5]_net_1\);
    
    \TFC_STRT_ADDR[4]\ : DFN1E1C0
      port map(D => \TFC_STRT_ADDR_T[4]_net_1\, CLK => CLK60MHZ, 
        CLR => P_USB_MASTER_EN_c_13, E => \REG_STATE_d_0[30]\, Q
         => \TFC_STRT_ADDR[4]_net_1\);
    
    \SM_BANK_SEL_RNITVGH[1]\ : NOR2A
      port map(A => N_463, B => \SM_BANK_SEL[1]_net_1\, Y => 
        N_143);
    
    \ELINK_ADDRA_14[5]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[5]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_5, E => un1_SM_BANK_SEL_1, Q => 
        \ELINK_ADDRA_14[5]_net_1\);
    
    \ELINK_DINA_6[2]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[2]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_16, E => un1_SM_BANK_SEL_10, Q => 
        \ELINK_DINA_6[2]_net_1\);
    
    \WR_XFER_TYPE_RNO_1[2]\ : NOR2A
      port map(A => N_1716, B => \WR_XFER_TYPE[2]_net_1\, Y => 
        N_1822);
    
    \ELINK_DINA_6[6]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[6]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_16, E => un1_SM_BANK_SEL_10, Q => 
        \ELINK_DINA_6[6]_net_1\);
    
    \ELINK_DINA_8[3]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[3]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_18, E => un1_SM_BANK_SEL_21, Q => 
        \ELINK_DINA_8[3]_net_1\);
    
    \N_WR_USB_ADBUS_0_iv_0_RNO[6]\ : NOR2A
      port map(A => \TFC_STOP_ADDR[6]_net_1\, B => N_1501, Y => 
        \TFC_STOP_ADDR_m[6]\);
    
    \ELINK_DINA_3[2]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[2]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_11, E => un1_SM_BANK_SEL_4, Q => 
        \ELINK_DINA_3[2]_net_1\);
    
    \ELINK_ADDRA_9[5]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[5]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_10, E => un1_SM_BANK_SEL_9, Q => 
        \ELINK_ADDRA_9[5]_net_1\);
    
    \TFC_STOP_ADDR[2]\ : DFN1E1C0
      port map(D => \TFC_STOP_ADDR_T[2]_net_1\, CLK => CLK60MHZ, 
        CLR => P_USB_MASTER_EN_c_8, E => \REG_STATE_d_0[30]\, Q
         => \TFC_STOP_ADDR[2]_net_1\);
    
    USB_TXE_B_RNIPOIA1 : OR2A
      port map(A => \USB_TXE_B\, B => N_255, Y => N_256);
    
    \RD_XFER_TYPE[3]\ : DFN1C0
      port map(D => \RD_XFER_TYPE_RNO[3]_net_1\, CLK => CLK60MHZ, 
        CLR => P_USB_MASTER_EN_c, Q => \RD_XFER_TYPE[3]_net_1\);
    
    \RD_USB_ADBUS_RNI4OCD2[4]\ : OR2
      port map(A => N_1903, B => N_1698, Y => N_1736);
    
    \ELINK_ADDRA_1[0]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[0]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_20, E => un1_SM_BANK_SEL_19, Q => 
        \ELINK_ADDRA_1[0]_net_1\);
    
    \ELINK_BLKA_RNO_0[6]\ : NOR2B
      port map(A => \SM_BANK_SEL[13]_net_1\, B => X_BLKA_i, Y => 
        X_BLKA_i_m_5);
    
    \WR_XFER_TYPE_RNI4KSS[7]\ : NOR2B
      port map(A => \WR_XFER_TYPE[7]_net_1\, B => 
        \WR_XFER_TYPE[1]_net_1\, Y => REG_STATE_tr72_6_1);
    
    \ELINK_DINA_8[6]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[6]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_18, E => un1_SM_BANK_SEL_21, Q => 
        \ELINK_DINA_8[6]_net_1\);
    
    \WR_USB_ADBUS_RNO_13[2]\ : NOR2B
      port map(A => \ELINK_DOUTA_16[2]\, B => un1_SM_BANK_SEL_39, 
        Y => \ELINK_DOUTA_16_m[2]\);
    
    \ELINK_RWA_RNO[13]\ : AOI1
      port map(A => \SM_BANK_SEL[6]_net_1\, B => un1_USB_RXF_B_m, 
        C => N_177, Y => \N_ELINK_RWA_0_iv[13]\);
    
    \SM_BANK_SEL_RNIUNN22[11]\ : NOR3A
      port map(A => \SM_BANK_SEL[11]_net_1\, B => N_312, C => 
        N_1566_i_i_0, Y => un1_SM_BANK_SEL_38);
    
    \SM_BANK_SEL[4]\ : DFN1E1C0
      port map(D => N_1832, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_7, E => un1_REG_STATE_30, Q => 
        \SM_BANK_SEL[4]_net_1\);
    
    \WR_XFER_TYPE_RNO[3]\ : NOR3
      port map(A => N_1826, B => N_1823, C => N_1825, Y => 
        \WR_XFER_TYPE_RNO[3]_net_1\);
    
    \SM_BANK_SEL_RNIQC73[16]\ : OR2
      port map(A => \N_ELINK_BLKA_10_0[10]\, B => N_618_1, Y => 
        N_620_10);
    
    \SM_BANK_SEL_RNIMRK6[10]\ : OR2
      port map(A => \SM_BANK_SEL[10]_net_1\, B => 
        \SM_BANK_SEL[9]_net_1\, Y => \N_ELINK_RWA_16_0[0]\);
    
    USB_TXE_B_RNIIHIA1 : NOR2A
      port map(A => N_1352_1, B => N_339, Y => N_456);
    
    \TFC_DINA[7]\ : DFN1E0C0
      port map(D => \N_TFC_DINA[7]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_4, E => N_142, Q => \TFC_DINA[7]_net_1\);
    
    \WR_USB_ADBUS_RNO[2]\ : OR3
      port map(A => \N_WR_USB_ADBUS_0_iv_22[2]\, B => 
        \N_WR_USB_ADBUS_0_iv_21[2]\, C => 
        \N_WR_USB_ADBUS_0_iv_26[2]\, Y => \N_WR_USB_ADBUS[2]\);
    
    \ELINK_DINA_12[3]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[3]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_12, E => un1_SM_BANK_SEL_7, Q => 
        \ELINK_DINA_12[3]_net_1\);
    
    \REG_STATE_0[3]\ : DFN1C0
      port map(D => \REG_STATE_0_RNIGPV6T1[0]_net_1\, CLK => 
        CLK60MHZ, CLR => P_USB_MASTER_EN_c_22_0, Q => 
        \REG_STATE_0[3]_net_1\);
    
    \RD_USB_ADBUS_RNIMAIK2[1]\ : NOR2A
      port map(A => \RD_USB_ADBUS[1]_net_1\, B => N_206, Y => 
        \N_TFC_DINA[1]\);
    
    \N_WR_USB_ADBUS_0_iv_0[2]\ : OR2
      port map(A => \TFC_STOP_ADDR_m[2]\, B => N_1562_i, Y => 
        \N_WR_USB_ADBUS_0_iv_0[2]_net_1\);
    
    \REG_STATE_RNI0J4O4[5]\ : NOR3B
      port map(A => REG_STATE_tr49_6, B => N_1351_8, C => N_252, 
        Y => N_1374);
    
    \REG_ADDR_RNO[2]\ : NOR2
      port map(A => REG_ADDR_n2_i_0, B => N_675, Y => N_2629);
    
    \REG_STATE_ns_i_i_o2_6[0]\ : OR2
      port map(A => N_275, B => 
        \REG_STATE_ns_i_i_o2_6_1[0]_net_1\, Y => N_244_1);
    
    REG_STATE_s23_i_2_RNO : OR2A
      port map(A => \REG_STATE[3]_net_1\, B => 
        \REG_STATE[5]_net_1\, Y => REG_STATE_s23_i_1);
    
    \RD_USB_ADBUS_RNI38BJ_0[4]\ : NOR2A
      port map(A => \RD_USB_ADBUS[4]_net_1\, B => 
        \RD_USB_ADBUS[5]_net_1\, Y => N_459);
    
    \ELINK_ADDRA_8[4]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[4]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_8, E => un1_SM_BANK_SEL_21, Q => 
        \ELINK_ADDRA_8[4]_net_1\);
    
    \ELINK_RWA[9]\ : DFN1E0P0
      port map(D => \N_ELINK_RWA_0_iv[9]\, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_6, E => \SM_BANK_SEL_0[20]_net_1\, 
        Q => \ELINK_RWA[9]_net_1\);
    
    \WR_XFER_TYPE_RNI0FP34[5]\ : NOR3B
      port map(A => REG_STATE_tr67_3, B => N_1404_7, C => N_252, 
        Y => REG_STATE_tr67_5);
    
    \REG_STATE_0_RNI6NBS2[3]\ : AO1
      port map(A => N_2606, B => N_287, C => N_417, Y => 
        \REG_STATE_ns_i_i_o2_10_0[2]\);
    
    \REG_STATE_ns_i_i_a2_0_RNIN0TJ41[0]\ : OR3A
      port map(A => N_511_1, B => N_388, C => 
        \REG_STATE_ns_i_i_2[0]\, Y => 
        \REG_STATE_ns_i_i_a2_0_RNIN0TJ41[0]_net_1\);
    
    \REG_ADDR_RNITPKG2[1]\ : NOR3C
      port map(A => REG_STATE_tr49_3, B => REG_STATE_tr49_2, C
         => REG_STATE_tr49_4, Y => REG_STATE_tr49_6);
    
    \WR_USB_ADBUS_RNO_9[6]\ : AO1
      port map(A => \ELINK_DOUTA_0[6]\, B => un1_SM_BANK_SEL_31, 
        C => \ELINK_DOUTA_13_m[6]\, Y => 
        \N_WR_USB_ADBUS_0_iv_13[6]\);
    
    \SM_BANK_SEL_RNI08VN[13]\ : OR3A
      port map(A => N_143, B => N_620_10, C => \N_ELINK_RWA_1[7]\, 
        Y => \N_ELINK_RWA_3[7]\);
    
    USB_RXF_B_0_RNIE0VR9 : OR2
      port map(A => N_1419, B => N_1737, Y => un1_REG_STATE_30);
    
    \TFC_STRT_ADDR[3]\ : DFN1E1C0
      port map(D => \TFC_STRT_ADDR_T[3]_net_1\, CLK => CLK60MHZ, 
        CLR => P_USB_MASTER_EN_c_13, E => \REG_STATE_d_0[30]\, Q
         => \TFC_STRT_ADDR[3]_net_1\);
    
    \TFC_STOP_ADDR[7]\ : DFN1E1C0
      port map(D => \TFC_STOP_ADDR_T[7]_net_1\, CLK => CLK60MHZ, 
        CLR => P_USB_MASTER_EN_c_8, E => \REG_STATE_d_0[30]\, Q
         => \TFC_STOP_ADDR[7]_net_1\);
    
    \ELINKS_STRT_ADDR[4]\ : DFN1E1C0
      port map(D => \ELINKS_STRT_ADDR_T[4]_net_1\, CLK => 
        CLK60MHZ, CLR => P_USB_MASTER_EN_c_17, E => 
        \REG_STATE_d[30]\, Q => \ELINKS_STRT_ADDR[4]_net_1\);
    
    \SM_BANK_SEL_RNI6GK1[16]\ : OR2
      port map(A => \SM_BANK_SEL[16]_net_1\, B => 
        \SM_BANK_SEL[21]_net_1\, Y => un1_SM_BANK_SEL_4);
    
    \WR_USB_ADBUS_RNO_9[0]\ : AO1
      port map(A => \ELINK_DOUTA_0[0]\, B => un1_SM_BANK_SEL_31, 
        C => \ELINK_DOUTA_16_m[0]\, Y => 
        \N_WR_USB_ADBUS_0_iv_14[0]\);
    
    \REG_STATE_0_RNIC10H4[0]\ : AO1
      port map(A => N_1744_i, B => N_1907, C => N_675_0, Y => 
        un1_REG_STATE_22);
    
    \WR_USB_ADBUS_RNO_19[5]\ : OR3A
      port map(A => N_1569, B => \ELINKS_STRT_ADDR_m[5]\, C => 
        \CHKSUM_m[5]\, Y => \N_WR_USB_ADBUS_0_iv_4[5]\);
    
    \WR_USB_ADBUS[6]\ : DFN1E0C0
      port map(D => \N_WR_USB_ADBUS[6]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_15, E => un1_REG_STATE_26, Q => 
        \WR_USB_ADBUS[6]_net_1\);
    
    \REG_STATE_ns_i_i_o2_6_1_RNO[0]\ : OA1B
      port map(A => N_449, B => N_450, C => 
        \REG_STATE_0[5]_net_1\, Y => N_487);
    
    \RD_XFER_TYPE[0]\ : DFN1C0
      port map(D => \RD_XFER_TYPE_RNO[0]_net_1\, CLK => CLK60MHZ, 
        CLR => P_USB_MASTER_EN_c, Q => \RD_XFER_TYPE[0]_net_1\);
    
    \ELINK_DINA_7[1]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[1]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_17, E => un1_SM_BANK_SEL_12, Q => 
        \ELINK_DINA_7[1]_net_1\);
    
    USB_RXF_B_0_RNI27AB1_0 : NOR3A
      port map(A => \REG_STATE_0[3]_net_1\, B => \USB_RXF_B_0\, C
         => \REG_STATE_0[4]_net_1\, Y => N_1907);
    
    \ELINK_ADDRA_12[2]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[2]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_2_0, E => un1_SM_BANK_SEL_7, Q => 
        \ELINK_ADDRA_12[2]_net_1\);
    
    \REG_ADDR_RNIN2HE[2]\ : OR2
      port map(A => \REG_ADDR[5]_net_1\, B => \REG_ADDR[2]_net_1\, 
        Y => REG_STATE_tr74_tz_tz_tz_2);
    
    \REG_ADDR_RNI9MA41[3]\ : OR3
      port map(A => \REG_ADDR[6]_net_1\, B => \REG_ADDR[3]_net_1\, 
        C => REG_STATE_tr74_tz_tz_tz_4, Y => 
        REG_STATE_tr74_tz_tz_tz_6);
    
    \SM_BANK_SEL_RNIL77M1[7]\ : OR3B
      port map(A => N_365, B => N_143, C => \N_ELINK_RWA_1[14]\, 
        Y => \N_ELINK_RWA_3[14]\);
    
    \REG_STATE_0_RNIF9MT1_1[4]\ : NOR3B
      port map(A => N_1359_2, B => N_1352_1, C => 
        \REG_STATE_0[4]_net_1\, Y => \REG_STATE_d[30]\);
    
    \ELINK_ADDRA_7[0]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[0]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_5, E => un1_SM_BANK_SEL_12, Q => 
        \ELINK_ADDRA_7[0]_net_1\);
    
    USB_RXF_B_RNIP2C35 : NOR3A
      port map(A => N_1351_i_i_a5_2, B => N_282, C => N_285, Y
         => N_358);
    
    U100_PATT_ELINK_BLK : DPRT_512X9_SRAM_0
      port map(ELINK_RWA_0 => \ELINK_RWA[0]_net_1\, 
        ELK_RX_SER_WORD_0(7) => ELK_RX_SER_WORD_0(7), 
        ELK_RX_SER_WORD_0(6) => ELK_RX_SER_WORD_0(6), 
        ELK_RX_SER_WORD_0(5) => ELK_RX_SER_WORD_0(5), 
        ELK_RX_SER_WORD_0(4) => ELK_RX_SER_WORD_0(4), 
        ELK_RX_SER_WORD_0(3) => ELK_RX_SER_WORD_0(3), 
        ELK_RX_SER_WORD_0(2) => ELK_RX_SER_WORD_0(2), 
        ELK_RX_SER_WORD_0(1) => ELK_RX_SER_WORD_0(1), 
        ELK_RX_SER_WORD_0(0) => ELK_RX_SER_WORD_0(0), 
        ELINK_DINA_0(7) => \ELINK_DINA_0[7]_net_1\, 
        ELINK_DINA_0(6) => \ELINK_DINA_0[6]_net_1\, 
        ELINK_DINA_0(5) => \ELINK_DINA_0[5]_net_1\, 
        ELINK_DINA_0(4) => \ELINK_DINA_0[4]_net_1\, 
        ELINK_DINA_0(3) => \ELINK_DINA_0[3]_net_1\, 
        ELINK_DINA_0(2) => \ELINK_DINA_0[2]_net_1\, 
        ELINK_DINA_0(1) => \ELINK_DINA_0[1]_net_1\, 
        ELINK_DINA_0(0) => \ELINK_DINA_0[0]_net_1\, ELINK_BLKA_0
         => \ELINK_BLKA[0]_net_1\, ELKS_ADDRB(7) => ELKS_ADDRB(7), 
        ELKS_ADDRB(6) => ELKS_ADDRB(6), ELKS_ADDRB(5) => 
        ELKS_ADDRB(5), ELKS_ADDRB(4) => ELKS_ADDRB(4), 
        ELKS_ADDRB(3) => ELKS_ADDRB(3), ELKS_ADDRB(2) => 
        ELKS_ADDRB(2), ELKS_ADDRB(1) => ELKS_ADDRB(1), 
        ELKS_ADDRB(0) => ELKS_ADDRB(0), ELINK_ADDRA_0(7) => 
        \ELINK_ADDRA_0[7]_net_1\, ELINK_ADDRA_0(6) => 
        \ELINK_ADDRA_0[6]_net_1\, ELINK_ADDRA_0(5) => 
        \ELINK_ADDRA_0[5]_net_1\, ELINK_ADDRA_0(4) => 
        \ELINK_ADDRA_0[4]_net_1\, ELINK_ADDRA_0(3) => 
        \ELINK_ADDRA_0[3]_net_1\, ELINK_ADDRA_0(2) => 
        \ELINK_ADDRA_0[2]_net_1\, ELINK_ADDRA_0(1) => 
        \ELINK_ADDRA_0[1]_net_1\, ELINK_ADDRA_0(0) => 
        \ELINK_ADDRA_0[0]_net_1\, PATT_ELK_DAT_0(7) => 
        PATT_ELK_DAT_0(7), PATT_ELK_DAT_0(6) => PATT_ELK_DAT_0(6), 
        PATT_ELK_DAT_0(5) => PATT_ELK_DAT_0(5), PATT_ELK_DAT_0(4)
         => PATT_ELK_DAT_0(4), PATT_ELK_DAT_0(3) => 
        PATT_ELK_DAT_0(3), PATT_ELK_DAT_0(2) => PATT_ELK_DAT_0(2), 
        PATT_ELK_DAT_0(1) => PATT_ELK_DAT_0(1), PATT_ELK_DAT_0(0)
         => PATT_ELK_DAT_0(0), ELINK_DOUTA_0(7) => 
        \ELINK_DOUTA_0[7]\, ELINK_DOUTA_0(6) => 
        \ELINK_DOUTA_0[6]\, ELINK_DOUTA_0(5) => 
        \ELINK_DOUTA_0[5]\, ELINK_DOUTA_0(4) => 
        \ELINK_DOUTA_0[4]\, ELINK_DOUTA_0(3) => 
        \ELINK_DOUTA_0[3]\, ELINK_DOUTA_0(2) => 
        \ELINK_DOUTA_0[2]\, ELINK_DOUTA_0(1) => 
        \ELINK_DOUTA_0[1]\, ELINK_DOUTA_0(0) => 
        \ELINK_DOUTA_0[0]\, ELKS_RWB => ELKS_RWB, 
        P_USB_MASTER_EN_c_0 => P_USB_MASTER_EN_c_0, CLK_40M_GL
         => CLK_40M_GL, CLK60MHZ => CLK60MHZ, ELKS_RAM_BLKB_EN
         => ELKS_RAM_BLKB_EN);
    
    \REG_STATE_RNIJVGL2[4]\ : OR2
      port map(A => N_2537_1, B => N_1784, Y => N_350);
    
    \ELINK_RWA_RNO_0[7]\ : OA1B
      port map(A => N_616_16, B => \N_ELINK_RWA_3[7]\, C => 
        \ELINK_RWA[7]_net_1\, Y => \ELINK_RWA_i_m[7]\);
    
    \REG_STATE_0_RNIE3U12[5]\ : AO1C
      port map(A => \REG_STATE_0[2]_net_1\, B => N_2515, C => 
        \REG_STATE_0[5]_net_1\, Y => \REG_STATE_ns_i_tz_0[5]\);
    
    \ELINK_DINA_18[6]\ : DFN1E0C0
      port map(D => \N_TFC_DINA[6]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_21, E => N_198, Q => 
        \ELINK_DINA_18[6]_net_1\);
    
    \ELINK_DINA_11[5]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[5]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_11, E => un1_SM_BANK_SEL_16, Q => 
        \ELINK_DINA_11[5]_net_1\);
    
    \WR_USB_ADBUS_RNO_17[5]\ : AO1A
      port map(A => N_1497, B => \TFC_STRT_ADDR[5]_net_1\, C => 
        \ELINKS_STOP_ADDR_m[5]\, Y => \N_WR_USB_ADBUS_0_iv_3[5]\);
    
    \RD_XFER_TYPE_RNIVRMR[4]\ : OR2
      port map(A => \RD_XFER_TYPE[4]_net_1\, B => 
        \RD_XFER_TYPE[5]_net_1\, Y => N_1367_i_i_o2_0_2);
    
    \ELINK_BLKA_RNO_0[0]\ : OA1B
      port map(A => N_616_16, B => \N_ELINK_RWA_3[0]\, C => 
        \ELINK_BLKA[0]_net_1\, Y => \ELINK_BLKA_i_m[0]\);
    
    \SM_BANK_SEL_RNO[19]\ : NOR3B
      port map(A => N_1882, B => N_1902, C => N_1700, Y => N_1848);
    
    \OP_MODE_T[7]\ : DFN1E1C0
      port map(D => \RD_USB_ADBUS[7]_net_1\, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_17, E => N_OP_MODE_T_0_sqmuxa, Q
         => \OP_MODE_T[7]_net_1\);
    
    \ELINK_ADDRA_0[0]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[0]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_18, E => un1_SM_BANK_SEL_6, Q => 
        \ELINK_ADDRA_0[0]_net_1\);
    
    \WR_USB_ADBUS_RNO_14[2]\ : NOR2B
      port map(A => \ELINK_DOUTA_5[2]\, B => un1_SM_BANK_SEL_35, 
        Y => \ELINK_DOUTA_5_m[2]\);
    
    \ELINK_BLKA_RNO[1]\ : AOI1
      port map(A => \SM_BANK_SEL[18]_net_1\, B => X_BLKA_i, C => 
        N_167, Y => \N_ELINK_BLKA_0_iv[1]\);
    
    \ELINK_DINA_13[2]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[2]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_14, E => un1_SM_BANK_SEL_2, Q => 
        \ELINK_DINA_13[2]_net_1\);
    
    \ELINK_ADDRA_0[1]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[1]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_18, E => un1_SM_BANK_SEL_6, Q => 
        \ELINK_ADDRA_0[1]_net_1\);
    
    \ELINK_BLKA_RNO[12]\ : AOI1
      port map(A => \SM_BANK_SEL[7]_net_1\, B => X_BLKA_i, C => 
        \ELINK_BLKA_i_m[12]\, Y => \N_ELINK_BLKA_0_iv[12]\);
    
    \WR_USB_ADBUS_RNO_19[2]\ : NOR2B
      port map(A => \ELINK_DOUTA_3[2]\, B => un1_SM_BANK_SEL_43, 
        Y => \ELINK_DOUTA_3_m[2]\);
    
    USB_RD_BI_RNO_8 : NOR3A
      port map(A => \REG_STATE_0[0]_net_1\, B => 
        \REG_STATE_0[2]_net_1\, C => \REG_STATE_0[3]_net_1\, Y
         => N_1868);
    
    \ELINKS_STOP_ADDR[4]\ : DFN1E1C0
      port map(D => \ELINKS_STOP_ADDR_T[4]_net_1\, CLK => 
        CLK60MHZ, CLR => P_USB_MASTER_EN_c_14, E => 
        \REG_STATE_d[30]\, Q => \ELINKS_STOP_ADDR[4]_net_1\);
    
    \WR_USB_ADBUS_RNO_30[1]\ : NOR3B
      port map(A => N_1352_1, B => \OP_MODE[1]_net_1\, C => 
        REG_STATE_s20_i_0, Y => \OP_MODE_m[1]\);
    
    \WR_USB_ADBUS_RNO_2[2]\ : OR3
      port map(A => \N_WR_USB_ADBUS_0_iv_18[2]\, B => 
        \N_WR_USB_ADBUS_0_iv_17[2]\, C => 
        \N_WR_USB_ADBUS_0_iv_24[2]\, Y => 
        \N_WR_USB_ADBUS_0_iv_26[2]\);
    
    \WR_USB_ADBUS_RNO_10[5]\ : OR2
      port map(A => \ELINK_DOUTA_6_m[5]\, B => 
        \ELINK_DOUTA_8_m[5]\, Y => \N_WR_USB_ADBUS_0_iv_13[5]\);
    
    \ELINK_DINA_12[1]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[1]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_12, E => un1_SM_BANK_SEL_7, Q => 
        \ELINK_DINA_12[1]_net_1\);
    
    \ELINK_DINA_1[3]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[3]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_7, E => un1_SM_BANK_SEL_19, Q => 
        \ELINK_DINA_1[3]_net_1\);
    
    \WR_USB_ADBUS_RNO_18[3]\ : OR3
      port map(A => \OP_MODE_m[3]\, B => \TFC_STOP_ADDR_m[3]\, C
         => \WR_XFER_TYPE_m[3]\, Y => \N_WR_USB_ADBUS_0_iv_2[3]\);
    
    \SM_BANK_SEL_RNIM873[18]\ : OR3
      port map(A => \SM_BANK_SEL[17]_net_1\, B => 
        \SM_BANK_SEL[18]_net_1\, C => N_616_2, Y => 
        \N_ELINK_RWA_1[0]\);
    
    \REG_ADDR_RNIMD2T[6]\ : NOR3C
      port map(A => \REG_ADDR[7]_net_1\, B => \REG_ADDR[6]_net_1\, 
        C => N_491, Y => REG_STATE_tr49_3);
    
    \ELINK_RWA_RNO_0[1]\ : OA1B
      port map(A => N_616_16, B => \N_ELINK_RWA_3[1]\, C => 
        \ELINK_RWA[1]_net_1\, Y => N_185);
    
    \RD_USB_ADBUS_RNIJQ0T[7]\ : NOR2B
      port map(A => \RD_USB_ADBUS[7]_net_1\, B => N_1352_5, Y => 
        N_USB_OE_BI_iv_0_i_a2_0_1);
    
    \ELINK_RWA[8]\ : DFN1E0P0
      port map(D => \N_ELINK_RWA_0_iv[8]\, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_6, E => \SM_BANK_SEL_0[20]_net_1\, 
        Q => \ELINK_RWA[8]_net_1\);
    
    \ELINK_RWA[5]\ : DFN1E0P0
      port map(D => \N_ELINK_RWA_0_iv[5]\, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_6, E => \SM_BANK_SEL_0[20]_net_1\, 
        Q => \ELINK_RWA[5]_net_1\);
    
    \ELINK_DINA_19[3]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[3]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_1, E => un1_SM_BANK_SEL_11, Q => 
        \ELINK_DINA_19[3]_net_1\);
    
    \SM_BANK_SEL_RNI399C[1]\ : NOR2
      port map(A => N_624_15, B => \SM_BANK_SEL[1]_net_1\, Y => 
        N_464);
    
    \ELINKS_STRT_ADDR_T[2]\ : DFN1E1C0
      port map(D => \RD_USB_ADBUS[2]_net_1\, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_21, E => 
        N_ELINKS_STRT_ADDR_T_0_sqmuxa, Q => 
        \ELINKS_STRT_ADDR_T[2]_net_1\);
    
    \REG_STATE_RNI04LF1[3]\ : NOR2A
      port map(A => N_1359_1, B => N_292, Y => N_418);
    
    \REG_STATE_ns_i_i_o2_6_1[0]\ : OR2
      port map(A => N_487, B => \REG_STATE_ns_i_i_o2_6_0[0]\, Y
         => \REG_STATE_ns_i_i_o2_6_1[0]_net_1\);
    
    \ELINK_RWA_RNO_0[4]\ : OA1B
      port map(A => N_616_16, B => \N_ELINK_RWA_1[4]\, C => 
        \ELINK_RWA[4]_net_1\, Y => \ELINK_RWA_i_m[4]\);
    
    \ELINK_DINA_14[0]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[0]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_16, E => un1_SM_BANK_SEL_1, Q => 
        \ELINK_DINA_14[0]_net_1\);
    
    \REG_STATE_RNI61O31[3]\ : OR2A
      port map(A => \REG_STATE[3]_net_1\, B => N_252, Y => N_255);
    
    \REG_STATE_RNI2KQN[1]\ : NOR2B
      port map(A => \REG_STATE[1]_net_1\, B => 
        \REG_STATE[5]_net_1\, Y => N_2600);
    
    \ELINK_BLKA[6]\ : DFN1E0P0
      port map(D => \N_ELINK_BLKA_0_iv[6]\, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_19, E => \SM_BANK_SEL[20]_net_1\, Q
         => \ELINK_BLKA[6]_net_1\);
    
    \WR_XFER_TYPE_RNO[2]\ : NOR3
      port map(A => N_1824, B => N_1823, C => N_1822, Y => 
        \WR_XFER_TYPE_RNO[2]_net_1\);
    
    \WR_USB_ADBUS_RNO_15[1]\ : NOR2B
      port map(A => \ELINK_DOUTA_18[1]\, B => un1_SM_BANK_SEL_25, 
        Y => \ELINK_DOUTA_18_m[1]\);
    
    USB_OE_BI_RNO_0 : AO1D
      port map(A => N_1879, B => N_1756, C => N_1862, Y => N_1669);
    
    ELK_N_ACTIVE_RNIP1UMP : NOR3A
      port map(A => \REG_STATE_ns_i_a2_0[3]\, B => N_359, C => 
        N_357, Y => N_2592);
    
    \WR_USB_ADBUS_RNO_7[3]\ : NOR2B
      port map(A => \ELINK_DOUTA_14[3]\, B => un1_SM_BANK_SEL_23, 
        Y => \ELINK_DOUTA_14_m[3]\);
    
    \WR_USB_ADBUS_RNO_21[0]\ : NOR2B
      port map(A => \ELINK_DOUTA_3[0]\, B => un1_SM_BANK_SEL_43, 
        Y => \ELINK_DOUTA_3_m[0]\);
    
    \REG_STATE_0[0]\ : DFN1C0
      port map(D => \REG_STATE_ns_i_i_a2_0_RNIN0TJ41[0]_net_1\, 
        CLK => CLK60MHZ, CLR => P_USB_MASTER_EN_c_22_0, Q => 
        \REG_STATE_0[0]_net_1\);
    
    ELK_N_ACTIVE : DFN1C0
      port map(D => \ELK_N_ACTIVE_RNO\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_22, Q => \ELK_N_ACTIVE\);
    
    \RD_USB_ADBUS[6]\ : DFN1C0
      port map(D => \N_RD_USB_ADBUS[6]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_22_0, Q => \RD_USB_ADBUS[6]_net_1\);
    
    \RD_USB_ADBUS_RNI38BJ_1[4]\ : NOR2
      port map(A => \RD_USB_ADBUS[4]_net_1\, B => 
        \RD_USB_ADBUS[5]_net_1\, Y => N_1351_i_i_a5_0);
    
    \ELINKS_STOP_ADDR_T[4]\ : DFN1E1C0
      port map(D => \RD_USB_ADBUS[4]_net_1\, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_7, E => 
        N_ELINKS_STOP_ADDR_T_0_sqmuxa, Q => 
        \ELINKS_STOP_ADDR_T[4]_net_1\);
    
    \WR_USB_ADBUS_RNO_33[7]\ : NOR2B
      port map(A => \ELINK_DOUTA_13[7]\, B => un1_SM_BANK_SEL_29, 
        Y => \ELINK_DOUTA_13_m[7]\);
    
    \REG_STATE_ns_i_i_o2_1_RNO_6[0]\ : NOR2A
      port map(A => \REG_STATE[2]_net_1\, B => N_287, Y => N_437);
    
    \REG_ADDR[4]\ : DFN1E1C0
      port map(D => REG_ADDR_n4, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_10, E => REG_ADDRe, Q => 
        \REG_ADDR[4]_net_1\);
    
    \WR_USB_ADBUS_RNO_14[3]\ : NOR2B
      port map(A => \ELINK_DOUTA_3[3]\, B => un1_SM_BANK_SEL_43, 
        Y => \ELINK_DOUTA_3_m[3]\);
    
    \ELINK_ADDRA_18[7]\ : DFN1E0C0
      port map(D => \N_TFC_ADDRA[7]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_12, E => N_198, Q => 
        \ELINK_ADDRA_18[7]_net_1\);
    
    \WR_USB_ADBUS_RNO_28[1]\ : NOR2B
      port map(A => \ELINK_DOUTA_5[1]\, B => un1_SM_BANK_SEL_35, 
        Y => \ELINK_DOUTA_5_m[1]\);
    
    \RD_USB_ADBUS_RNIOCIK2[3]\ : NOR2A
      port map(A => \RD_USB_ADBUS[3]_net_1\, B => N_206, Y => 
        \N_TFC_DINA[3]\);
    
    \OP_MODE[0]\ : DFN1E1C0
      port map(D => \OP_MODE_T[0]_net_1\, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_15, E => \REG_STATE_d[30]\, Q => 
        \OP_MODE[0]_net_1\);
    
    \ELINK_RWA[14]\ : DFN1E0P0
      port map(D => \N_ELINK_RWA_0_iv[14]\, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_12, E => \SM_BANK_SEL_0[20]_net_1\, 
        Q => \ELINK_RWA[14]_net_1\);
    
    \SM_BANK_SEL_RNIF5P72[3]\ : NOR3A
      port map(A => \SM_BANK_SEL[3]_net_1\, B => N_312, C => 
        N_1566_i_i_0, Y => un1_SM_BANK_SEL_39);
    
    \N_TFC_ADDRA_0_o2[7]\ : OR2
      port map(A => N_429, B => \N_TFC_ADDRA_0_o2_0[7]\, Y => 
        N_261);
    
    \ELINK_DINA_13[4]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[4]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_14, E => un1_SM_BANK_SEL_2, Q => 
        \ELINK_DINA_13[4]_net_1\);
    
    \WR_USB_ADBUS_RNO_3[2]\ : NOR2B
      port map(A => \ELINK_DOUTA_17[2]\, B => un1_SM_BANK_SEL_40, 
        Y => \ELINK_DOUTA_17_m[2]\);
    
    USB_RXF_B_0_RNIKK3L1 : AO1A
      port map(A => \REG_STATE_0[4]_net_1\, B => \USB_RXF_B_0\, C
         => N_2600, Y => \REG_STATE_ns_i_1_tz_0[3]\);
    
    \SM_BANK_SEL_RNIAECN[5]\ : NOR3A
      port map(A => N_462, B => \SM_BANK_SEL[6]_net_1\, C => 
        \SM_BANK_SEL[5]_net_1\, Y => N_477);
    
    \WR_USB_ADBUS_RNO_20[3]\ : NOR2A
      port map(A => \TFC_DOUTA[3]\, B => N_243, Y => 
        \TFC_DOUTA_m[3]\);
    
    \REG_STATE_ns_i_i_o2_6_RNISP5I5[0]\ : OA1
      port map(A => N_244_1, B => N_504, C => 
        \REG_STATE_ns_i_i_a5_1_3[0]\, Y => N_388);
    
    \WR_USB_ADBUS_RNO_30[4]\ : NOR2B
      port map(A => \ELINK_DOUTA_18[4]\, B => un1_SM_BANK_SEL_25, 
        Y => \ELINK_DOUTA_18_m[4]\);
    
    \WR_USB_ADBUS_RNO_2[7]\ : OR3
      port map(A => \N_WR_USB_ADBUS_0_iv_14[7]\, B => 
        \N_WR_USB_ADBUS_0_iv_13[7]\, C => 
        \N_WR_USB_ADBUS_0_iv_22[7]\, Y => 
        \N_WR_USB_ADBUS_0_iv_25[7]\);
    
    \REG_STATE_RNIVPN31[0]\ : NOR2A
      port map(A => N_268, B => \REG_STATE[0]_net_1\, Y => N_379);
    
    \WR_USB_ADBUS_RNO_19[1]\ : OR3A
      port map(A => N_1569, B => \ELINKS_STRT_ADDR_m[1]\, C => 
        \CHKSUM_m[1]\, Y => \N_WR_USB_ADBUS_0_iv_4[1]\);
    
    \TFC_STRT_ADDR_T[1]\ : DFN1E1C0
      port map(D => \RD_USB_ADBUS[1]_net_1\, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_4, E => N_TFC_STRT_ADDR_T_0_sqmuxa, 
        Q => \TFC_STRT_ADDR_T[1]_net_1\);
    
    \OP_MODE[1]\ : DFN1E1C0
      port map(D => \OP_MODE_T[1]_net_1\, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_15, E => \REG_STATE_d[30]\, Q => 
        \OP_MODE[1]_net_1\);
    
    \WR_XFER_TYPE[5]\ : DFN1C0
      port map(D => \WR_XFER_TYPE_RNO[5]_net_1\, CLK => CLK60MHZ, 
        CLR => P_USB_MASTER_EN_c, Q => \WR_XFER_TYPE[5]_net_1\);
    
    \WR_USB_ADBUS_RNO_30[0]\ : NOR2B
      port map(A => \ELINK_DOUTA_18[0]\, B => un1_SM_BANK_SEL_25, 
        Y => \ELINK_DOUTA_18_m[0]\);
    
    \REG_ADDR_RNI2FA41[4]\ : NOR2B
      port map(A => REG_ADDR_c3, B => \REG_ADDR[4]_net_1\, Y => 
        REG_ADDR_c4);
    
    \CHKSUM[5]\ : DFN1E1C0
      port map(D => N_230, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_3, E => un1_REG_STATE_22, Q => 
        \CHKSUM[5]_net_1\);
    
    \RD_USB_ADBUS_RNIIP0T[6]\ : NOR2B
      port map(A => \RD_USB_ADBUS[6]_net_1\, B => N_1359_6, Y => 
        N_1367_i_i_a2_0);
    
    \CHKSUM_RNO[0]\ : NOR2A
      port map(A => \RD_USB_ADBUS[0]_net_1\, B => N_675, Y => 
        N_1593);
    
    \SM_BANK_SEL_RNIBNN91[10]\ : OR3B
      port map(A => N_461, B => N_477, C => \N_ELINK_RWA_16_0[0]\, 
        Y => N_616_16);
    
    \ELINKS_STRT_ADDR_T[5]\ : DFN1E1C0
      port map(D => \RD_USB_ADBUS[5]_net_1\, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_21, E => 
        N_ELINKS_STRT_ADDR_T_0_sqmuxa, Q => 
        \ELINKS_STRT_ADDR_T[5]_net_1\);
    
    \SM_BANK_SEL_RNO[15]\ : NOR3C
      port map(A => N_1882, B => N_1359_6, C => N_1902, Y => 
        N_1843);
    
    \ELINK_DINA_16[6]\ : DFN1E0C0
      port map(D => \N_TFC_DINA[6]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_18, E => N_200, Q => 
        \ELINK_DINA_16[6]_net_1\);
    
    \ELINK_DINA_3[0]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[0]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_11, E => un1_SM_BANK_SEL_4, Q => 
        \ELINK_DINA_3[0]_net_1\);
    
    \ELINK_BLKA[4]\ : DFN1E0P0
      port map(D => \N_ELINK_BLKA_0_iv[4]\, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_19, E => \SM_BANK_SEL[20]_net_1\, Q
         => \ELINK_BLKA[4]_net_1\);
    
    \ELINKS_STRT_ADDR_T[1]\ : DFN1E1C0
      port map(D => \RD_USB_ADBUS[1]_net_1\, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_21, E => 
        N_ELINKS_STRT_ADDR_T_0_sqmuxa, Q => 
        \ELINKS_STRT_ADDR_T[1]_net_1\);
    
    \WR_XFER_TYPE_RNO[0]\ : NOR3
      port map(A => N_1816, B => N_1818, C => N_1817, Y => 
        \WR_XFER_TYPE_RNO[0]_net_1\);
    
    \REG_STATE_RNI904KE[2]\ : AO1
      port map(A => \REG_STATE_ns_i_i_a5_1_3[0]\, B => N_504, C
         => N_384, Y => \REG_STATE_ns_i_i_0[2]\);
    
    \ELINK_ADDRA_7[7]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[7]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_6, E => un1_SM_BANK_SEL_12, Q => 
        \ELINK_ADDRA_7[7]_net_1\);
    
    USB_RD_BI_RNO_6 : NOR2B
      port map(A => un1_REG_STATE_40_i_a2_0, B => N_1877_1, Y => 
        N_1877);
    
    \RD_USB_ADBUS[3]\ : DFN1C0
      port map(D => \N_RD_USB_ADBUS[3]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_22, Q => \RD_USB_ADBUS[3]_net_1\);
    
    \SM_BANK_SEL_RNI5FK1[15]\ : OR2
      port map(A => \SM_BANK_SEL[15]_net_1\, B => 
        \SM_BANK_SEL[21]_net_1\, Y => un1_SM_BANK_SEL_8);
    
    \WR_USB_ADBUS_RNO_17[6]\ : NOR2B
      port map(A => \ELINK_DOUTA_6[6]\, B => un1_SM_BANK_SEL_30, 
        Y => \ELINK_DOUTA_6_m[6]\);
    
    \ELINK_DINA_15[7]\ : DFN1E0C0
      port map(D => \N_TFC_DINA[7]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_17, E => N_199, Q => 
        \ELINK_DINA_15[7]_net_1\);
    
    \ELINKS_STOP_ADDR_T[1]\ : DFN1E1C0
      port map(D => \RD_USB_ADBUS[1]_net_1\, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_7, E => 
        N_ELINKS_STOP_ADDR_T_0_sqmuxa, Q => 
        \ELINKS_STOP_ADDR_T[1]_net_1\);
    
    \ELINK_ADDRA_9[6]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[6]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_10, E => un1_SM_BANK_SEL_9, Q => 
        \ELINK_ADDRA_9[6]_net_1\);
    
    \WR_USB_ADBUS_RNO_12[1]\ : NOR2B
      port map(A => \ELINK_DOUTA_2[1]\, B => un1_SM_BANK_SEL_32, 
        Y => \ELINK_DOUTA_2_m[1]\);
    
    \TFC_STOP_ADDR_T[3]\ : DFN1E1C0
      port map(D => \RD_USB_ADBUS[3]_net_1\, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_15, E => N_TFC_STOP_ADDR_T_0_sqmuxa, 
        Q => \TFC_STOP_ADDR_T[3]_net_1\);
    
    \ELINK_RWA[16]\ : DFN1E0P0
      port map(D => \N_ELINK_RWA_0_iv[16]\, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_12, E => \SM_BANK_SEL_0[20]_net_1\, 
        Q => \ELINK_RWA[16]_net_1\);
    
    \WR_USB_ADBUS_RNO_13[0]\ : NOR2B
      port map(A => \ELINK_DOUTA_9[0]\, B => un1_SM_BANK_SEL_42, 
        Y => \ELINK_DOUTA_9_m[0]\);
    
    \N_TFC_ADDRA_0_o2_2[7]\ : OR2
      port map(A => \SM_BANK_SEL[20]_net_1\, B => \ELK_N_ACTIVE\, 
        Y => N_251);
    
    un1_N_WR_USB_ADBUS_0_sqmuxa_i : OR2
      port map(A => N_78, B => \un1_N_WR_USB_ADBUS_0_sqmuxa_i_0\, 
        Y => N_243);
    
    \REG_STATE[5]\ : DFN1C0
      port map(D => \USB_TXE_B_RNIV2O4Q\, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_22_0, Q => \REG_STATE[5]_net_1\);
    
    \ELINK_BLKA_RNO_0[1]\ : OA1B
      port map(A => N_616_16, B => \N_ELINK_RWA_3[1]\, C => 
        \ELINK_BLKA[1]_net_1\, Y => N_167);
    
    \ELINK_ADDRA_0[7]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[7]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_19, E => un1_SM_BANK_SEL_6, Q => 
        \ELINK_ADDRA_0[7]_net_1\);
    
    \WR_USB_ADBUS_RNO_12[6]\ : NOR2B
      port map(A => \ELINK_DOUTA_18[6]\, B => un1_SM_BANK_SEL_25, 
        Y => \ELINK_DOUTA_18_m[6]\);
    
    \SM_BANK_SEL_RNO[3]\ : NOR3B
      port map(A => un1_N_ELK_N_ACTIVE_0_sqmuxa_15_0_a2_0_0, B
         => N_1902, C => N_1697, Y => N_1849);
    
    \RD_USB_ADBUS_RNIVD4K6[4]\ : AO1A
      port map(A => N_282, B => \REG_STATE_ns_i_i_a5_0_1_0[2]\, C
         => \REG_STATE_ns_i_i_a5_1[2]\, Y => N_1294_tz);
    
    \REG_STATE_RNI4KDN1[2]\ : NOR2A
      port map(A => N_1862_1, B => N_1700, Y => 
        un1_REG_STATE_39_i_a2_0);
    
    \REG_STATE_ns_i_8_tz_1[4]\ : OR2
      port map(A => \REG_STATE_ns_i_a4_1_0[4]_net_1\, B => 
        \REG_STATE_ns_i_8_tz_0[4]_net_1\, Y => 
        \REG_STATE_ns_i_8_tz_1[4]_net_1\);
    
    \REG_STATE_0_RNI3HUOT[5]\ : OA1
      port map(A => \REG_STATE_ns_i_a4_0[1]\, B => N_1282_tz, C
         => N_2587, Y => \REG_STATE_ns_i_4[1]\);
    
    \RD_XFER_TYPE_RNO_0[7]\ : NOR2A
      port map(A => \RD_USB_ADBUS[7]_net_1\, B => N_1694, Y => 
        N_1808);
    
    \ELINKS_STOP_ADDR[5]\ : DFN1E1C0
      port map(D => \ELINKS_STOP_ADDR_T[5]_net_1\, CLK => 
        CLK60MHZ, CLR => P_USB_MASTER_EN_c_14, E => 
        \REG_STATE_d[30]\, Q => \ELINKS_STOP_ADDR[5]_net_1\);
    
    \REG_STATE[0]\ : DFN1C0
      port map(D => \REG_STATE_ns_i_i_a2_0_RNIN0TJ41[0]_net_1\, 
        CLK => CLK60MHZ, CLR => P_USB_MASTER_EN_c_22_0, Q => 
        \REG_STATE[0]_net_1\);
    
    \ELINK_DINA_10[1]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[1]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_9, E => un1_SM_BANK_SEL_20, Q => 
        \ELINK_DINA_10[1]_net_1\);
    
    \WR_XFER_TYPE_RNO_0[3]\ : NOR2
      port map(A => N_1716, B => \RD_USB_ADBUS[3]_net_1\, Y => 
        N_1826);
    
    \ELINK_DINA_4[2]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[2]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_13, E => un1_SM_BANK_SEL_8, Q => 
        \ELINK_DINA_4[2]_net_1\);
    
    \TFC_ADDRA[6]\ : DFN1E0C0
      port map(D => \N_TFC_ADDRA[6]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_10, E => N_142, Q => 
        \TFC_ADDRA[6]_net_1\);
    
    \REG_STATE_ns_i_i_o2_6_1_RNO_1[0]\ : NOR2B
      port map(A => N_1352_2, B => N_414_1, Y => N_449);
    
    \ELINK_ADDRA_16[0]\ : DFN1E0C0
      port map(D => \N_TFC_ADDRA[0]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_8, E => N_200, Q => 
        \ELINK_ADDRA_16[0]_net_1\);
    
    \WR_USB_ADBUS_RNO_14[7]\ : NOR2B
      port map(A => \ELINK_DOUTA_3[7]\, B => un1_SM_BANK_SEL_43, 
        Y => \ELINK_DOUTA_3_m[7]\);
    
    \ELINK_RWA_RNO_0[15]\ : AOI1
      port map(A => \N_ELINK_RWA_0_iv_0_o2_i_a5_0[15]\, B => 
        N_503, C => \ELINK_RWA[15]_net_1\, Y => N_175);
    
    \WR_USB_ADBUS_RNO_34[1]\ : NOR2B
      port map(A => \CHKSUM[1]_net_1\, B => un1_REG_STATE_4, Y
         => \CHKSUM_m[1]\);
    
    \WR_USB_ADBUS_RNO_20[6]\ : AO1A
      port map(A => N_1497, B => \TFC_STRT_ADDR[6]_net_1\, C => 
        \ELINKS_STOP_ADDR_m[6]\, Y => \N_WR_USB_ADBUS_0_iv_3[6]\);
    
    \RD_USB_ADBUS_RNIRCVLB[7]\ : AOI1B
      port map(A => REG_STATE_tr67_5, B => N_1404_8, C => 
        N_1387_i, Y => \REG_STATE_ns_i_a2_0[4]\);
    
    \WR_USB_ADBUS_RNO_15[0]\ : NOR2B
      port map(A => \ELINK_DOUTA_12[0]\, B => un1_SM_BANK_SEL_33, 
        Y => \ELINK_DOUTA_12_m[0]\);
    
    \RD_XFER_TYPE_RNO_0[0]\ : NOR2A
      port map(A => \RD_USB_ADBUS[0]_net_1\, B => N_1694, Y => 
        N_1794);
    
    ELK_N_ACTIVE_RNO_0 : OA1
      port map(A => \USB_RXF_B_0\, B => N_1694, C => 
        \ELK_N_ACTIVE\, Y => N_1873);
    
    \ELINK_DINA_7[5]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[5]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_17, E => un1_SM_BANK_SEL_12, Q => 
        \ELINK_DINA_7[5]_net_1\);
    
    \WR_USB_ADBUS_RNO_21[2]\ : AO1
      port map(A => \ELINK_DOUTA_8[2]\, B => un1_SM_BANK_SEL_38, 
        C => \ELINK_DOUTA_9_m[2]\, Y => 
        \N_WR_USB_ADBUS_0_iv_9[2]\);
    
    \ELINK_DINA_2[4]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[4]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_9, E => un1_SM_BANK_SEL_5, Q => 
        \ELINK_DINA_2[4]_net_1\);
    
    \ELINK_DINA_10[3]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[3]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_9, E => un1_SM_BANK_SEL_20, Q => 
        \ELINK_DINA_10[3]_net_1\);
    
    \CHKSUM_RNO[5]\ : NOR2A
      port map(A => \RD_USB_ADBUS[5]_net_1\, B => N_675, Y => 
        N_230);
    
    \WR_USB_ADBUS_RNO_16[5]\ : AO1
      port map(A => \ELINK_DOUTA_4[5]\, B => un1_SM_BANK_SEL_28, 
        C => \ELINK_DOUTA_5_m[5]\, Y => 
        \N_WR_USB_ADBUS_0_iv_12[5]\);
    
    \ELINK_DINA_1[0]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[0]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_7, E => un1_SM_BANK_SEL_19, Q => 
        \ELINK_DINA_1[0]_net_1\);
    
    \ELINK_DINA_9[0]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[0]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_19, E => un1_SM_BANK_SEL_9, Q => 
        \ELINK_DINA_9[0]_net_1\);
    
    \SM_BANK_SEL_RNO[4]\ : NOR3B
      port map(A => \RD_USB_ADBUS[2]_net_1\, B => N_1892, C => 
        N_290, Y => N_1832);
    
    \WR_USB_ADBUS[4]\ : DFN1E0C0
      port map(D => \N_WR_USB_ADBUS[4]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_15, E => un1_REG_STATE_26, Q => 
        \WR_USB_ADBUS[4]_net_1\);
    
    \ELINK_BLKA_RNO[6]\ : OA1C
      port map(A => N_622, B => \ELINK_BLKA[6]_net_1\, C => 
        X_BLKA_i_m_5, Y => \N_ELINK_BLKA_0_iv[6]\);
    
    \TFC_ADDRA[2]\ : DFN1E0C0
      port map(D => \N_TFC_ADDRA[2]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_9, E => N_142, Q => 
        \TFC_ADDRA[2]_net_1\);
    
    \OP_MODE[2]\ : DFN1E1C0
      port map(D => \OP_MODE_T[2]_net_1\, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_15, E => \REG_STATE_d[30]\, Q => 
        \OP_MODE[2]_net_1\);
    
    USB_TRIEN_B_RNO : AO1A
      port map(A => N_1749, B => N_1917, C => N_675_0, Y => 
        un1_REG_STATE_23);
    
    \TFC_STOP_ADDR_T[6]\ : DFN1E1C0
      port map(D => \RD_USB_ADBUS[6]_net_1\, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_15, E => N_TFC_STOP_ADDR_T_0_sqmuxa, 
        Q => \TFC_STOP_ADDR_T[6]_net_1\);
    
    \REG_ADDR_RNILMPL[8]\ : NOR3B
      port map(A => \REG_ADDR[2]_net_1\, B => \REG_ADDR[3]_net_1\, 
        C => \REG_ADDR[8]_net_1\, Y => REG_STATE_tr49_2);
    
    \RD_USB_ADBUS_RNIH2N32[4]\ : NOR3B
      port map(A => N_1351_i_i_a5_0, B => N_465, C => N_1700, Y
         => N_1351_i_i_a5_2);
    
    \RD_XFER_TYPE_RNINJMR_1[0]\ : NOR2A
      port map(A => \RD_XFER_TYPE[0]_net_1\, B => 
        \RD_XFER_TYPE[1]_net_1\, Y => N_1370_i_i_a5_0);
    
    \WR_USB_ADBUS_RNO_5[7]\ : OR3
      port map(A => \ELINK_DOUTA_3_m[7]\, B => 
        \ELINK_DOUTA_18_m[7]\, C => \N_WR_USB_ADBUS_0_iv_12[7]\, 
        Y => \N_WR_USB_ADBUS_0_iv_20[7]\);
    
    \ELINK_DINA_11[1]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[1]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_11, E => un1_SM_BANK_SEL_16, Q => 
        \ELINK_DINA_11[1]_net_1\);
    
    \REG_STATE[3]\ : DFN1C0
      port map(D => \REG_STATE_0_RNIGPV6T1[0]_net_1\, CLK => 
        CLK60MHZ, CLR => P_USB_MASTER_EN_c_22_0, Q => 
        \REG_STATE[3]_net_1\);
    
    \RD_XFER_TYPE_RNILOOSL[0]\ : NOR3A
      port map(A => \REG_STATE_ns_i_a2_0[1]\, B => N_359, C => 
        N_358, Y => N_2587);
    
    \WR_USB_ADBUS_RNO_33[2]\ : NOR2A
      port map(A => \ELINKS_STRT_ADDR[2]_net_1\, B => N_1499, Y
         => \ELINKS_STRT_ADDR_m[2]\);
    
    \WR_USB_ADBUS_RNO_6[0]\ : AO1
      port map(A => \ELINK_DOUTA_6[0]\, B => un1_SM_BANK_SEL_30, 
        C => \ELINK_DOUTA_7_m[0]\, Y => 
        \N_WR_USB_ADBUS_0_iv_8[0]\);
    
    \RD_USB_ADBUS_RNI5KNJ2[6]\ : OR2
      port map(A => N_1695, B => N_1694, Y => N_1697);
    
    \SM_BANK_SEL_RNIBKJ1[16]\ : OR2
      port map(A => \SM_BANK_SEL[16]_net_1\, B => 
        \SM_BANK_SEL[17]_net_1\, Y => \N_ELINK_BLKA_10_0[10]\);
    
    \TFC_STRT_ADDR_T[3]\ : DFN1E1C0
      port map(D => \RD_USB_ADBUS[3]_net_1\, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_4, E => N_TFC_STRT_ADDR_T_0_sqmuxa, 
        Q => \TFC_STRT_ADDR_T[3]_net_1\);
    
    \WR_XFER_TYPE_RNI0FP34_0[5]\ : NOR3B
      port map(A => REG_STATE_tr72_6_3, B => N_1404_7, C => N_252, 
        Y => REG_STATE_tr72_6_5);
    
    \TFC_STRT_ADDR_T[4]\ : DFN1E1C0
      port map(D => \RD_USB_ADBUS[4]_net_1\, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_4, E => N_TFC_STRT_ADDR_T_0_sqmuxa, 
        Q => \TFC_STRT_ADDR_T[4]_net_1\);
    
    \ELINK_RWA_RNO[2]\ : AOI1
      port map(A => \SM_BANK_SEL[17]_net_1\, B => un1_USB_RXF_B_m, 
        C => \ELINK_RWA_i_m[2]\, Y => \N_ELINK_RWA_0_iv[2]\);
    
    \ELINK_ADDRA_0[3]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[3]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_18, E => un1_SM_BANK_SEL_6, Q => 
        \ELINK_ADDRA_0[3]_net_1\);
    
    \REG_STATE_RNIU1LF1[3]\ : NOR2B
      port map(A => N_1359_2, B => N_1359_1, Y => N_1367_i_i_a2_3);
    
    \REG_ADDR_RNO[5]\ : XA1B
      port map(A => REG_ADDR_c4, B => \REG_ADDR[5]_net_1\, C => 
        N_675_0, Y => REG_ADDR_n5);
    
    \ELINK_RWA_RNO_0[19]\ : NOR2B
      port map(A => \SM_BANK_SEL[0]_net_1\, B => un1_USB_RXF_B_m, 
        Y => N_170);
    
    \ELINK_ADDRA_6[6]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[6]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_4, E => un1_SM_BANK_SEL_10, Q => 
        \ELINK_ADDRA_6[6]_net_1\);
    
    \WR_USB_ADBUS_RNO_28[6]\ : OR3
      port map(A => \N_WR_USB_ADBUS_0_iv_0[6]_net_1\, B => 
        \OP_MODE_m[6]\, C => \ELINKS_STRT_ADDR_m[6]\, Y => 
        \N_WR_USB_ADBUS_0_iv_2[6]\);
    
    \REG_STATE_RNI5G241[2]\ : NOR2A
      port map(A => \REG_STATE[2]_net_1\, B => N_1695, Y => 
        N_1862_1);
    
    \ELINK_RWA_RNO_0[17]\ : NOR2B
      port map(A => \SM_BANK_SEL[2]_net_1\, B => un1_USB_RXF_B_m, 
        Y => N_174);
    
    \ELINK_DINA_19[5]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[5]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_1, E => un1_SM_BANK_SEL_11, Q => 
        \ELINK_DINA_19[5]_net_1\);
    
    \ELINK_DINA_12[6]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[6]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_12, E => un1_SM_BANK_SEL_7, Q => 
        \ELINK_DINA_12[6]_net_1\);
    
    \ELINK_ADDRA_5[4]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[4]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_3, E => un1_SM_BANK_SEL_15, Q => 
        \ELINK_ADDRA_5[4]_net_1\);
    
    \WR_USB_ADBUS_RNO_17[1]\ : AO1A
      port map(A => N_1497, B => \TFC_STRT_ADDR[1]_net_1\, C => 
        \ELINKS_STOP_ADDR_m[1]\, Y => \N_WR_USB_ADBUS_0_iv_3[1]\);
    
    \OP_MODE_T[2]\ : DFN1E1C0
      port map(D => \RD_USB_ADBUS[2]_net_1\, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_17, E => N_OP_MODE_T_0_sqmuxa, Q
         => \OP_MODE_T[2]_net_1\);
    
    \RD_USB_ADBUS_RNIVNN03[4]\ : AO1
      port map(A => N_1903, B => N_1352_4, C => N_1698, Y => 
        N_1772);
    
    \WR_USB_ADBUS_RNO_22[2]\ : OR3
      port map(A => \ELINK_DOUTA_13_m[2]\, B => 
        \ELINK_DOUTA_12_m[2]\, C => \N_WR_USB_ADBUS_0_iv_12[2]\, 
        Y => \N_WR_USB_ADBUS_0_iv_20[2]\);
    
    \SM_BANK_SEL_RNI6O63[14]\ : OR3
      port map(A => \SM_BANK_SEL[13]_net_1\, B => 
        \SM_BANK_SEL[14]_net_1\, C => N_616_4, Y => N_616_11);
    
    \WR_USB_ADBUS_RNO_24[0]\ : NOR2B
      port map(A => \ELINK_DOUTA_17[0]\, B => un1_SM_BANK_SEL_40, 
        Y => \ELINK_DOUTA_17_m[0]\);
    
    \WR_USB_ADBUS_RNO_19[4]\ : AO1
      port map(A => \CHKSUM[4]_net_1\, B => un1_REG_STATE_4, C
         => \N_WR_USB_ADBUS_0_iv_3[4]\, Y => 
        \N_WR_USB_ADBUS_0_iv_5[4]\);
    
    \ELINK_ADDRA_3[0]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[0]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_1, E => un1_SM_BANK_SEL_4, Q => 
        \ELINK_ADDRA_3[0]_net_1\);
    
    \ELINK_ADDRA_11[4]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[4]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_2, E => un1_SM_BANK_SEL_16, Q => 
        \ELINK_ADDRA_11[4]_net_1\);
    
    \RD_USB_ADBUS_RNI7HSK4[7]\ : NOR3C
      port map(A => N_465, B => N_1367_i_i_a2_2, C => 
        N_1367_i_i_a2_3, Y => N_480);
    
    \ELINK_ADDRA_13[0]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[0]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_3, E => un1_SM_BANK_SEL_2, Q => 
        \ELINK_ADDRA_13[0]_net_1\);
    
    \TFC_STRT_ADDR[6]\ : DFN1E1C0
      port map(D => \TFC_STRT_ADDR_T[6]_net_1\, CLK => CLK60MHZ, 
        CLR => P_USB_MASTER_EN_c_13, E => \REG_STATE_d_0[30]\, Q
         => \TFC_STRT_ADDR[6]_net_1\);
    
    \WR_XFER_TYPE[0]\ : DFN1C0
      port map(D => \WR_XFER_TYPE_RNO[0]_net_1\, CLK => CLK60MHZ, 
        CLR => P_USB_MASTER_EN_c, Q => \WR_XFER_TYPE[0]_net_1\);
    
    \REG_STATE_RNI6VOT[2]\ : NOR2A
      port map(A => N_2613, B => \REG_STATE[2]_net_1\, Y => 
        \REG_STATE_ns_i_a4_7_0[4]\);
    
    \ELINK_BLKA_RNO_0[9]\ : NOR2B
      port map(A => \SM_BANK_SEL[10]_net_1\, B => X_BLKA_i, Y => 
        N_164);
    
    \REG_STATE[4]\ : DFN1C0
      port map(D => \REG_STATE_RNIMO53U3[2]_net_1\, CLK => 
        CLK60MHZ, CLR => P_USB_MASTER_EN_c_22_0, Q => 
        \REG_STATE[4]_net_1\);
    
    \SM_BANK_SEL[19]\ : DFN1E1C0
      port map(D => N_1848, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_1_0, E => un1_REG_STATE_30, Q => 
        \SM_BANK_SEL[19]_net_1\);
    
    \ELINK_ADDRA_4[3]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[3]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_2_0, E => un1_SM_BANK_SEL_8, Q => 
        \ELINK_ADDRA_4[3]_net_1\);
    
    \WR_XFER_TYPE_RNO_1[0]\ : NOR3A
      port map(A => \RD_USB_ADBUS[1]_net_1\, B => 
        \WR_XFER_TYPE[0]_net_1\, C => \RD_USB_ADBUS[5]_net_1\, Y
         => N_1818);
    
    \REG_STATE_RNIU1LF1[0]\ : NOR2
      port map(A => N_1739, B => N_268, Y => N_1351_8);
    
    \REG_STATE_RNI0SAF5[4]\ : OR3
      port map(A => N_2570, B => N_1877_1, C => N_2566, Y => 
        \REG_STATE_ns_i_1[4]\);
    
    \ELINK_DINA_13[3]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[3]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_14, E => un1_SM_BANK_SEL_2, Q => 
        \ELINK_DINA_13[3]_net_1\);
    
    \WR_USB_ADBUS_RNO_9[1]\ : AO1
      port map(A => \ELINK_DOUTA_7[1]\, B => un1_SM_BANK_SEL_37, 
        C => \ELINK_DOUTA_9_m[1]\, Y => 
        \N_WR_USB_ADBUS_0_iv_14[1]\);
    
    \REG_STATE_RNITEQN_1[0]\ : NOR2A
      port map(A => \REG_STATE[1]_net_1\, B => 
        \REG_STATE[0]_net_1\, Y => N_1352_1);
    
    \ELINK_ADDRA_19[4]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[4]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_13, E => un1_SM_BANK_SEL_11, Q => 
        \ELINK_ADDRA_19[4]_net_1\);
    
    \WR_USB_ADBUS_RNO_37[5]\ : NOR2B
      port map(A => \ELINK_DOUTA_13[5]\, B => un1_SM_BANK_SEL_29, 
        Y => \ELINK_DOUTA_13_m[5]\);
    
    \SM_BANK_SEL_RNICN9D[8]\ : NOR2A
      port map(A => N_469, B => \SM_BANK_SEL[8]_net_1\, Y => 
        N_365);
    
    \REG_STATE_RNIVGQN_1[0]\ : OR2A
      port map(A => \REG_STATE[3]_net_1\, B => 
        \REG_STATE[0]_net_1\, Y => N_287);
    
    \ELINK_ADDRA_9[1]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[1]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_10, E => un1_SM_BANK_SEL_9, Q => 
        \ELINK_ADDRA_9[1]_net_1\);
    
    \ELINK_BLKA_RNO[11]\ : OA1B
      port map(A => N_393, B => \ELINK_BLKA[11]_net_1\, C => 
        N_162, Y => \N_ELINK_BLKA_0_iv[11]\);
    
    \ELINKS_STRT_ADDR_T[6]\ : DFN1E1C0
      port map(D => \RD_USB_ADBUS[6]_net_1\, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_21, E => 
        N_ELINKS_STRT_ADDR_T_0_sqmuxa, Q => 
        \ELINKS_STRT_ADDR_T[6]_net_1\);
    
    \WR_USB_ADBUS_RNO_34[2]\ : NOR2B
      port map(A => \ELINK_DOUTA_19[2]\, B => un1_SM_BANK_SEL_41, 
        Y => \ELINK_DOUTA_19_m[2]\);
    
    \TFC_STRT_ADDR[2]\ : DFN1E1C0
      port map(D => \TFC_STRT_ADDR_T[2]_net_1\, CLK => CLK60MHZ, 
        CLR => P_USB_MASTER_EN_c_13, E => \REG_STATE_d_0[30]\, Q
         => \TFC_STRT_ADDR[2]_net_1\);
    
    \REG_STATE_RNIR359F1[2]\ : OR3A
      port map(A => N_264, B => \REG_STATE_ns_i_1[4]\, C => 
        \REG_STATE_ns_i_8[4]\, Y => \REG_STATE_ns_i_3[4]\);
    
    \REG_STATE_ns_i_i_o2_6_1_RNO_3[0]\ : NOR2A
      port map(A => N_274, B => N_287, Y => N_450);
    
    USB_RXF_B_0_RNI1JC64 : AO1D
      port map(A => N_1694, B => \USB_RXF_B_0\, C => N_675_0, Y
         => N_1737);
    
    un1_REG_STATE_4_0_a2 : AND2
      port map(A => N_1690_i, B => un1_REG_STATE_4_0_a2_1, Y => 
        N_1781);
    
    \SM_BANK_SEL_RNO[10]\ : NOR3B
      port map(A => N_1892, B => N_1351_4, C => 
        \RD_USB_ADBUS[2]_net_1\, Y => N_1839);
    
    \WR_USB_ADBUS_RNO_13[1]\ : NOR2B
      port map(A => \ELINK_DOUTA_1[1]\, B => un1_SM_BANK_SEL_36, 
        Y => \ELINK_DOUTA_1_m[1]\);
    
    \REG_STATE_RNI0DIR1[4]\ : OR2
      port map(A => N_1691, B => N_2497, Y => N_1694);
    
    \ELINK_ADDRA_0[2]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[2]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_18, E => un1_SM_BANK_SEL_6, Q => 
        \ELINK_ADDRA_0[2]_net_1\);
    
    \ELINK_ADDRA_16[4]\ : DFN1E0C0
      port map(D => \N_TFC_ADDRA[4]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_8, E => N_200, Q => 
        \ELINK_ADDRA_16[4]_net_1\);
    
    \WR_USB_ADBUS_RNO_30[5]\ : NOR3B
      port map(A => N_1730_i, B => \ELINKS_STOP_ADDR[5]_net_1\, C
         => N_1726, Y => \ELINKS_STOP_ADDR_m[5]\);
    
    USB_RXF_B_0_RNI27AB1_1 : NOR3
      port map(A => \REG_STATE_0[3]_net_1\, B => \USB_RXF_B_0\, C
         => \REG_STATE_0[4]_net_1\, Y => 
        \REG_STATE_ns_i_a4_6_1[4]\);
    
    \SM_BANK_SEL_RNIEV0C2[4]\ : NOR3A
      port map(A => \SM_BANK_SEL[4]_net_1\, B => N_312_0, C => 
        N_1566_i_i_0, Y => un1_SM_BANK_SEL_24);
    
    \WR_USB_ADBUS_RNO_6[2]\ : NOR2B
      port map(A => \ELINK_DOUTA_15[2]\, B => un1_SM_BANK_SEL_24, 
        Y => \ELINK_DOUTA_15_m[2]\);
    
    \WR_USB_ADBUS_RNO[6]\ : OR3
      port map(A => \N_WR_USB_ADBUS_0_iv_23[6]\, B => 
        \N_WR_USB_ADBUS_0_iv_22[6]\, C => 
        \N_WR_USB_ADBUS_0_iv_24[6]\, Y => \N_WR_USB_ADBUS[6]\);
    
    \REG_STATE_RNIM3OI[5]\ : NOR2A
      port map(A => \REG_STATE[5]_net_1\, B => \USB_TXE_B\, Y => 
        N_433_1);
    
    \REG_ADDR[3]\ : DFN1E1C0
      port map(D => REG_ADDR_n3, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_10, E => REG_ADDRe, Q => 
        \REG_ADDR[3]_net_1\);
    
    \RD_USB_ADBUS_RNI2S3U2[5]\ : OA1
      port map(A => \RD_USB_ADBUS[5]_net_1\, B => N_1881, C => 
        un1_REG_STATE_39_i_a2_0, Y => N_1862);
    
    \REG_STATE_ns_i_i_o2_6_1_RNO_2[0]\ : NOR2
      port map(A => \REG_STATE[5]_net_1\, B => N_292, Y => 
        \REG_STATE_ns_i_i_a2_5_0[0]\);
    
    \ELINK_BLKA_RNO[5]\ : AOI1
      port map(A => \SM_BANK_SEL[14]_net_1\, B => X_BLKA_i, C => 
        N_165, Y => \N_ELINK_BLKA_0_iv[5]\);
    
    \WR_USB_ADBUS_RNO_17[3]\ : AO1A
      port map(A => N_1497, B => \TFC_STRT_ADDR[3]_net_1\, C => 
        \ELINKS_STOP_ADDR_m[3]\, Y => \N_WR_USB_ADBUS_0_iv_3[3]\);
    
    \REG_ADDR_RNIKLPL[8]\ : NOR3A
      port map(A => \REG_ADDR[8]_net_1\, B => \REG_ADDR[1]_net_1\, 
        C => \REG_ADDR[3]_net_1\, Y => REG_STATE_tr73_4);
    
    \ELINK_ADDRA_4[0]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[0]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_2, E => un1_SM_BANK_SEL_8, Q => 
        \ELINK_ADDRA_4[0]_net_1\);
    
    \ELINK_ADDRA_16[5]\ : DFN1E0C0
      port map(D => \N_TFC_ADDRA[5]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_9, E => N_200, Q => 
        \ELINK_ADDRA_16[5]_net_1\);
    
    \WR_USB_ADBUS_RNO_18[0]\ : NOR2B
      port map(A => \ELINK_DOUTA_5[0]\, B => un1_SM_BANK_SEL_35, 
        Y => \ELINK_DOUTA_5_m[0]\);
    
    \ELINK_DINA_3[5]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[5]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_11, E => un1_SM_BANK_SEL_4, Q => 
        \ELINK_DINA_3[5]_net_1\);
    
    \ELINK_ADDRA_8[6]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[6]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_8, E => un1_SM_BANK_SEL_21, Q => 
        \ELINK_ADDRA_8[6]_net_1\);
    
    \REG_STATE_RNI1JQN[3]\ : OR2A
      port map(A => \REG_STATE[2]_net_1\, B => 
        \REG_STATE[3]_net_1\, Y => N_268);
    
    \REG_STATE_0_RNIF9MT1_0[4]\ : NOR3B
      port map(A => N_1359_2, B => N_1352_1, C => 
        \REG_STATE_0[4]_net_1\, Y => \REG_STATE_d_0[30]\);
    
    U113_PATT_ELINK_BLK : DPRT_512X9_SRAM_13
      port map(ELINK_RWA_0 => \ELINK_RWA[13]_net_1\, 
        ELK_RX_SER_WORD_13(7) => ELK_RX_SER_WORD_13(7), 
        ELK_RX_SER_WORD_13(6) => ELK_RX_SER_WORD_13(6), 
        ELK_RX_SER_WORD_13(5) => ELK_RX_SER_WORD_13(5), 
        ELK_RX_SER_WORD_13(4) => ELK_RX_SER_WORD_13(4), 
        ELK_RX_SER_WORD_13(3) => ELK_RX_SER_WORD_13(3), 
        ELK_RX_SER_WORD_13(2) => ELK_RX_SER_WORD_13(2), 
        ELK_RX_SER_WORD_13(1) => ELK_RX_SER_WORD_13(1), 
        ELK_RX_SER_WORD_13(0) => ELK_RX_SER_WORD_13(0), 
        ELINK_DINA_13(7) => \ELINK_DINA_13[7]_net_1\, 
        ELINK_DINA_13(6) => \ELINK_DINA_13[6]_net_1\, 
        ELINK_DINA_13(5) => \ELINK_DINA_13[5]_net_1\, 
        ELINK_DINA_13(4) => \ELINK_DINA_13[4]_net_1\, 
        ELINK_DINA_13(3) => \ELINK_DINA_13[3]_net_1\, 
        ELINK_DINA_13(2) => \ELINK_DINA_13[2]_net_1\, 
        ELINK_DINA_13(1) => \ELINK_DINA_13[1]_net_1\, 
        ELINK_DINA_13(0) => \ELINK_DINA_13[0]_net_1\, 
        ELINK_BLKA_0 => \ELINK_BLKA[13]_net_1\, ELKS_ADDRB_0_d0
         => ELKS_ADDRB(0), ELKS_ADDRB_1 => ELKS_ADDRB(1), 
        ELKS_ADDRB_3 => ELKS_ADDRB(3), ELKS_ADDRB_5 => 
        ELKS_ADDRB(5), ELKS_ADDRB_7 => ELKS_ADDRB(7), 
        ELKS_ADDRB_0_0 => ELKS_ADDRB_0_0, ELKS_ADDRB_0_2 => 
        ELKS_ADDRB_0_2, ELKS_ADDRB_0_4 => ELKS_ADDRB_0_4, 
        ELINK_ADDRA_13(7) => \ELINK_ADDRA_13[7]_net_1\, 
        ELINK_ADDRA_13(6) => \ELINK_ADDRA_13[6]_net_1\, 
        ELINK_ADDRA_13(5) => \ELINK_ADDRA_13[5]_net_1\, 
        ELINK_ADDRA_13(4) => \ELINK_ADDRA_13[4]_net_1\, 
        ELINK_ADDRA_13(3) => \ELINK_ADDRA_13[3]_net_1\, 
        ELINK_ADDRA_13(2) => \ELINK_ADDRA_13[2]_net_1\, 
        ELINK_ADDRA_13(1) => \ELINK_ADDRA_13[1]_net_1\, 
        ELINK_ADDRA_13(0) => \ELINK_ADDRA_13[0]_net_1\, 
        PATT_ELK_DAT_13(7) => PATT_ELK_DAT_13(7), 
        PATT_ELK_DAT_13(6) => PATT_ELK_DAT_13(6), 
        PATT_ELK_DAT_13(5) => PATT_ELK_DAT_13(5), 
        PATT_ELK_DAT_13(4) => PATT_ELK_DAT_13(4), 
        PATT_ELK_DAT_13(3) => PATT_ELK_DAT_13(3), 
        PATT_ELK_DAT_13(2) => PATT_ELK_DAT_13(2), 
        PATT_ELK_DAT_13(1) => PATT_ELK_DAT_13(1), 
        PATT_ELK_DAT_13(0) => PATT_ELK_DAT_13(0), 
        ELINK_DOUTA_13(7) => \ELINK_DOUTA_13[7]\, 
        ELINK_DOUTA_13(6) => \ELINK_DOUTA_13[6]\, 
        ELINK_DOUTA_13(5) => \ELINK_DOUTA_13[5]\, 
        ELINK_DOUTA_13(4) => \ELINK_DOUTA_13[4]\, 
        ELINK_DOUTA_13(3) => \ELINK_DOUTA_13[3]\, 
        ELINK_DOUTA_13(2) => \ELINK_DOUTA_13[2]\, 
        ELINK_DOUTA_13(1) => \ELINK_DOUTA_13[1]\, 
        ELINK_DOUTA_13(0) => \ELINK_DOUTA_13[0]\, ELKS_RWB => 
        ELKS_RWB, P_USB_MASTER_EN_c_0 => P_USB_MASTER_EN_c_0, 
        CLK_40M_GL => CLK_40M_GL, CLK60MHZ => CLK60MHZ, 
        ELKS_RAM_BLKB_EN => ELKS_RAM_BLKB_EN);
    
    \SI_CNT[0]\ : DFN1E1C0
      port map(D => N_2625, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_5, E => SI_CNTe, Q => \SI_CNT[0]_net_1\);
    
    \REG_STATE_0_RNI6SJO1[5]\ : NOR3A
      port map(A => N_312, B => N_339, C => 
        \REG_STATE_0[5]_net_1\, Y => N_2539);
    
    USB_TXE_B_RNIKF203 : OA1
      port map(A => REG_STATE_tr74_tz_tz_tz_5, B => 
        REG_STATE_tr74_tz_tz_tz_6, C => REG_STATE_tr74_0, Y => 
        REG_STATE_tr74_1);
    
    \RD_XFER_TYPE_RNO[7]\ : AO1
      port map(A => \RD_XFER_TYPE[7]_net_1\, B => N_1703, C => 
        N_1808, Y => \RD_XFER_TYPE_RNO[7]_net_1\);
    
    \ELINK_RWA[6]\ : DFN1E0P0
      port map(D => \N_ELINK_RWA_0_iv[6]\, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_6, E => \SM_BANK_SEL_0[20]_net_1\, 
        Q => \ELINK_RWA[6]_net_1\);
    
    \ELINK_BLKA[7]\ : DFN1E0P0
      port map(D => \N_ELINK_BLKA_0_iv[7]\, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_19, E => \SM_BANK_SEL[20]_net_1\, Q
         => \ELINK_BLKA[7]_net_1\);
    
    USB_RXF_B_RNIQMBQL : AO1
      port map(A => N_510, B => N_285, C => N_471, Y => N_311);
    
    \REG_STATE_0_RNISQSJ1_0[1]\ : NOR3
      port map(A => \REG_STATE_0[2]_net_1\, B => 
        \REG_STATE_0[1]_net_1\, C => N_287, Y => N_2546);
    
    \RD_XFER_TYPE_RNO[6]\ : AO1
      port map(A => \RD_XFER_TYPE[6]_net_1\, B => N_1703, C => 
        N_1806, Y => \RD_XFER_TYPE_RNO[6]_net_1\);
    
    \RD_XFER_TYPE_RNO_0[3]\ : NOR2A
      port map(A => \RD_USB_ADBUS[3]_net_1\, B => N_1694, Y => 
        N_1800);
    
    \ELINK_ADDRA_19[7]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[7]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_13, E => un1_SM_BANK_SEL_11, Q => 
        \ELINK_ADDRA_19[7]_net_1\);
    
    \ELINK_ADDRA_7[2]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[2]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_6, E => un1_SM_BANK_SEL_12, Q => 
        \ELINK_ADDRA_7[2]_net_1\);
    
    \RD_USB_ADBUS_RNIQO682[6]\ : NOR3C
      port map(A => N_1351_3, B => N_459, C => N_1367_i_i_a2_0, Y
         => N_1367_i_i_a2_2);
    
    \ELINK_ADDRA_1[3]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[3]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_20, E => un1_SM_BANK_SEL_19, Q => 
        \ELINK_ADDRA_1[3]_net_1\);
    
    \WR_USB_ADBUS_RNO_35[1]\ : NOR2B
      port map(A => \ELINK_DOUTA_0[1]\, B => un1_SM_BANK_SEL_31, 
        Y => \ELINK_DOUTA_0_m[1]\);
    
    \RD_USB_ADBUS_RNISGIK2[7]\ : NOR2A
      port map(A => \RD_USB_ADBUS[7]_net_1\, B => N_206, Y => 
        \N_TFC_DINA[7]\);
    
    \RD_XFER_TYPE_RNO[5]\ : AO1
      port map(A => \RD_XFER_TYPE[5]_net_1\, B => N_1703, C => 
        N_1804, Y => \RD_XFER_TYPE_RNO[5]_net_1\);
    
    \ELINK_DINA_3[4]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[4]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_11, E => un1_SM_BANK_SEL_4, Q => 
        \ELINK_DINA_3[4]_net_1\);
    
    \ELINK_ADDRA_10[5]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[5]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_22, E => un1_SM_BANK_SEL_20, Q => 
        \ELINK_ADDRA_10[5]_net_1\);
    
    \N_TFC_ADDRA_0_o2_RNO_7[7]\ : MX2A
      port map(A => \REG_STATE_0[0]_net_1\, B => 
        \REG_STATE_0[4]_net_1\, S => \REG_STATE_0[1]_net_1\, Y
         => N_259);
    
    \CHKSUM[4]\ : DFN1E1C0
      port map(D => N_232, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_3, E => un1_REG_STATE_22, Q => 
        \CHKSUM[4]_net_1\);
    
    \WR_USB_ADBUS_RNO_1[0]\ : OR3
      port map(A => \N_WR_USB_ADBUS_0_iv_8[0]\, B => 
        \N_WR_USB_ADBUS_0_iv_7[0]\, C => 
        \N_WR_USB_ADBUS_0_iv_17[0]\, Y => 
        \N_WR_USB_ADBUS_0_iv_23[0]\);
    
    \RD_USB_ADBUS_RNIRVAJ_0[0]\ : OR2B
      port map(A => \RD_USB_ADBUS[0]_net_1\, B => 
        \RD_USB_ADBUS[1]_net_1\, Y => N_290);
    
    \WR_USB_ADBUS[7]\ : DFN1E0C0
      port map(D => \N_WR_USB_ADBUS[7]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_15, E => un1_REG_STATE_26, Q => 
        \WR_USB_ADBUS[7]_net_1\);
    
    \ELINK_RWA_RNO_0[0]\ : OA1B
      port map(A => N_616_16, B => \N_ELINK_RWA_3[0]\, C => 
        \ELINK_RWA[0]_net_1\, Y => \ELINK_RWA_i_m[0]\);
    
    \TFC_STOP_ADDR[3]\ : DFN1E1C0
      port map(D => \TFC_STOP_ADDR_T[3]_net_1\, CLK => CLK60MHZ, 
        CLR => P_USB_MASTER_EN_c_8, E => \REG_STATE_d_0[30]\, Q
         => \TFC_STOP_ADDR[3]_net_1\);
    
    \WR_USB_ADBUS_RNO_34[3]\ : NOR2B
      port map(A => \CHKSUM[3]_net_1\, B => un1_REG_STATE_4, Y
         => \CHKSUM_m[3]\);
    
    \WR_USB_ADBUS_RNO_27[0]\ : NOR2B
      port map(A => \ELINK_DOUTA_19[0]\, B => un1_SM_BANK_SEL_41, 
        Y => \ELINK_DOUTA_19_m[0]\);
    
    \WR_USB_ADBUS_RNO_25[2]\ : OR3
      port map(A => \N_WR_USB_ADBUS_0_iv_0[2]_net_1\, B => 
        \OP_MODE_m[2]\, C => \ELINKS_STRT_ADDR_m[2]\, Y => 
        \N_WR_USB_ADBUS_0_iv_2[2]\);
    
    \SM_BANK_SEL_RNIU2E6[16]\ : OR3
      port map(A => N_616_2, B => N_618_1, C => N_616_11, Y => 
        \N_ELINK_RWA_1[2]\);
    
    \REG_ADDR_RNO_0[2]\ : AX1E
      port map(A => \REG_ADDR[0]_net_1\, B => \REG_ADDR[1]_net_1\, 
        C => \REG_ADDR[2]_net_1\, Y => REG_ADDR_n2_i_0);
    
    \OP_MODE_T[3]\ : DFN1E1C0
      port map(D => \RD_USB_ADBUS[3]_net_1\, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_17, E => N_OP_MODE_T_0_sqmuxa, Q
         => \OP_MODE_T[3]_net_1\);
    
    \WR_XFER_TYPE_RNO[4]\ : NOR3B
      port map(A => N_1763, B => N_1716, C => N_1827, Y => 
        \WR_XFER_TYPE_RNO[4]_net_1\);
    
    \REG_STATE_0_RNI6SJO1_0[5]\ : AO1A
      port map(A => N_287, B => \REG_STATE_0[5]_net_1\, C => 
        N_1749, Y => un1_REG_STATE_26_0_0);
    
    \ELINK_BLKA[14]\ : DFN1E0P0
      port map(D => \N_ELINK_BLKA_0_iv[14]\, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_20, E => \SM_BANK_SEL[20]_net_1\, Q
         => \ELINK_BLKA[14]_net_1\);
    
    \WR_USB_ADBUS_RNO_21[3]\ : NOR2B
      port map(A => \ELINK_DOUTA_19[3]\, B => un1_SM_BANK_SEL_41, 
        Y => \ELINK_DOUTA_19_m[3]\);
    
    \REG_STATE_ns_i_i_a2_0_2_RNO_1[0]\ : NOR3A
      port map(A => N_1778, B => N_292, C => N_1359_1, Y => N_413);
    
    \REG_ADDR_RNIQVCP[7]\ : NOR3B
      port map(A => N_261, B => \REG_ADDR[7]_net_1\, C => 
        \SM_BANK_SEL_0[21]_net_1\, Y => \N_TFC_ADDRA[7]\);
    
    \ELINK_BLKA[18]\ : DFN1E0P0
      port map(D => N_63, CLK => CLK60MHZ, PRE => 
        P_USB_MASTER_EN_c_20, E => \SM_BANK_SEL[20]_net_1\, Q => 
        \ELINK_BLKA[18]_net_1\);
    
    \ELINK_DINA_4[5]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[5]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_13, E => un1_SM_BANK_SEL_8, Q => 
        \ELINK_DINA_4[5]_net_1\);
    
    \ELINK_ADDRA_15[4]\ : DFN1E0C0
      port map(D => \N_TFC_ADDRA[4]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_6, E => N_199, Q => 
        \ELINK_ADDRA_15[4]_net_1\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \ELINK_ADDRA_3[2]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[2]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_1, E => un1_SM_BANK_SEL_4, Q => 
        \ELINK_ADDRA_3[2]_net_1\);
    
    \SM_BANK_SEL_RNILRL6[6]\ : OR2
      port map(A => \SM_BANK_SEL[6]_net_1\, B => 
        \SM_BANK_SEL[21]_net_1\, Y => un1_SM_BANK_SEL_2);
    
    \REG_STATE_0_RNIKIRD2[3]\ : OR2
      port map(A => N_2622, B => \REG_STATE_ns_i_a4_1_0[3]\, Y
         => N_1259_tz);
    
    U112_PATT_ELINK_BLK : DPRT_512X9_SRAM_12
      port map(ELINK_RWA_0 => \ELINK_RWA[12]_net_1\, 
        ELK_RX_SER_WORD_12(7) => ELK_RX_SER_WORD_12(7), 
        ELK_RX_SER_WORD_12(6) => ELK_RX_SER_WORD_12(6), 
        ELK_RX_SER_WORD_12(5) => ELK_RX_SER_WORD_12(5), 
        ELK_RX_SER_WORD_12(4) => ELK_RX_SER_WORD_12(4), 
        ELK_RX_SER_WORD_12(3) => ELK_RX_SER_WORD_12(3), 
        ELK_RX_SER_WORD_12(2) => ELK_RX_SER_WORD_12(2), 
        ELK_RX_SER_WORD_12(1) => ELK_RX_SER_WORD_12(1), 
        ELK_RX_SER_WORD_12(0) => ELK_RX_SER_WORD_12(0), 
        ELINK_DINA_12(7) => \ELINK_DINA_12[7]_net_1\, 
        ELINK_DINA_12(6) => \ELINK_DINA_12[6]_net_1\, 
        ELINK_DINA_12(5) => \ELINK_DINA_12[5]_net_1\, 
        ELINK_DINA_12(4) => \ELINK_DINA_12[4]_net_1\, 
        ELINK_DINA_12(3) => \ELINK_DINA_12[3]_net_1\, 
        ELINK_DINA_12(2) => \ELINK_DINA_12[2]_net_1\, 
        ELINK_DINA_12(1) => \ELINK_DINA_12[1]_net_1\, 
        ELINK_DINA_12(0) => \ELINK_DINA_12[0]_net_1\, 
        ELINK_BLKA_0 => \ELINK_BLKA[12]_net_1\, ELKS_ADDRB_0_d0
         => ELKS_ADDRB(0), ELKS_ADDRB_1 => ELKS_ADDRB(1), 
        ELKS_ADDRB_3 => ELKS_ADDRB(3), ELKS_ADDRB_5 => 
        ELKS_ADDRB(5), ELKS_ADDRB_7 => ELKS_ADDRB(7), 
        ELKS_ADDRB_0_0 => ELKS_ADDRB_0_0, ELKS_ADDRB_0_2 => 
        ELKS_ADDRB_0_2, ELKS_ADDRB_0_4 => ELKS_ADDRB_0_4, 
        ELINK_ADDRA_12(7) => \ELINK_ADDRA_12[7]_net_1\, 
        ELINK_ADDRA_12(6) => \ELINK_ADDRA_12[6]_net_1\, 
        ELINK_ADDRA_12(5) => \ELINK_ADDRA_12[5]_net_1\, 
        ELINK_ADDRA_12(4) => \ELINK_ADDRA_12[4]_net_1\, 
        ELINK_ADDRA_12(3) => \ELINK_ADDRA_12[3]_net_1\, 
        ELINK_ADDRA_12(2) => \ELINK_ADDRA_12[2]_net_1\, 
        ELINK_ADDRA_12(1) => \ELINK_ADDRA_12[1]_net_1\, 
        ELINK_ADDRA_12(0) => \ELINK_ADDRA_12[0]_net_1\, 
        PATT_ELK_DAT_12(7) => PATT_ELK_DAT_12(7), 
        PATT_ELK_DAT_12(6) => PATT_ELK_DAT_12(6), 
        PATT_ELK_DAT_12(5) => PATT_ELK_DAT_12(5), 
        PATT_ELK_DAT_12(4) => PATT_ELK_DAT_12(4), 
        PATT_ELK_DAT_12(3) => PATT_ELK_DAT_12(3), 
        PATT_ELK_DAT_12(2) => PATT_ELK_DAT_12(2), 
        PATT_ELK_DAT_12(1) => PATT_ELK_DAT_12(1), 
        PATT_ELK_DAT_12(0) => PATT_ELK_DAT_12(0), 
        ELINK_DOUTA_12(7) => \ELINK_DOUTA_12[7]\, 
        ELINK_DOUTA_12(6) => \ELINK_DOUTA_12[6]\, 
        ELINK_DOUTA_12(5) => \ELINK_DOUTA_12[5]\, 
        ELINK_DOUTA_12(4) => \ELINK_DOUTA_12[4]\, 
        ELINK_DOUTA_12(3) => \ELINK_DOUTA_12[3]\, 
        ELINK_DOUTA_12(2) => \ELINK_DOUTA_12[2]\, 
        ELINK_DOUTA_12(1) => \ELINK_DOUTA_12[1]\, 
        ELINK_DOUTA_12(0) => \ELINK_DOUTA_12[0]\, ELKS_RWB => 
        ELKS_RWB, P_USB_MASTER_EN_c_0 => P_USB_MASTER_EN_c_0, 
        CLK_40M_GL => CLK_40M_GL, CLK60MHZ => CLK60MHZ, 
        ELKS_RAM_BLKB_EN => ELKS_RAM_BLKB_EN);
    
    \WR_USB_ADBUS_RNO_1[6]\ : OR3
      port map(A => \N_WR_USB_ADBUS_0_iv_7[6]\, B => 
        \N_WR_USB_ADBUS_0_iv_6[6]\, C => 
        \N_WR_USB_ADBUS_0_iv_16[6]\, Y => 
        \N_WR_USB_ADBUS_0_iv_22[6]\);
    
    \ELINK_ADDRA_4[1]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[1]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_2, E => un1_SM_BANK_SEL_8, Q => 
        \ELINK_ADDRA_4[1]_net_1\);
    
    \ELINK_ADDRA_11[5]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[5]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_2, E => un1_SM_BANK_SEL_16, Q => 
        \ELINK_ADDRA_11[5]_net_1\);
    
    \WR_USB_ADBUS_RNO_28[7]\ : NOR2B
      port map(A => \ELINK_DOUTA_5[7]\, B => un1_SM_BANK_SEL_35, 
        Y => \ELINK_DOUTA_5_m[7]\);
    
    \TFC_STRT_ADDR[7]\ : DFN1E1C0
      port map(D => \TFC_STRT_ADDR_T[7]_net_1\, CLK => CLK60MHZ, 
        CLR => P_USB_MASTER_EN_c_13, E => \REG_STATE_d_0[30]\, Q
         => \TFC_STRT_ADDR[7]_net_1\);
    
    \ELINK_ADDRA_18[6]\ : DFN1E0C0
      port map(D => \N_TFC_ADDRA[6]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_12, E => N_198, Q => 
        \ELINK_ADDRA_18[6]_net_1\);
    
    \SM_BANK_SEL[5]\ : DFN1E1C0
      port map(D => N_1845, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_7, E => un1_REG_STATE_30, Q => 
        \SM_BANK_SEL[5]_net_1\);
    
    \RD_USB_ADBUS_RNIR0NJ3[6]\ : NOR2A
      port map(A => \REG_STATE_ns_i_i_a5_1_2[0]\, B => N_282, Y
         => \REG_STATE_ns_i_i_a5_1_3[0]\);
    
    \ELINK_ADDRA_6[7]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[7]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_4, E => un1_SM_BANK_SEL_10, Q => 
        \ELINK_ADDRA_6[7]_net_1\);
    
    \ELINK_ADDRA_2[5]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[5]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_21, E => un1_SM_BANK_SEL_5, Q => 
        \ELINK_ADDRA_2[5]_net_1\);
    
    USB_TXE_B_RNIV2O4Q : OR2B
      port map(A => N_2581, B => N_2454_tz, Y => 
        \USB_TXE_B_RNIV2O4Q\);
    
    \ELINK_DINA_10[2]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[2]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_9, E => un1_SM_BANK_SEL_20, Q => 
        \ELINK_DINA_10[2]_net_1\);
    
    \CHKSUM[7]\ : DFN1E1C0
      port map(D => N_226, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_4, E => un1_REG_STATE_22, Q => 
        \CHKSUM[7]_net_1\);
    
    \WR_USB_ADBUS_RNO_22[4]\ : NOR2B
      port map(A => \ELINK_DOUTA_16[4]\, B => un1_SM_BANK_SEL_39, 
        Y => \ELINK_DOUTA_16_m[4]\);
    
    \WR_XFER_TYPE[3]\ : DFN1C0
      port map(D => \WR_XFER_TYPE_RNO[3]_net_1\, CLK => CLK60MHZ, 
        CLR => P_USB_MASTER_EN_c, Q => \WR_XFER_TYPE[3]_net_1\);
    
    \WR_USB_ADBUS_RNO_1[2]\ : OR3
      port map(A => \ELINK_DOUTA_15_m[2]\, B => \TFC_DOUTA_m[2]\, 
        C => \N_WR_USB_ADBUS_0_iv_14[2]\, Y => 
        \N_WR_USB_ADBUS_0_iv_21[2]\);
    
    \REG_ADDR_RNIV1JB1[5]\ : NOR2B
      port map(A => REG_ADDR_c4, B => \REG_ADDR[5]_net_1\, Y => 
        REG_ADDR_c5);
    
    \REG_STATE_RNI3LQN[3]\ : OR2B
      port map(A => \REG_STATE[3]_net_1\, B => 
        \REG_STATE[4]_net_1\, Y => N_1726);
    
    \ELINK_DINA_9[2]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[2]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_19, E => un1_SM_BANK_SEL_9, Q => 
        \ELINK_DINA_9[2]_net_1\);
    
    \CHKSUM[0]\ : DFN1E1C0
      port map(D => N_1593, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_3, E => un1_REG_STATE_22, Q => 
        \CHKSUM[0]_net_1\);
    
    \REG_STATE_0_RNI5OTL2[5]\ : OA1A
      port map(A => \REG_STATE_0[4]_net_1\, B => N_2577, C => 
        \REG_STATE_0[5]_net_1\, Y => N_457);
    
    \SM_BANK_SEL_RNID1N12[0]\ : NOR3C
      port map(A => N_463, B => N_464, C => 
        \N_ELINK_BLKA_0_iv_0_o2_i_a5_2[9]\, Y => N_392);
    
    \ELINK_DINA_6[3]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[3]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_16, E => un1_SM_BANK_SEL_10, Q => 
        \ELINK_DINA_6[3]_net_1\);
    
    \WR_USB_ADBUS[1]\ : DFN1E0C0
      port map(D => \N_WR_USB_ADBUS[1]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_15, E => un1_REG_STATE_26, Q => 
        \WR_USB_ADBUS[1]_net_1\);
    
    \ELINK_RWA[3]\ : DFN1E0P0
      port map(D => \N_ELINK_RWA_0_iv[3]\, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_6, E => \SM_BANK_SEL_0[20]_net_1\, 
        Q => \ELINK_RWA[3]_net_1\);
    
    \SM_BANK_SEL_RNIGML6[1]\ : NOR2
      port map(A => \SM_BANK_SEL[1]_net_1\, B => 
        \SM_BANK_SEL[21]_net_1\, Y => N_198);
    
    ELK_N_ACTIVE_RNIGTNG9 : NOR3C
      port map(A => N_480, B => N_277, C => N_256, Y => N_384);
    
    \ELINK_ADDRA_17[0]\ : DFN1E0C0
      port map(D => \N_TFC_ADDRA[0]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_10, E => N_197, Q => 
        \ELINK_ADDRA_17[0]_net_1\);
    
    \REG_STATE_0_RNIT92S[0]\ : OR2A
      port map(A => \REG_STATE_0[0]_net_1\, B => 
        \REG_STATE_0[3]_net_1\, Y => N_312_0);
    
    \REG_STATE_RNIKJIA1[0]\ : NOR2A
      port map(A => N_2571_1, B => N_339, Y => 
        \REG_STATE_ns_i_a4_8_0_a5_0[4]\);
    
    \SM_BANK_SEL[1]\ : DFN1E1C0
      port map(D => N_1850, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_7, E => un1_REG_STATE_30, Q => 
        \SM_BANK_SEL[1]_net_1\);
    
    \REG_STATE_0_RNIFS5H2[5]\ : NOR3A
      port map(A => N_2498, B => \REG_STATE_0[5]_net_1\, C => 
        N_312, Y => \REG_STATE_ns_i_a4_0[4]\);
    
    \ELINK_DINA_3[1]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[1]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_11, E => un1_SM_BANK_SEL_4, Q => 
        \ELINK_DINA_3[1]_net_1\);
    
    \SI_CNT_RNI5TT8[3]\ : NOR2B
      port map(A => \SI_CNT[3]_net_1\, B => \SI_CNT[2]_net_1\, Y
         => \REG_STATE_ns_i_a2_2_0[4]\);
    
    \ELINK_ADDRA_13[6]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[6]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_3, E => un1_SM_BANK_SEL_2, Q => 
        \ELINK_ADDRA_13[6]_net_1\);
    
    \ELINKS_STOP_ADDR_T[3]\ : DFN1E1C0
      port map(D => \RD_USB_ADBUS[3]_net_1\, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_7, E => 
        N_ELINKS_STOP_ADDR_T_0_sqmuxa, Q => 
        \ELINKS_STOP_ADDR_T[3]_net_1\);
    
    \ELINK_DINA_17[7]\ : DFN1E0C0
      port map(D => \N_TFC_DINA[7]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_19, E => N_197, Q => 
        \ELINK_DINA_17[7]_net_1\);
    
    \ELINK_ADDRA_11[7]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[7]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_2, E => un1_SM_BANK_SEL_16, Q => 
        \ELINK_ADDRA_11[7]_net_1\);
    
    \WR_USB_ADBUS_RNO_32[1]\ : NOR2B
      port map(A => \WR_XFER_TYPE[1]_net_1\, B => N_398, Y => 
        \WR_XFER_TYPE_m[1]\);
    
    \ELINK_BLKA[16]\ : DFN1E0P0
      port map(D => \N_ELINK_BLKA_0_iv[16]\, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_20, E => \SM_BANK_SEL[20]_net_1\, Q
         => \ELINK_BLKA[16]_net_1\);
    
    \ELINK_ADDRA_3[7]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[7]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_1_0, E => un1_SM_BANK_SEL_4, Q => 
        \ELINK_ADDRA_3[7]_net_1\);
    
    \REG_STATE_ns_i_8_tz_0[4]\ : OR2
      port map(A => \REG_STATE_ns_i_a4_2_0[4]\, B => 
        \REG_STATE_ns_i_a4_5_1[4]\, Y => 
        \REG_STATE_ns_i_8_tz_0[4]_net_1\);
    
    \ELINK_DINA_1[7]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[7]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_7, E => un1_SM_BANK_SEL_19, Q => 
        \ELINK_DINA_1[7]_net_1\);
    
    \WR_XFER_TYPE_RNO_2[0]\ : OA1C
      port map(A => N_1736, B => N_1702, C => 
        \WR_XFER_TYPE[0]_net_1\, Y => N_1817);
    
    \WR_USB_ADBUS_RNO_33[0]\ : NOR2A
      port map(A => \ELINKS_STRT_ADDR[0]_net_1\, B => N_1499, Y
         => \ELINKS_STRT_ADDR_m[0]\);
    
    \WR_USB_ADBUS_RNO_5[2]\ : AO1
      port map(A => \ELINK_DOUTA_2[2]\, B => un1_SM_BANK_SEL_32, 
        C => \ELINK_DOUTA_18_m[2]\, Y => 
        \N_WR_USB_ADBUS_0_iv_16[2]\);
    
    \WR_USB_ADBUS_RNO_13[6]\ : NOR2B
      port map(A => \ELINK_DOUTA_16[6]\, B => un1_SM_BANK_SEL_39, 
        Y => \ELINK_DOUTA_16_m[6]\);
    
    \ELINK_DINA_1[6]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[6]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_7, E => un1_SM_BANK_SEL_19, Q => 
        \ELINK_DINA_1[6]_net_1\);
    
    \WR_USB_ADBUS_RNO_32[6]\ : NOR2A
      port map(A => \ELINKS_STRT_ADDR[6]_net_1\, B => N_1499, Y
         => \ELINKS_STRT_ADDR_m[6]\);
    
    \ELINK_ADDRA_6[3]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[3]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_4, E => un1_SM_BANK_SEL_10, Q => 
        \ELINK_ADDRA_6[3]_net_1\);
    
    \WR_USB_ADBUS_RNO_22[7]\ : AO1
      port map(A => \ELINK_DOUTA_15[7]\, B => un1_SM_BANK_SEL_24, 
        C => \ELINK_DOUTA_0_m[7]\, Y => 
        \N_WR_USB_ADBUS_0_iv_8[7]\);
    
    \ELINK_ADDRA_3[4]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[4]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_1, E => un1_SM_BANK_SEL_4, Q => 
        \ELINK_ADDRA_3[4]_net_1\);
    
    \TFC_ADDRA[5]\ : DFN1E0C0
      port map(D => \N_TFC_ADDRA[5]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_10, E => N_142, Q => 
        \TFC_ADDRA[5]_net_1\);
    
    \REG_STATE_0_RNIBSOBC[2]\ : OR3
      port map(A => \REG_STATE_ns_i_i_o2_10_3[2]\, B => 
        \REG_STATE_ns_i_i_o2_10_2[2]\, C => N_349, Y => 
        \REG_STATE_ns_i_i_o2_10_5[2]\);
    
    \REG_ADDR_RNIG0CL[6]\ : NOR3
      port map(A => \REG_ADDR[6]_net_1\, B => \REG_ADDR[7]_net_1\, 
        C => \USB_TXE_B\, Y => REG_STATE_tr73_6);
    
    \TFC_DINA[6]\ : DFN1E0C0
      port map(D => \N_TFC_DINA[6]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_4, E => N_142, Q => \TFC_DINA[6]_net_1\);
    
    \ELINK_ADDRA_2[6]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[6]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_21, E => un1_SM_BANK_SEL_5, Q => 
        \ELINK_ADDRA_2[6]_net_1\);
    
    \ELINK_RWA_RNO[12]\ : AOI1
      port map(A => \SM_BANK_SEL[7]_net_1\, B => un1_USB_RXF_B_m, 
        C => \ELINK_RWA_i_m[12]\, Y => \N_ELINK_RWA_0_iv[12]\);
    
    \WR_USB_ADBUS_RNO_34[7]\ : NOR3B
      port map(A => N_1352_1, B => \OP_MODE[7]_net_1\, C => 
        REG_STATE_s20_i_0, Y => \OP_MODE_m[7]\);
    
    \REG_STATE_RNITEQN[0]\ : OR2A
      port map(A => \REG_STATE[0]_net_1\, B => 
        \REG_STATE[1]_net_1\, Y => N_1739);
    
    \WR_USB_ADBUS_RNO_25[3]\ : NOR2B
      port map(A => \ELINK_DOUTA_11[3]\, B => un1_SM_BANK_SEL_26, 
        Y => \ELINK_DOUTA_11_m[3]\);
    
    \REG_STATE_0_RNIFLMOT[5]\ : OA1
      port map(A => \REG_STATE_ns_i_a4_0_0[3]\, B => N_1259_tz, C
         => N_2592, Y => \REG_STATE_ns_i_1_0[3]\);
    
    \REG_STATE_0[1]\ : DFN1C0
      port map(D => \USB_TXE_B_RNI75TNL2\, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_22_0, Q => \REG_STATE_0[1]_net_1\);
    
    \ELINK_ADDRA_14[2]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[2]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_5, E => un1_SM_BANK_SEL_1, Q => 
        \ELINK_ADDRA_14[2]_net_1\);
    
    \ELINK_DINA_7[2]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[2]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_17, E => un1_SM_BANK_SEL_12, Q => 
        \ELINK_DINA_7[2]_net_1\);
    
    USB_RXF_B_RNIDHQ11 : NOR2A
      port map(A => N_1352_4, B => \USB_RXF_B\, Y => N_385_1);
    
    \REG_STATE_0_RNIFI3A1[1]\ : AO1B
      port map(A => \REG_STATE_0[1]_net_1\, B => 
        \REG_STATE_0[2]_net_1\, C => \REG_STATE_0[5]_net_1\, Y
         => N_1566_i_i_0);
    
    \TFC_ADDRA[0]\ : DFN1E0C0
      port map(D => \N_TFC_ADDRA[0]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_9, E => N_142, Q => 
        \TFC_ADDRA[0]_net_1\);
    
    \REG_STATE_0_RNI1R5C2[2]\ : NOR3C
      port map(A => N_TFC_STRT_ADDR_T_0_sqmuxa_0_a2_0, B => 
        \REG_STATE_0[2]_net_1\, C => N_470, Y => 
        N_TFC_STRT_ADDR_T_0_sqmuxa);
    
    \WR_USB_ADBUS_RNO_36[5]\ : NOR2B
      port map(A => \ELINK_DOUTA_0[5]\, B => un1_SM_BANK_SEL_31, 
        Y => \ELINK_DOUTA_0_m[5]\);
    
    \REG_STATE_RNITEQN_0[0]\ : NOR2B
      port map(A => \REG_STATE[0]_net_1\, B => 
        \REG_STATE[1]_net_1\, Y => N_1359_1);
    
    USB_TRIEN_B : DFI1E1P0
      port map(D => N_675_0, CLK => CLK60MHZ, E => 
        un1_REG_STATE_23, PRE => P_USB_MASTER_EN_c_16, QN => 
        TrienAux);
    
    \WR_USB_ADBUS_RNO_28[2]\ : NOR2B
      port map(A => \ELINK_DOUTA_13[2]\, B => un1_SM_BANK_SEL_29, 
        Y => \ELINK_DOUTA_13_m[2]\);
    
    U111_PATT_ELINK_BLK : DPRT_512X9_SRAM_11
      port map(ELINK_RWA_0 => \ELINK_RWA[11]_net_1\, 
        ELK_RX_SER_WORD_11(7) => ELK_RX_SER_WORD_11(7), 
        ELK_RX_SER_WORD_11(6) => ELK_RX_SER_WORD_11(6), 
        ELK_RX_SER_WORD_11(5) => ELK_RX_SER_WORD_11(5), 
        ELK_RX_SER_WORD_11(4) => ELK_RX_SER_WORD_11(4), 
        ELK_RX_SER_WORD_11(3) => ELK_RX_SER_WORD_11(3), 
        ELK_RX_SER_WORD_11(2) => ELK_RX_SER_WORD_11(2), 
        ELK_RX_SER_WORD_11(1) => ELK_RX_SER_WORD_11(1), 
        ELK_RX_SER_WORD_11(0) => ELK_RX_SER_WORD_11(0), 
        ELINK_DINA_11(7) => \ELINK_DINA_11[7]_net_1\, 
        ELINK_DINA_11(6) => \ELINK_DINA_11[6]_net_1\, 
        ELINK_DINA_11(5) => \ELINK_DINA_11[5]_net_1\, 
        ELINK_DINA_11(4) => \ELINK_DINA_11[4]_net_1\, 
        ELINK_DINA_11(3) => \ELINK_DINA_11[3]_net_1\, 
        ELINK_DINA_11(2) => \ELINK_DINA_11[2]_net_1\, 
        ELINK_DINA_11(1) => \ELINK_DINA_11[1]_net_1\, 
        ELINK_DINA_11(0) => \ELINK_DINA_11[0]_net_1\, 
        ELINK_BLKA_0 => \ELINK_BLKA[11]_net_1\, ELKS_ADDRB_0_d0
         => ELKS_ADDRB(0), ELKS_ADDRB_1 => ELKS_ADDRB(1), 
        ELKS_ADDRB_3 => ELKS_ADDRB(3), ELKS_ADDRB_5 => 
        ELKS_ADDRB(5), ELKS_ADDRB_7 => ELKS_ADDRB(7), 
        ELKS_ADDRB_0_0 => ELKS_ADDRB_0_0, ELKS_ADDRB_0_2 => 
        ELKS_ADDRB_0_2, ELKS_ADDRB_0_4 => ELKS_ADDRB_0_4, 
        ELINK_ADDRA_11(7) => \ELINK_ADDRA_11[7]_net_1\, 
        ELINK_ADDRA_11(6) => \ELINK_ADDRA_11[6]_net_1\, 
        ELINK_ADDRA_11(5) => \ELINK_ADDRA_11[5]_net_1\, 
        ELINK_ADDRA_11(4) => \ELINK_ADDRA_11[4]_net_1\, 
        ELINK_ADDRA_11(3) => \ELINK_ADDRA_11[3]_net_1\, 
        ELINK_ADDRA_11(2) => \ELINK_ADDRA_11[2]_net_1\, 
        ELINK_ADDRA_11(1) => \ELINK_ADDRA_11[1]_net_1\, 
        ELINK_ADDRA_11(0) => \ELINK_ADDRA_11[0]_net_1\, 
        PATT_ELK_DAT_11(7) => PATT_ELK_DAT_11(7), 
        PATT_ELK_DAT_11(6) => PATT_ELK_DAT_11(6), 
        PATT_ELK_DAT_11(5) => PATT_ELK_DAT_11(5), 
        PATT_ELK_DAT_11(4) => PATT_ELK_DAT_11(4), 
        PATT_ELK_DAT_11(3) => PATT_ELK_DAT_11(3), 
        PATT_ELK_DAT_11(2) => PATT_ELK_DAT_11(2), 
        PATT_ELK_DAT_11(1) => PATT_ELK_DAT_11(1), 
        PATT_ELK_DAT_11(0) => PATT_ELK_DAT_11(0), 
        ELINK_DOUTA_11(7) => \ELINK_DOUTA_11[7]\, 
        ELINK_DOUTA_11(6) => \ELINK_DOUTA_11[6]\, 
        ELINK_DOUTA_11(5) => \ELINK_DOUTA_11[5]\, 
        ELINK_DOUTA_11(4) => \ELINK_DOUTA_11[4]\, 
        ELINK_DOUTA_11(3) => \ELINK_DOUTA_11[3]\, 
        ELINK_DOUTA_11(2) => \ELINK_DOUTA_11[2]\, 
        ELINK_DOUTA_11(1) => \ELINK_DOUTA_11[1]\, 
        ELINK_DOUTA_11(0) => \ELINK_DOUTA_11[0]\, ELKS_RWB => 
        ELKS_RWB, P_USB_MASTER_EN_c_0 => P_USB_MASTER_EN_c_0, 
        CLK_40M_GL => CLK_40M_GL, CLK60MHZ => CLK60MHZ, 
        ELKS_RAM_BLKB_EN => ELKS_RAM_BLKB_EN);
    
    \TFC_ADDRA[1]\ : DFN1E0C0
      port map(D => \N_TFC_ADDRA[1]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_9, E => N_142, Q => 
        \TFC_ADDRA[1]_net_1\);
    
    \SM_BANK_SEL_RNO[14]\ : NOR3C
      port map(A => N_1882, B => N_1359_6, C => N_1351_4, Y => 
        N_1841);
    
    \REG_STATE_RNI5NQN[5]\ : OR2A
      port map(A => \REG_STATE[4]_net_1\, B => 
        \REG_STATE[5]_net_1\, Y => N_252);
    
    \ELINKS_STRT_ADDR_T[0]\ : DFN1E1C0
      port map(D => \RD_USB_ADBUS[0]_net_1\, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_21, E => 
        N_ELINKS_STRT_ADDR_T_0_sqmuxa, Q => 
        \ELINKS_STRT_ADDR_T[0]_net_1\);
    
    \WR_USB_ADBUS_RNO_23[5]\ : NOR2B
      port map(A => \ELINK_DOUTA_9[5]\, B => un1_SM_BANK_SEL_42, 
        Y => \ELINK_DOUTA_9_m[5]\);
    
    \REG_STATE_RNI0DIR1_0[4]\ : NOR2A
      port map(A => N_1710_i_0, B => N_1691, Y => N_675_0);
    
    USB_RXF_B_RNIGJ4U1 : OR2A
      port map(A => N_1351_8, B => \USB_RXF_B\, Y => N_285);
    
    \RD_USB_ADBUS_RNIGN0T[4]\ : NOR2
      port map(A => N_1700, B => \RD_USB_ADBUS[4]_net_1\, Y => 
        N_1903);
    
    \SI_CNT[3]\ : DFN1E1C0
      port map(D => SI_CNT_n3, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_5, E => SI_CNTe, Q => \SI_CNT[3]_net_1\);
    
    \ELINK_RWA[12]\ : DFN1E0P0
      port map(D => \N_ELINK_RWA_0_iv[12]\, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_11, E => \SM_BANK_SEL_0[20]_net_1\, 
        Q => \ELINK_RWA[12]_net_1\);
    
    \ELINK_ADDRA_6[2]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[2]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_4, E => un1_SM_BANK_SEL_10, Q => 
        \ELINK_ADDRA_6[2]_net_1\);
    
    \REG_STATE_0_RNI28RP1[1]\ : OA1
      port map(A => \REG_STATE_0[3]_net_1\, B => N_2617, C => 
        \REG_STATE_0[1]_net_1\, Y => N_2577);
    
    \WR_USB_ADBUS_RNO_23[3]\ : NOR2B
      port map(A => \ELINK_DOUTA_9[3]\, B => un1_SM_BANK_SEL_42, 
        Y => \ELINK_DOUTA_9_m[3]\);
    
    U116_PATT_ELINK_BLK : DPRT_512X9_SRAM_16
      port map(ELINK_RWA_0 => \ELINK_RWA[16]_net_1\, 
        ELK_RX_SER_WORD_16(7) => ELK_RX_SER_WORD_16(7), 
        ELK_RX_SER_WORD_16(6) => ELK_RX_SER_WORD_16(6), 
        ELK_RX_SER_WORD_16(5) => ELK_RX_SER_WORD_16(5), 
        ELK_RX_SER_WORD_16(4) => ELK_RX_SER_WORD_16(4), 
        ELK_RX_SER_WORD_16(3) => ELK_RX_SER_WORD_16(3), 
        ELK_RX_SER_WORD_16(2) => ELK_RX_SER_WORD_16(2), 
        ELK_RX_SER_WORD_16(1) => ELK_RX_SER_WORD_16(1), 
        ELK_RX_SER_WORD_16(0) => ELK_RX_SER_WORD_16(0), 
        ELINK_DINA_16(7) => \ELINK_DINA_16[7]_net_1\, 
        ELINK_DINA_16(6) => \ELINK_DINA_16[6]_net_1\, 
        ELINK_DINA_16(5) => \ELINK_DINA_16[5]_net_1\, 
        ELINK_DINA_16(4) => \ELINK_DINA_16[4]_net_1\, 
        ELINK_DINA_16(3) => \ELINK_DINA_16[3]_net_1\, 
        ELINK_DINA_16(2) => \ELINK_DINA_16[2]_net_1\, 
        ELINK_DINA_16(1) => \ELINK_DINA_16[1]_net_1\, 
        ELINK_DINA_16(0) => \ELINK_DINA_16[0]_net_1\, 
        ELINK_BLKA_0 => \ELINK_BLKA[16]_net_1\, ELKS_ADDRB_0_d0
         => ELKS_ADDRB(0), ELKS_ADDRB_1 => ELKS_ADDRB(1), 
        ELKS_ADDRB_3 => ELKS_ADDRB(3), ELKS_ADDRB_5 => 
        ELKS_ADDRB(5), ELKS_ADDRB_7 => ELKS_ADDRB(7), 
        ELKS_ADDRB_0_0 => ELKS_ADDRB_0_0, ELKS_ADDRB_0_2 => 
        ELKS_ADDRB_0_2, ELKS_ADDRB_0_4 => ELKS_ADDRB_0_4, 
        ELINK_ADDRA_16(7) => \ELINK_ADDRA_16[7]_net_1\, 
        ELINK_ADDRA_16(6) => \ELINK_ADDRA_16[6]_net_1\, 
        ELINK_ADDRA_16(5) => \ELINK_ADDRA_16[5]_net_1\, 
        ELINK_ADDRA_16(4) => \ELINK_ADDRA_16[4]_net_1\, 
        ELINK_ADDRA_16(3) => \ELINK_ADDRA_16[3]_net_1\, 
        ELINK_ADDRA_16(2) => \ELINK_ADDRA_16[2]_net_1\, 
        ELINK_ADDRA_16(1) => \ELINK_ADDRA_16[1]_net_1\, 
        ELINK_ADDRA_16(0) => \ELINK_ADDRA_16[0]_net_1\, 
        PATT_ELK_DAT_16(7) => PATT_ELK_DAT_16(7), 
        PATT_ELK_DAT_16(6) => PATT_ELK_DAT_16(6), 
        PATT_ELK_DAT_16(5) => PATT_ELK_DAT_16(5), 
        PATT_ELK_DAT_16(4) => PATT_ELK_DAT_16(4), 
        PATT_ELK_DAT_16(3) => PATT_ELK_DAT_16(3), 
        PATT_ELK_DAT_16(2) => PATT_ELK_DAT_16(2), 
        PATT_ELK_DAT_16(1) => PATT_ELK_DAT_16(1), 
        PATT_ELK_DAT_16(0) => PATT_ELK_DAT_16(0), 
        ELINK_DOUTA_16(7) => \ELINK_DOUTA_16[7]\, 
        ELINK_DOUTA_16(6) => \ELINK_DOUTA_16[6]\, 
        ELINK_DOUTA_16(5) => \ELINK_DOUTA_16[5]\, 
        ELINK_DOUTA_16(4) => \ELINK_DOUTA_16[4]\, 
        ELINK_DOUTA_16(3) => \ELINK_DOUTA_16[3]\, 
        ELINK_DOUTA_16(2) => \ELINK_DOUTA_16[2]\, 
        ELINK_DOUTA_16(1) => \ELINK_DOUTA_16[1]\, 
        ELINK_DOUTA_16(0) => \ELINK_DOUTA_16[0]\, ELKS_RWB => 
        ELKS_RWB, P_USB_MASTER_EN_c_0 => P_USB_MASTER_EN_c_0, 
        CLK_40M_GL => CLK_40M_GL, CLK60MHZ => CLK60MHZ, 
        ELKS_RAM_BLKB_EN => ELKS_RAM_BLKB_EN);
    
    \TFC_STRT_ADDR[5]\ : DFN1E1C0
      port map(D => \TFC_STRT_ADDR_T[5]_net_1\, CLK => CLK60MHZ, 
        CLR => P_USB_MASTER_EN_c_13, E => \REG_STATE_d_0[30]\, Q
         => \TFC_STRT_ADDR[5]_net_1\);
    
    \REG_STATE_RNIVU1F2[2]\ : NOR2B
      port map(A => N_1782_1, B => N_1907, Y => 
        N_TFC_STOP_ADDR_T_0_sqmuxa);
    
    \ELINK_ADDRA_17[1]\ : DFN1E0C0
      port map(D => \N_TFC_ADDRA[1]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_10, E => N_197, Q => 
        \ELINK_ADDRA_17[1]_net_1\);
    
    \WR_USB_ADBUS_RNO_9[7]\ : AO1
      port map(A => \ELINK_DOUTA_7[7]\, B => un1_SM_BANK_SEL_37, 
        C => \ELINK_DOUTA_9_m[7]\, Y => 
        \N_WR_USB_ADBUS_0_iv_14[7]\);
    
    \ELINK_RWA[0]\ : DFN1E0P0
      port map(D => \N_ELINK_RWA_0_iv[0]\, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_6, E => \SM_BANK_SEL_0[20]_net_1\, 
        Q => \ELINK_RWA[0]_net_1\);
    
    \ELINK_RWA_RNO_0[18]\ : OA1B
      port map(A => N_624_15, B => \N_ELINK_RWA_0_iv_0_o2_0[18]\, 
        C => \ELINK_RWA[18]_net_1\, Y => N_171);
    
    USB_RD_BI_RNO : NOR3
      port map(A => N_USB_RD_BI_i_5, B => N_1867, C => N_1866, Y
         => N_1673);
    
    \REG_ADDR_RNIKPCP[1]\ : NOR3B
      port map(A => N_261, B => \REG_ADDR[1]_net_1\, C => 
        \SM_BANK_SEL_0[21]_net_1\, Y => \N_TFC_ADDRA[1]\);
    
    \WR_USB_ADBUS_RNO_4[1]\ : AO1
      port map(A => \ELINK_DOUTA_16[1]\, B => un1_SM_BANK_SEL_39, 
        C => \ELINK_DOUTA_1_m[1]\, Y => 
        \N_WR_USB_ADBUS_0_iv_9[1]\);
    
    U4C_REGCROSS : CLK60M_TO_40M_4_1
      port map(ELINKS_STRT_ADDR(7) => \ELINKS_STRT_ADDR[7]_net_1\, 
        ELINKS_STRT_ADDR(6) => \ELINKS_STRT_ADDR[6]_net_1\, 
        ELINKS_STRT_ADDR(5) => \ELINKS_STRT_ADDR[5]_net_1\, 
        ELINKS_STRT_ADDR(4) => \ELINKS_STRT_ADDR[4]_net_1\, 
        ELINKS_STRT_ADDR(3) => \ELINKS_STRT_ADDR[3]_net_1\, 
        ELINKS_STRT_ADDR(2) => \ELINKS_STRT_ADDR[2]_net_1\, 
        ELINKS_STRT_ADDR(1) => \ELINKS_STRT_ADDR[1]_net_1\, 
        ELINKS_STRT_ADDR(0) => \ELINKS_STRT_ADDR[0]_net_1\, 
        ELKS_STRT_ADDR(7) => ELKS_STRT_ADDR(7), ELKS_STRT_ADDR(6)
         => ELKS_STRT_ADDR(6), ELKS_STRT_ADDR(5) => 
        ELKS_STRT_ADDR(5), ELKS_STRT_ADDR(4) => ELKS_STRT_ADDR(4), 
        ELKS_STRT_ADDR(3) => ELKS_STRT_ADDR(3), ELKS_STRT_ADDR(2)
         => ELKS_STRT_ADDR(2), ELKS_STRT_ADDR(1) => 
        ELKS_STRT_ADDR(1), ELKS_STRT_ADDR(0) => ELKS_STRT_ADDR(0), 
        P_MASTER_POR_B_c_28 => P_MASTER_POR_B_c_28, 
        P_MASTER_POR_B_c_22_0 => P_MASTER_POR_B_c_22_0, 
        P_MASTER_POR_B_c_33 => P_MASTER_POR_B_c_33, 
        P_MASTER_POR_B_c_21 => P_MASTER_POR_B_c_21, 
        P_MASTER_POR_B_c_32 => P_MASTER_POR_B_c_32, CLK_40M_GL
         => CLK_40M_GL);
    
    \ELINK_ADDRA_16[6]\ : DFN1E0C0
      port map(D => \N_TFC_ADDRA[6]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_9, E => N_200, Q => 
        \ELINK_ADDRA_16[6]_net_1\);
    
    \SM_BANK_SEL_RNI49E6[12]\ : OR2
      port map(A => \N_ELINK_RWA_15_1[8]\, B => N_620_10, Y => 
        N_624_15);
    
    \RD_XFER_TYPE_RNO[1]\ : AO1
      port map(A => \RD_XFER_TYPE[1]_net_1\, B => N_1703, C => 
        N_1796, Y => \RD_XFER_TYPE_RNO[1]_net_1\);
    
    \ELINK_ADDRA_3[6]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[6]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_1, E => un1_SM_BANK_SEL_4, Q => 
        \ELINK_ADDRA_3[6]_net_1\);
    
    \REG_STATE_RNI3LQN_0[3]\ : OR2A
      port map(A => \REG_STATE[3]_net_1\, B => 
        \REG_STATE[4]_net_1\, Y => N_292);
    
    \REG_ADDR[2]\ : DFN1E1C0
      port map(D => N_2629, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_10, E => REG_ADDRe, Q => 
        \REG_ADDR[2]_net_1\);
    
    \ELINK_ADDRA_5[5]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[5]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_3, E => un1_SM_BANK_SEL_15, Q => 
        \ELINK_ADDRA_5[5]_net_1\);
    
    \ELINK_DINA_8[0]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[0]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_18, E => un1_SM_BANK_SEL_21, Q => 
        \ELINK_DINA_8[0]_net_1\);
    
    \ELINK_DINA_5[0]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[0]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_14, E => un1_SM_BANK_SEL_15, Q => 
        \ELINK_DINA_5[0]_net_1\);
    
    \ELINKS_STOP_ADDR[1]\ : DFN1E1C0
      port map(D => \ELINKS_STOP_ADDR_T[1]_net_1\, CLK => 
        CLK60MHZ, CLR => P_USB_MASTER_EN_c_14, E => 
        \REG_STATE_d_0[30]\, Q => \ELINKS_STOP_ADDR[1]_net_1\);
    
    \ELINK_RWA[19]\ : DFN1E0P0
      port map(D => \N_ELINK_RWA_0_iv[19]\, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_12, E => \SM_BANK_SEL_0[20]_net_1\, 
        Q => \ELINK_RWA[19]_net_1\);
    
    \ELINK_DINA_16[5]\ : DFN1E0C0
      port map(D => \N_TFC_DINA[5]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_18, E => N_200, Q => 
        \ELINK_DINA_16[5]_net_1\);
    
    \ELINK_ADDRA_5[1]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[1]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_3, E => un1_SM_BANK_SEL_15, Q => 
        \ELINK_ADDRA_5[1]_net_1\);
    
    \ELINKS_STOP_ADDR[7]\ : DFN1E1C0
      port map(D => \ELINKS_STOP_ADDR_T[7]_net_1\, CLK => 
        CLK60MHZ, CLR => P_USB_MASTER_EN_c_14, E => 
        \REG_STATE_d[30]\, Q => \ELINKS_STOP_ADDR[7]_net_1\);
    
    \ELINK_ADDRA_13[4]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[4]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_3, E => un1_SM_BANK_SEL_2, Q => 
        \ELINK_ADDRA_13[4]_net_1\);
    
    \ELINK_DINA_7[3]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[3]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_17, E => un1_SM_BANK_SEL_12, Q => 
        \ELINK_DINA_7[3]_net_1\);
    
    \SM_BANK_SEL_RNI3TN22[16]\ : NOR3A
      port map(A => \SM_BANK_SEL[16]_net_1\, B => N_312, C => 
        N_1566_i_i_0, Y => un1_SM_BANK_SEL_43);
    
    \REG_STATE_ns_i_a4_1_0[4]\ : NOR2A
      port map(A => N_2606, B => N_379, Y => 
        \REG_STATE_ns_i_a4_1_0[4]_net_1\);
    
    \ELINK_DINA_15[4]\ : DFN1E0C0
      port map(D => \N_TFC_DINA[4]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_16, E => N_199, Q => 
        \ELINK_DINA_15[4]_net_1\);
    
    \REG_ADDR_RNIL0HE[5]\ : NOR2
      port map(A => \REG_ADDR[0]_net_1\, B => \REG_ADDR[5]_net_1\, 
        Y => REG_STATE_tr73_1);
    
    ELK_N_ACTIVE_RNIGJ8H3 : AO1A
      port map(A => N_273, B => N_262_i, C => \ELK_N_ACTIVE\, Y
         => N_277);
    
    \ELINK_BLKA[12]\ : DFN1E0P0
      port map(D => \N_ELINK_BLKA_0_iv[12]\, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_20, E => \SM_BANK_SEL[20]_net_1\, Q
         => \ELINK_BLKA[12]_net_1\);
    
    \ELINK_ADDRA_6[5]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[5]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_4, E => un1_SM_BANK_SEL_10, Q => 
        \ELINK_ADDRA_6[5]_net_1\);
    
    \ELINK_ADDRA_5[0]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[0]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_3, E => un1_SM_BANK_SEL_15, Q => 
        \ELINK_ADDRA_5[0]_net_1\);
    
    \ELINK_ADDRA_4[4]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[4]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_2_0, E => un1_SM_BANK_SEL_8, Q => 
        \ELINK_ADDRA_4[4]_net_1\);
    
    \SM_BANK_SEL_RNIF01C2[5]\ : NOR3A
      port map(A => \SM_BANK_SEL[5]_net_1\, B => N_312_0, C => 
        N_1566_i_i_0, Y => un1_SM_BANK_SEL_23);
    
    USB_RXF_B_0 : DFN1P0
      port map(D => P_USB_RXF_B_c, CLK => CLK60MHZ, PRE => 
        P_USB_MASTER_EN_c, Q => \USB_RXF_B_0\);
    
    \ELINK_ADDRA_7[4]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[4]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_6, E => un1_SM_BANK_SEL_12, Q => 
        \ELINK_ADDRA_7[4]_net_1\);
    
    \WR_XFER_TYPE_RNO_0[2]\ : NOR2
      port map(A => N_1716, B => \RD_USB_ADBUS[2]_net_1\, Y => 
        N_1824);
    
    \ELINK_RWA_RNO[15]\ : AOI1
      port map(A => \SM_BANK_SEL[4]_net_1\, B => un1_USB_RXF_B_m, 
        C => N_175, Y => \N_ELINK_RWA_0_iv[15]\);
    
    \ELINK_DINA_14[5]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[5]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_16, E => un1_SM_BANK_SEL_1, Q => 
        \ELINK_DINA_14[5]_net_1\);
    
    \WR_USB_ADBUS_RNO_2[1]\ : OR3
      port map(A => \N_WR_USB_ADBUS_0_iv_14[1]\, B => 
        \N_WR_USB_ADBUS_0_iv_13[1]\, C => 
        \N_WR_USB_ADBUS_0_iv_22[1]\, Y => 
        \N_WR_USB_ADBUS_0_iv_25[1]\);
    
    \RD_USB_ADBUS[4]\ : DFN1C0
      port map(D => \N_RD_USB_ADBUS[4]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_22, Q => \RD_USB_ADBUS[4]_net_1\);
    
    \RD_XFER_TYPE_RNIRON38[0]\ : NOR3B
      port map(A => N_480, B => N_1370_i_i_a5_0, C => N_273, Y
         => N_359);
    
    \WR_USB_ADBUS_RNO_1[7]\ : OR3
      port map(A => \N_WR_USB_ADBUS_0_iv_6[7]\, B => 
        \ELINK_DOUTA_14_m[7]\, C => \N_WR_USB_ADBUS_0_iv_18[7]\, 
        Y => \N_WR_USB_ADBUS_0_iv_23[7]\);
    
    \SM_BANK_SEL_RNIP0VN[18]\ : OR3A
      port map(A => N_143, B => N_616_11, C => \N_ELINK_RWA_1[0]\, 
        Y => \N_ELINK_RWA_3[0]\);
    
    \REG_ADDR_RNIP4HE[3]\ : NOR2B
      port map(A => \REG_ADDR[6]_net_1\, B => \REG_ADDR[3]_net_1\, 
        Y => N_1398_i_0_a2_1);
    
    \ELINK_BLKA[9]\ : DFN1E0P0
      port map(D => \N_ELINK_BLKA_0_iv[9]\, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_19, E => \SM_BANK_SEL[20]_net_1\, Q
         => \ELINK_BLKA[9]_net_1\);
    
    \RD_USB_ADBUS_RNIMT0T[6]\ : OR2
      port map(A => N_293, B => \RD_USB_ADBUS[6]_net_1\, Y => 
        N_1729);
    
    \ELINK_BLKA_RNO_0[11]\ : NOR2B
      port map(A => \SM_BANK_SEL[8]_net_1\, B => X_BLKA_i, Y => 
        N_162);
    
    \WR_USB_ADBUS_RNO_22[5]\ : AO1
      port map(A => \ELINK_DOUTA_15[5]\, B => un1_SM_BANK_SEL_24, 
        C => \ELINK_DOUTA_0_m[5]\, Y => 
        \N_WR_USB_ADBUS_0_iv_8[5]\);
    
    \REG_STATE_ns_i_i_a2_0_2_RNO_0[0]\ : NOR3A
      port map(A => \USB_RXF_B_0\, B => N_413, C => N_412, Y => 
        \REG_STATE_ns_i_i_a2_0_1[0]\);
    
    \ELINK_ADDRA_18[3]\ : DFN1E0C0
      port map(D => \N_TFC_ADDRA[3]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_12, E => N_198, Q => 
        \ELINK_ADDRA_18[3]_net_1\);
    
    \WR_USB_ADBUS_RNO_0[0]\ : OR3
      port map(A => \N_WR_USB_ADBUS_0_iv_10[0]\, B => 
        \N_WR_USB_ADBUS_0_iv_9[0]\, C => 
        \N_WR_USB_ADBUS_0_iv_20[0]\, Y => 
        \N_WR_USB_ADBUS_0_iv_24[0]\);
    
    \RD_USB_ADBUS_RNIRFIK2[6]\ : NOR2A
      port map(A => \RD_USB_ADBUS[6]_net_1\, B => N_206, Y => 
        \N_TFC_DINA[6]\);
    
    USB_TXE_B_RNIU9JI6 : AO1
      port map(A => \USB_TXE_B\, B => N_2520, C => 
        \REG_STATE_ns_i_tz_1[5]\, Y => N_2454_tz);
    
    \WR_USB_ADBUS_RNO_26[1]\ : NOR2B
      port map(A => \ELINK_DOUTA_10[1]\, B => un1_SM_BANK_SEL_34, 
        Y => \ELINK_DOUTA_10_m[1]\);
    
    \ELINK_ADDRA_12[5]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[5]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_2_0, E => un1_SM_BANK_SEL_7, Q => 
        \ELINK_ADDRA_12[5]_net_1\);
    
    \ELINK_ADDRA_2[3]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[3]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_21, E => un1_SM_BANK_SEL_5, Q => 
        \ELINK_ADDRA_2[3]_net_1\);
    
    \REG_STATE_0_RNITKSV81[5]\ : AO1
      port map(A => N_510, B => N_1398_i_0_0, C => N_311, Y => 
        N_513);
    
    \WR_USB_ADBUS_RNO_33[1]\ : NOR2A
      port map(A => \ELINKS_STRT_ADDR[1]_net_1\, B => N_1499, Y
         => \ELINKS_STRT_ADDR_m[1]\);
    
    USB_WR_BI_RNO_0 : OA1
      port map(A => N_1352_1, B => N_1744_i, C => 
        \REG_STATE_0[4]_net_1\, Y => N_1779);
    
    \ELINK_DINA_15[2]\ : DFN1E0C0
      port map(D => \N_TFC_DINA[2]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_16, E => N_199, Q => 
        \ELINK_DINA_15[2]_net_1\);
    
    \WR_USB_ADBUS_RNO_20[2]\ : AO1
      port map(A => \ELINK_DOUTA_10[2]\, B => un1_SM_BANK_SEL_34, 
        C => \ELINK_DOUTA_11_m[2]\, Y => 
        \N_WR_USB_ADBUS_0_iv_10[2]\);
    
    \WR_USB_ADBUS_RNO_27[7]\ : AO1
      port map(A => \ELINK_DOUTA_12[7]\, B => un1_SM_BANK_SEL_33, 
        C => \ELINK_DOUTA_13_m[7]\, Y => 
        \N_WR_USB_ADBUS_0_iv_16[7]\);
    
    \TFC_STOP_ADDR[5]\ : DFN1E1C0
      port map(D => \TFC_STOP_ADDR_T[5]_net_1\, CLK => CLK60MHZ, 
        CLR => P_USB_MASTER_EN_c_8, E => \REG_STATE_d_0[30]\, Q
         => \TFC_STOP_ADDR[5]_net_1\);
    
    \TFC_DINA[0]\ : DFN1E0C0
      port map(D => \N_TFC_DINA[0]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_4, E => N_142, Q => \TFC_DINA[0]_net_1\);
    
    \ELINK_ADDRA_3[3]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[3]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_1, E => un1_SM_BANK_SEL_4, Q => 
        \ELINK_ADDRA_3[3]_net_1\);
    
    \WR_USB_ADBUS_RNO_29[3]\ : NOR3B
      port map(A => N_1730_i, B => \ELINKS_STOP_ADDR[3]_net_1\, C
         => N_1726, Y => \ELINKS_STOP_ADDR_m[3]\);
    
    \ELINK_BLKA_RNO[19]\ : OA1C
      port map(A => N_130, B => \ELINK_BLKA[19]_net_1\, C => 
        X_BLKA_i_m_18, Y => \N_ELINK_BLKA_0_iv[19]\);
    
    \SM_BANK_SEL_RNINSK6[9]\ : NOR2
      port map(A => \SM_BANK_SEL[9]_net_1\, B => 
        \SM_BANK_SEL[11]_net_1\, Y => 
        \N_ELINK_BLKA_0_iv_0_o2_i_a5_0[9]\);
    
    \WR_USB_ADBUS_RNO_29[0]\ : OR3
      port map(A => \N_WR_USB_ADBUS_0_iv_0[0]_net_1\, B => 
        \OP_MODE_m[0]\, C => \ELINKS_STRT_ADDR_m[0]\, Y => 
        \N_WR_USB_ADBUS_0_iv_2[0]\);
    
    \TFC_STOP_ADDR_T[4]\ : DFN1E1C0
      port map(D => \RD_USB_ADBUS[4]_net_1\, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_15, E => N_TFC_STOP_ADDR_T_0_sqmuxa, 
        Q => \TFC_STOP_ADDR_T[4]_net_1\);
    
    \REG_ADDR_RNIILOT[1]\ : NOR3B
      port map(A => \REG_ADDR[0]_net_1\, B => \REG_ADDR[1]_net_1\, 
        C => \USB_RXF_B_0\, Y => REG_STATE_tr49_4);
    
    \TFC_DINA[4]\ : DFN1E0C0
      port map(D => \N_TFC_DINA[4]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_4, E => N_142, Q => \TFC_DINA[4]_net_1\);
    
    \REG_STATE_0_RNIGAMT1[2]\ : NOR3A
      port map(A => N_1499_2_i_0, B => N_257, C => 
        \REG_STATE_0[2]_net_1\, Y => N_454);
    
    \REG_STATE_RNITNN31_0[2]\ : NOR2A
      port map(A => N_1352_1, B => \REG_STATE[2]_net_1\, Y => 
        N_1782_1);
    
    \REG_STATE_RNI2TN31[4]\ : OR2A
      port map(A => N_1690_i, B => \REG_STATE[4]_net_1\, Y => 
        N_1691);
    
    \RD_USB_ADBUS_RNIV3BJ_1[3]\ : NOR2A
      port map(A => \RD_USB_ADBUS[3]_net_1\, B => 
        \RD_USB_ADBUS[2]_net_1\, Y => N_1352_5);
    
    \ELINKS_STOP_ADDR[6]\ : DFN1E1C0
      port map(D => \ELINKS_STOP_ADDR_T[6]_net_1\, CLK => 
        CLK60MHZ, CLR => P_USB_MASTER_EN_c_14, E => 
        \REG_STATE_d[30]\, Q => \ELINKS_STOP_ADDR[6]_net_1\);
    
    \WR_USB_ADBUS_RNO_8[2]\ : AO1
      port map(A => \ELINK_DOUTA_0[2]\, B => un1_SM_BANK_SEL_31, 
        C => \ELINK_DOUTA_16_m[2]\, Y => 
        \N_WR_USB_ADBUS_0_iv_14[2]\);
    
    \REG_STATE_0[4]\ : DFN1C0
      port map(D => \REG_STATE_RNIMO53U3[2]_net_1\, CLK => 
        CLK60MHZ, CLR => P_USB_MASTER_EN_c_22_0, Q => 
        \REG_STATE_0[4]_net_1\);
    
    \SM_BANK_SEL_RNIU06G[0]\ : OR2
      port map(A => \SM_BANK_SEL[0]_net_1\, B => 
        \SM_BANK_SEL_0[21]_net_1\, Y => un1_SM_BANK_SEL_11);
    
    \SM_BANK_SEL[9]\ : DFN1E1C0
      port map(D => N_1847, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_8, E => un1_REG_STATE_30, Q => 
        \SM_BANK_SEL[9]_net_1\);
    
    \ELINK_DINA_3[3]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[3]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_11, E => un1_SM_BANK_SEL_4, Q => 
        \ELINK_DINA_3[3]_net_1\);
    
    U103_PATT_ELINK_BLK : DPRT_512X9_SRAM_3
      port map(ELINK_RWA_0 => \ELINK_RWA[3]_net_1\, 
        ELK_RX_SER_WORD_3(7) => ELK_RX_SER_WORD_3(7), 
        ELK_RX_SER_WORD_3(6) => ELK_RX_SER_WORD_3(6), 
        ELK_RX_SER_WORD_3(5) => ELK_RX_SER_WORD_3(5), 
        ELK_RX_SER_WORD_3(4) => ELK_RX_SER_WORD_3(4), 
        ELK_RX_SER_WORD_3(3) => ELK_RX_SER_WORD_3(3), 
        ELK_RX_SER_WORD_3(2) => ELK_RX_SER_WORD_3(2), 
        ELK_RX_SER_WORD_3(1) => ELK_RX_SER_WORD_3(1), 
        ELK_RX_SER_WORD_3(0) => ELK_RX_SER_WORD_3(0), 
        ELINK_DINA_3(7) => \ELINK_DINA_3[7]_net_1\, 
        ELINK_DINA_3(6) => \ELINK_DINA_3[6]_net_1\, 
        ELINK_DINA_3(5) => \ELINK_DINA_3[5]_net_1\, 
        ELINK_DINA_3(4) => \ELINK_DINA_3[4]_net_1\, 
        ELINK_DINA_3(3) => \ELINK_DINA_3[3]_net_1\, 
        ELINK_DINA_3(2) => \ELINK_DINA_3[2]_net_1\, 
        ELINK_DINA_3(1) => \ELINK_DINA_3[1]_net_1\, 
        ELINK_DINA_3(0) => \ELINK_DINA_3[0]_net_1\, ELINK_BLKA_0
         => \ELINK_BLKA[3]_net_1\, ELKS_ADDRB_0_d0 => 
        ELKS_ADDRB(0), ELKS_ADDRB_1 => ELKS_ADDRB(1), 
        ELKS_ADDRB_3 => ELKS_ADDRB(3), ELKS_ADDRB_5 => 
        ELKS_ADDRB(5), ELKS_ADDRB_7 => ELKS_ADDRB(7), 
        ELKS_ADDRB_0_0 => ELKS_ADDRB_0_0, ELKS_ADDRB_0_2 => 
        ELKS_ADDRB_0_2, ELKS_ADDRB_0_4 => ELKS_ADDRB_0_4, 
        ELINK_ADDRA_3(7) => \ELINK_ADDRA_3[7]_net_1\, 
        ELINK_ADDRA_3(6) => \ELINK_ADDRA_3[6]_net_1\, 
        ELINK_ADDRA_3(5) => \ELINK_ADDRA_3[5]_net_1\, 
        ELINK_ADDRA_3(4) => \ELINK_ADDRA_3[4]_net_1\, 
        ELINK_ADDRA_3(3) => \ELINK_ADDRA_3[3]_net_1\, 
        ELINK_ADDRA_3(2) => \ELINK_ADDRA_3[2]_net_1\, 
        ELINK_ADDRA_3(1) => \ELINK_ADDRA_3[1]_net_1\, 
        ELINK_ADDRA_3(0) => \ELINK_ADDRA_3[0]_net_1\, 
        PATT_ELK_DAT_3(7) => PATT_ELK_DAT_3(7), PATT_ELK_DAT_3(6)
         => PATT_ELK_DAT_3(6), PATT_ELK_DAT_3(5) => 
        PATT_ELK_DAT_3(5), PATT_ELK_DAT_3(4) => PATT_ELK_DAT_3(4), 
        PATT_ELK_DAT_3(3) => PATT_ELK_DAT_3(3), PATT_ELK_DAT_3(2)
         => PATT_ELK_DAT_3(2), PATT_ELK_DAT_3(1) => 
        PATT_ELK_DAT_3(1), PATT_ELK_DAT_3(0) => PATT_ELK_DAT_3(0), 
        ELINK_DOUTA_3(7) => \ELINK_DOUTA_3[7]\, ELINK_DOUTA_3(6)
         => \ELINK_DOUTA_3[6]\, ELINK_DOUTA_3(5) => 
        \ELINK_DOUTA_3[5]\, ELINK_DOUTA_3(4) => 
        \ELINK_DOUTA_3[4]\, ELINK_DOUTA_3(3) => 
        \ELINK_DOUTA_3[3]\, ELINK_DOUTA_3(2) => 
        \ELINK_DOUTA_3[2]\, ELINK_DOUTA_3(1) => 
        \ELINK_DOUTA_3[1]\, ELINK_DOUTA_3(0) => 
        \ELINK_DOUTA_3[0]\, ELKS_RWB => ELKS_RWB, 
        P_USB_MASTER_EN_c_0 => P_USB_MASTER_EN_c_0, CLK_40M_GL
         => CLK_40M_GL, CLK60MHZ => CLK60MHZ, ELKS_RAM_BLKB_EN
         => ELKS_RAM_BLKB_EN);
    
    \RD_USB_ADBUS_RNIDK0T[5]\ : NOR2
      port map(A => N_1352_4, B => \RD_USB_ADBUS[5]_net_1\, Y => 
        N_356);
    
    USB_RXF_B_RNIN32A2 : NOR3B
      port map(A => N_1499_2_i_0, B => \REG_STATE_ns_i_a4_3_0[4]\, 
        C => N_268, Y => N_2566);
    
    \ELINK_RWA_RNO[5]\ : AOI1
      port map(A => \SM_BANK_SEL[14]_net_1\, B => un1_USB_RXF_B_m, 
        C => N_183, Y => \N_ELINK_RWA_0_iv[5]\);
    
    \WR_USB_ADBUS_RNO_11[0]\ : OR3
      port map(A => \ELINK_DOUTA_17_m[0]\, B => 
        \ELINK_DOUTA_1_m[0]\, C => \N_WR_USB_ADBUS_0_iv_16[0]\, Y
         => \N_WR_USB_ADBUS_0_iv_22[0]\);
    
    \SM_BANK_SEL[0]\ : DFN1E1C0
      port map(D => N_1834, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_7, E => un1_REG_STATE_30, Q => 
        \SM_BANK_SEL[0]_net_1\);
    
    \WR_XFER_TYPE_RNIUDSS_0[0]\ : NOR2
      port map(A => \WR_XFER_TYPE[0]_net_1\, B => 
        \WR_XFER_TYPE[2]_net_1\, Y => REG_STATE_tr72_6_0);
    
    \REG_STATE[1]\ : DFN1C0
      port map(D => \USB_TXE_B_RNI75TNL2\, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_22_0, Q => \REG_STATE[1]_net_1\);
    
    \ELINK_ADDRA_6[4]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[4]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_4, E => un1_SM_BANK_SEL_10, Q => 
        \ELINK_ADDRA_6[4]_net_1\);
    
    \RD_USB_ADBUS[0]\ : DFN1C0
      port map(D => \N_RD_USB_ADBUS[0]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_22, Q => \RD_USB_ADBUS[0]_net_1\);
    
    \SM_BANK_SEL_RNI1CL1[21]\ : NOR2
      port map(A => \SM_BANK_SEL[21]_net_1\, B => 
        \SM_BANK_SEL[20]_net_1\, Y => N_142);
    
    \RD_XFER_TYPE_RNO_0[4]\ : NOR2A
      port map(A => \RD_USB_ADBUS[4]_net_1\, B => N_1694, Y => 
        N_1802);
    
    \WR_USB_ADBUS_RNO_0[6]\ : OR3
      port map(A => \N_WR_USB_ADBUS_0_iv_9[6]\, B => 
        \N_WR_USB_ADBUS_0_iv_8[6]\, C => 
        \N_WR_USB_ADBUS_0_iv_19[6]\, Y => 
        \N_WR_USB_ADBUS_0_iv_23[6]\);
    
    \WR_USB_ADBUS_RNO_18[1]\ : OR3
      port map(A => \OP_MODE_m[1]\, B => \TFC_STOP_ADDR_m[1]\, C
         => \WR_XFER_TYPE_m[1]\, Y => \N_WR_USB_ADBUS_0_iv_2[1]\);
    
    \WR_USB_ADBUS_RNO_25[5]\ : NOR2B
      port map(A => \ELINK_DOUTA_8[5]\, B => un1_SM_BANK_SEL_38, 
        Y => \ELINK_DOUTA_8_m[5]\);
    
    \SI_CNT_RNO[0]\ : NOR2
      port map(A => \SI_CNT[0]_net_1\, B => N_678, Y => N_2625);
    
    \SM_BANK_SEL_RNIBS0C2[1]\ : NOR3A
      port map(A => \SM_BANK_SEL[1]_net_1\, B => N_312_0, C => 
        N_1566_i_i_0, Y => un1_SM_BANK_SEL_25);
    
    \WR_USB_ADBUS_RNO_28[5]\ : AO1
      port map(A => \ELINK_DOUTA_12[5]\, B => un1_SM_BANK_SEL_33, 
        C => \ELINK_DOUTA_13_m[5]\, Y => 
        \N_WR_USB_ADBUS_0_iv_16[5]\);
    
    \WR_USB_ADBUS_RNO_26[6]\ : AO1
      port map(A => \ELINK_DOUTA_2[6]\, B => un1_SM_BANK_SEL_32, 
        C => \ELINK_DOUTA_15_m[6]\, Y => 
        \N_WR_USB_ADBUS_0_iv_15[6]\);
    
    \ELINK_BLKA_RNO[4]\ : AOI1
      port map(A => \SM_BANK_SEL[15]_net_1\, B => X_BLKA_i, C => 
        \ELINK_BLKA_i_m[4]\, Y => \N_ELINK_BLKA_0_iv[4]\);
    
    \WR_USB_ADBUS_RNO_2[6]\ : OR3
      port map(A => \N_WR_USB_ADBUS_0_iv_13[6]\, B => 
        \N_WR_USB_ADBUS_0_iv_12[6]\, C => 
        \N_WR_USB_ADBUS_0_iv_21[6]\, Y => 
        \N_WR_USB_ADBUS_0_iv_24[6]\);
    
    \ELINK_DINA_5[1]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[1]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_14, E => un1_SM_BANK_SEL_15, Q => 
        \ELINK_DINA_5[1]_net_1\);
    
    \WR_USB_ADBUS_RNO_10[3]\ : AO1
      port map(A => \ELINK_DOUTA_6[3]\, B => un1_SM_BANK_SEL_30, 
        C => \ELINK_DOUTA_8_m[3]\, Y => 
        \N_WR_USB_ADBUS_0_iv_13[3]\);
    
    \ELINK_ADDRA_5[2]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[2]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_3, E => un1_SM_BANK_SEL_15, Q => 
        \ELINK_ADDRA_5[2]_net_1\);
    
    \ELINK_ADDRA_7[3]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[3]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_6, E => un1_SM_BANK_SEL_12, Q => 
        \ELINK_ADDRA_7[3]_net_1\);
    
    \WR_XFER_TYPE_RNO_1[1]\ : NOR3A
      port map(A => \RD_USB_ADBUS[0]_net_1\, B => 
        \WR_XFER_TYPE[1]_net_1\, C => \RD_USB_ADBUS[5]_net_1\, Y
         => N_1821);
    
    \WR_USB_ADBUS_RNO_9[3]\ : AO1
      port map(A => \ELINK_DOUTA_7[3]\, B => un1_SM_BANK_SEL_37, 
        C => \ELINK_DOUTA_9_m[3]\, Y => 
        \N_WR_USB_ADBUS_0_iv_14[3]\);
    
    \OP_MODE[6]\ : DFN1E1C0
      port map(D => \OP_MODE_T[6]_net_1\, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_15, E => \REG_STATE_d[30]\, Q => 
        \OP_MODE[6]_net_1\);
    
    \N_TFC_ADDRA_0_o2_RNO_2[7]\ : AO1
      port map(A => \N_TFC_ADDRA_0_a2_6_0[7]\, B => N_1352_1, C
         => N_424, Y => N_253);
    
    USB_RD_BI_RNO_7 : NOR3B
      port map(A => N_USB_RD_BI_i_a2_4_1, B => 
        N_USB_RD_BI_i_a2_4_3, C => N_1695, Y => N_1869);
    
    \ELINK_ADDRA_5[3]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[3]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_3, E => un1_SM_BANK_SEL_15, Q => 
        \ELINK_ADDRA_5[3]_net_1\);
    
    U102_PATT_ELINK_BLK : DPRT_512X9_SRAM_2
      port map(ELINK_RWA_0 => \ELINK_RWA[2]_net_1\, 
        ELK_RX_SER_WORD_2(7) => ELK_RX_SER_WORD_2(7), 
        ELK_RX_SER_WORD_2(6) => ELK_RX_SER_WORD_2(6), 
        ELK_RX_SER_WORD_2(5) => ELK_RX_SER_WORD_2(5), 
        ELK_RX_SER_WORD_2(4) => ELK_RX_SER_WORD_2(4), 
        ELK_RX_SER_WORD_2(3) => ELK_RX_SER_WORD_2(3), 
        ELK_RX_SER_WORD_2(2) => ELK_RX_SER_WORD_2(2), 
        ELK_RX_SER_WORD_2(1) => ELK_RX_SER_WORD_2(1), 
        ELK_RX_SER_WORD_2(0) => ELK_RX_SER_WORD_2(0), 
        ELINK_DINA_2(7) => \ELINK_DINA_2[7]_net_1\, 
        ELINK_DINA_2(6) => \ELINK_DINA_2[6]_net_1\, 
        ELINK_DINA_2(5) => \ELINK_DINA_2[5]_net_1\, 
        ELINK_DINA_2(4) => \ELINK_DINA_2[4]_net_1\, 
        ELINK_DINA_2(3) => \ELINK_DINA_2[3]_net_1\, 
        ELINK_DINA_2(2) => \ELINK_DINA_2[2]_net_1\, 
        ELINK_DINA_2(1) => \ELINK_DINA_2[1]_net_1\, 
        ELINK_DINA_2(0) => \ELINK_DINA_2[0]_net_1\, ELINK_BLKA_0
         => \ELINK_BLKA[2]_net_1\, ELKS_ADDRB(7) => ELKS_ADDRB(7), 
        ELKS_ADDRB(6) => ELKS_ADDRB(6), ELKS_ADDRB(5) => 
        ELKS_ADDRB(5), ELKS_ADDRB(4) => ELKS_ADDRB(4), 
        ELKS_ADDRB(3) => ELKS_ADDRB(3), ELKS_ADDRB(2) => 
        ELKS_ADDRB(2), ELKS_ADDRB(1) => ELKS_ADDRB(1), 
        ELKS_ADDRB(0) => ELKS_ADDRB(0), ELINK_ADDRA_2(7) => 
        \ELINK_ADDRA_2[7]_net_1\, ELINK_ADDRA_2(6) => 
        \ELINK_ADDRA_2[6]_net_1\, ELINK_ADDRA_2(5) => 
        \ELINK_ADDRA_2[5]_net_1\, ELINK_ADDRA_2(4) => 
        \ELINK_ADDRA_2[4]_net_1\, ELINK_ADDRA_2(3) => 
        \ELINK_ADDRA_2[3]_net_1\, ELINK_ADDRA_2(2) => 
        \ELINK_ADDRA_2[2]_net_1\, ELINK_ADDRA_2(1) => 
        \ELINK_ADDRA_2[1]_net_1\, ELINK_ADDRA_2(0) => 
        \ELINK_ADDRA_2[0]_net_1\, PATT_ELK_DAT_2(7) => 
        PATT_ELK_DAT_2(7), PATT_ELK_DAT_2(6) => PATT_ELK_DAT_2(6), 
        PATT_ELK_DAT_2(5) => PATT_ELK_DAT_2(5), PATT_ELK_DAT_2(4)
         => PATT_ELK_DAT_2(4), PATT_ELK_DAT_2(3) => 
        PATT_ELK_DAT_2(3), PATT_ELK_DAT_2(2) => PATT_ELK_DAT_2(2), 
        PATT_ELK_DAT_2(1) => PATT_ELK_DAT_2(1), PATT_ELK_DAT_2(0)
         => PATT_ELK_DAT_2(0), ELINK_DOUTA_2(7) => 
        \ELINK_DOUTA_2[7]\, ELINK_DOUTA_2(6) => 
        \ELINK_DOUTA_2[6]\, ELINK_DOUTA_2(5) => 
        \ELINK_DOUTA_2[5]\, ELINK_DOUTA_2(4) => 
        \ELINK_DOUTA_2[4]\, ELINK_DOUTA_2(3) => 
        \ELINK_DOUTA_2[3]\, ELINK_DOUTA_2(2) => 
        \ELINK_DOUTA_2[2]\, ELINK_DOUTA_2(1) => 
        \ELINK_DOUTA_2[1]\, ELINK_DOUTA_2(0) => 
        \ELINK_DOUTA_2[0]\, ELKS_RWB => ELKS_RWB, 
        P_USB_MASTER_EN_c_0 => P_USB_MASTER_EN_c_0, CLK_40M_GL
         => CLK_40M_GL, CLK60MHZ => CLK60MHZ, ELKS_RAM_BLKB_EN
         => ELKS_RAM_BLKB_EN);
    
    \WR_XFER_TYPE_RNIM29L[5]\ : NOR2
      port map(A => \WR_XFER_TYPE[5]_net_1\, B => \USB_TXE_B\, Y
         => N_1404_7);
    
    \SM_BANK_SEL_RNIGM4B[11]\ : OR2
      port map(A => \SM_BANK_SEL[11]_net_1\, B => 
        \SM_BANK_SEL_0[21]_net_1\, Y => un1_SM_BANK_SEL_21);
    
    \WR_XFER_TYPE_RNO_0[0]\ : NOR3A
      port map(A => N_1736, B => \RD_USB_ADBUS[0]_net_1\, C => 
        N_1702, Y => N_1816);
    
    \RD_USB_ADBUS_RNIRVAJ_3[0]\ : NOR2
      port map(A => \RD_USB_ADBUS[0]_net_1\, B => 
        \RD_USB_ADBUS[1]_net_1\, Y => N_1902);
    
    \ELINK_RWA[13]\ : DFN1E0P0
      port map(D => \N_ELINK_RWA_0_iv[13]\, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_11, E => \SM_BANK_SEL_0[20]_net_1\, 
        Q => \ELINK_RWA[13]_net_1\);
    
    \REG_STATE_ns_i_i_a2_0_2_RNO_2[0]\ : NOR3A
      port map(A => N_274, B => \REG_STATE_0[0]_net_1\, C => 
        N_255, Y => N_412);
    
    \REG_STATE_0_RNI46385[1]\ : OR3
      port map(A => N_2539, B => N_2546, C => N_2537, Y => 
        \REG_STATE_ns_i_1[1]\);
    
    \REG_ADDR_RNINSCP[4]\ : NOR3B
      port map(A => N_261, B => \REG_ADDR[4]_net_1\, C => 
        \SM_BANK_SEL_0[21]_net_1\, Y => \N_TFC_ADDRA[4]\);
    
    \ELINK_ADDRA_15[2]\ : DFN1E0C0
      port map(D => \N_TFC_ADDRA[2]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_6, E => N_199, Q => 
        \ELINK_ADDRA_15[2]_net_1\);
    
    \SM_BANK_SEL_RNO[5]\ : NOR3C
      port map(A => \RD_USB_ADBUS[2]_net_1\, B => N_1892, C => 
        N_1352_4, Y => N_1845);
    
    \WR_USB_ADBUS_RNO_5[1]\ : OR3
      port map(A => \ELINK_DOUTA_3_m[1]\, B => 
        \ELINK_DOUTA_18_m[1]\, C => \N_WR_USB_ADBUS_0_iv_12[1]\, 
        Y => \N_WR_USB_ADBUS_0_iv_20[1]\);
    
    \RD_USB_ADBUS_RNIQO682_0[6]\ : AO1
      port map(A => N_293, B => N_1700, C => N_282, Y => 
        N_1387_i_0_2);
    
    USB_RD_BI_RNO_15 : NOR2A
      port map(A => \REG_STATE[4]_net_1\, B => \USB_RXF_B\, Y => 
        N_1864);
    
    \ELINK_RWA_RNO[3]\ : AOI1
      port map(A => \SM_BANK_SEL[16]_net_1\, B => un1_USB_RXF_B_m, 
        C => \ELINK_RWA_i_m[3]\, Y => \N_ELINK_RWA_0_iv[3]\);
    
    \ELINK_BLKA_RNO[8]\ : AOI1
      port map(A => \SM_BANK_SEL[11]_net_1\, B => X_BLKA_i, C => 
        \ELINK_BLKA_i_m[8]\, Y => \N_ELINK_BLKA_0_iv[8]\);
    
    \RD_USB_ADBUS_RNIEQBG1[7]\ : NOR3B
      port map(A => N_290, B => \RD_USB_ADBUS[7]_net_1\, C => 
        N_1700, Y => N_488);
    
    \ELINK_ADDRA_10[3]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[3]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_22, E => un1_SM_BANK_SEL_20, Q => 
        \ELINK_ADDRA_10[3]_net_1\);
    
    \TFC_STOP_ADDR[1]\ : DFN1E1C0
      port map(D => \TFC_STOP_ADDR_T[1]_net_1\, CLK => CLK60MHZ, 
        CLR => P_USB_MASTER_EN_c_8, E => \REG_STATE_d_0[30]\, Q
         => \TFC_STOP_ADDR[1]_net_1\);
    
    \ELINK_ADDRA_16[7]\ : DFN1E0C0
      port map(D => \N_TFC_ADDRA[7]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_9, E => N_200, Q => 
        \ELINK_ADDRA_16[7]_net_1\);
    
    \N_TFC_ADDRA_0_o2_RNO_0[7]\ : AO1A
      port map(A => \REG_STATE_0[3]_net_1\, B => N_253, C => 
        N_432, Y => N_260);
    
    \ELINK_RWA_RNO_0[2]\ : NOR2A
      port map(A => N_618, B => \ELINK_RWA[2]_net_1\, Y => 
        \ELINK_RWA_i_m[2]\);
    
    \ELINK_RWA[2]\ : DFN1E0P0
      port map(D => \N_ELINK_RWA_0_iv[2]\, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_6, E => \SM_BANK_SEL_0[20]_net_1\, 
        Q => \ELINK_RWA[2]_net_1\);
    
    \ELINK_DINA_12[4]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[4]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_12, E => un1_SM_BANK_SEL_7, Q => 
        \ELINK_DINA_12[4]_net_1\);
    
    \ELINK_RWA_RNO[0]\ : AOI1
      port map(A => \SM_BANK_SEL[19]_net_1\, B => un1_USB_RXF_B_m, 
        C => \ELINK_RWA_i_m[0]\, Y => \N_ELINK_RWA_0_iv[0]\);
    
    \ELINK_BLKA_RNO[15]\ : AOI1B
      port map(A => \SM_BANK_SEL[4]_net_1\, B => X_BLKA_i, C => 
        N_65_tz, Y => N_65);
    
    \SM_BANK_SEL_RNIVJV62[14]\ : NOR3A
      port map(A => \SM_BANK_SEL[14]_net_1\, B => N_312_0, C => 
        N_1566_i_i_0, Y => un1_SM_BANK_SEL_35);
    
    \WR_USB_ADBUS_RNO_9[5]\ : AO1
      port map(A => \ELINK_DOUTA_7[5]\, B => un1_SM_BANK_SEL_37, 
        C => \ELINK_DOUTA_9_m[5]\, Y => 
        \N_WR_USB_ADBUS_0_iv_14[5]\);
    
    \ELINK_DINA_11[3]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[3]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_11, E => un1_SM_BANK_SEL_16, Q => 
        \ELINK_DINA_11[3]_net_1\);
    
    \REG_STATE_RNI3LQN_1[3]\ : OR2
      port map(A => \REG_STATE[3]_net_1\, B => 
        \REG_STATE[4]_net_1\, Y => N_1751);
    
    \WR_USB_ADBUS_RNO_29[6]\ : NOR3B
      port map(A => N_1730_i, B => \ELINKS_STOP_ADDR[6]_net_1\, C
         => N_1726, Y => \ELINKS_STOP_ADDR_m[6]\);
    
    \WR_USB_ADBUS_RNO[1]\ : OR3
      port map(A => \N_WR_USB_ADBUS_0_iv_24[1]\, B => 
        \N_WR_USB_ADBUS_0_iv_23[1]\, C => 
        \N_WR_USB_ADBUS_0_iv_25[1]\, Y => \N_WR_USB_ADBUS[1]\);
    
    \REG_STATE_RNI1JQN[1]\ : NOR2A
      port map(A => \REG_STATE[1]_net_1\, B => 
        \REG_STATE[4]_net_1\, Y => N_1879_1);
    
    \ELINK_ADDRA_18[4]\ : DFN1E0C0
      port map(D => \N_TFC_ADDRA[4]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_12, E => N_198, Q => 
        \ELINK_ADDRA_18[4]_net_1\);
    
    \SM_BANK_SEL_RNIPB7M1[0]\ : OR2B
      port map(A => N_463, B => N_394, Y => 
        \N_ELINK_RWA_0_iv_0_o2_0[18]\);
    
    USB_RXF_B_RNI8TTF3 : OA1
      port map(A => N_2467, B => N_2622, C => \USB_RXF_B\, Y => 
        N_471);
    
    \ELINK_ADDRA_14[3]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[3]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_5, E => un1_SM_BANK_SEL_1, Q => 
        \ELINK_ADDRA_14[3]_net_1\);
    
    \ELINK_ADDRA_15[5]\ : DFN1E0C0
      port map(D => \N_TFC_ADDRA[5]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_6, E => N_199, Q => 
        \ELINK_ADDRA_15[5]_net_1\);
    
    \ELINK_DINA_19[2]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[2]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_0, E => un1_SM_BANK_SEL_11, Q => 
        \ELINK_DINA_19[2]_net_1\);
    
    USB_RD_BI_RNO_9 : OR3
      port map(A => N_USB_RD_BI_i_1, B => N_1865, C => N_1744_i, 
        Y => N_USB_RD_BI_i_4);
    
    \ELINK_DINA_0[7]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[7]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_5, E => un1_SM_BANK_SEL_6, Q => 
        \ELINK_DINA_0[7]_net_1\);
    
    \RD_XFER_TYPE[5]\ : DFN1C0
      port map(D => \RD_XFER_TYPE_RNO[5]_net_1\, CLK => CLK60MHZ, 
        CLR => P_USB_MASTER_EN_c, Q => \RD_XFER_TYPE[5]_net_1\);
    
    \WR_USB_ADBUS_RNO_10[6]\ : AO1
      port map(A => \ELINK_DOUTA_11[6]\, B => un1_SM_BANK_SEL_26, 
        C => \ELINK_DOUTA_12_m[6]\, Y => 
        \N_WR_USB_ADBUS_0_iv_12[6]\);
    
    \ELINK_BLKA_RNO_0[15]\ : AO1
      port map(A => \N_ELINK_RWA_0_iv_0_o2_i_a5_0[15]\, B => 
        N_503, C => \ELINK_BLKA[15]_net_1\, Y => N_65_tz);
    
    USB_RXF_B_RNI3K6I2 : NOR3B
      port map(A => N_USB_OE_BI_iv_0_i_a2_0_1, B => N_385_1, C
         => N_293, Y => \REG_STATE_ns_i_i_a5_1_2[0]\);
    
    \ELINK_ADDRA_7[6]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[6]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_6, E => un1_SM_BANK_SEL_12, Q => 
        \ELINK_ADDRA_7[6]_net_1\);
    
    \CHKSUM_RNO[6]\ : NOR2A
      port map(A => \RD_USB_ADBUS[6]_net_1\, B => N_675, Y => 
        N_228);
    
    \RD_XFER_TYPE_RNO[2]\ : AO1
      port map(A => \RD_XFER_TYPE[2]_net_1\, B => N_1703, C => 
        N_1798, Y => \RD_XFER_TYPE_RNO[2]_net_1\);
    
    USB_TXE_B_RNI1TKL8 : OAI1
      port map(A => REG_STATE_tr74_1, B => REG_STATE_tr67_5, C
         => N_1404_8, Y => \REG_STATE_ns_i_a2_0[1]\);
    
    USB_RD_BI_RNO_4 : NOR2B
      port map(A => N_1862_1, B => N_1728, Y => N_1866);
    
    \WR_XFER_TYPE[2]\ : DFN1C0
      port map(D => \WR_XFER_TYPE_RNO[2]_net_1\, CLK => CLK60MHZ, 
        CLR => P_USB_MASTER_EN_c, Q => \WR_XFER_TYPE[2]_net_1\);
    
    \WR_USB_ADBUS_RNO_11[2]\ : OR3
      port map(A => \N_WR_USB_ADBUS_0_iv_10[2]\, B => 
        \N_WR_USB_ADBUS_0_iv_9[2]\, C => 
        \N_WR_USB_ADBUS_0_iv_20[2]\, Y => 
        \N_WR_USB_ADBUS_0_iv_24[2]\);
    
    \WR_USB_ADBUS[5]\ : DFN1E0C0
      port map(D => \N_WR_USB_ADBUS[5]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_15, E => un1_REG_STATE_26, Q => 
        \WR_USB_ADBUS[5]_net_1\);
    
    \ELINK_BLKA_RNO[16]\ : AOI1
      port map(A => \SM_BANK_SEL[3]_net_1\, B => X_BLKA_i, C => 
        \ELINK_BLKA_i_m[16]\, Y => \N_ELINK_BLKA_0_iv[16]\);
    
    \REG_STATE_0_RNIAD3A1[0]\ : NOR3B
      port map(A => \REG_STATE_0[0]_net_1\, B => 
        \REG_STATE_0[1]_net_1\, C => \REG_STATE_0[2]_net_1\, Y
         => N_1730_i);
    
    \WR_XFER_TYPE_RNO_0[5]\ : NOR2A
      port map(A => N_1698, B => N_1702, Y => N_1829);
    
    \REG_STATE_RNI4CAV2[3]\ : AO1A
      port map(A => N_379, B => N_2602, C => 
        \REG_STATE_ns_i_a4_7_0[1]\, Y => N_1278_tz);
    
    \WR_USB_ADBUS_RNO_21[5]\ : NOR2B
      port map(A => \ELINK_DOUTA_19[5]\, B => un1_SM_BANK_SEL_41, 
        Y => \ELINK_DOUTA_19_m[5]\);
    
    \USB_SIWU_BI\ : DFN1E1P0
      port map(D => N_678, CLK => CLK60MHZ, PRE => 
        P_USB_MASTER_EN_c_8, E => un1_REG_STATE_18, Q => 
        USB_SIWU_BI);
    
    \WR_USB_ADBUS_RNO_1[1]\ : OR3
      port map(A => \N_WR_USB_ADBUS_0_iv_6[1]\, B => 
        \ELINK_DOUTA_14_m[1]\, C => \N_WR_USB_ADBUS_0_iv_18[1]\, 
        Y => \N_WR_USB_ADBUS_0_iv_23[1]\);
    
    \SM_BANK_SEL_RNI6GE7[10]\ : NOR3
      port map(A => \SM_BANK_SEL[11]_net_1\, B => 
        \SM_BANK_SEL[10]_net_1\, C => \SM_BANK_SEL[9]_net_1\, Y
         => N_469);
    
    \REG_STATE_RNI3UN31[2]\ : NOR2A
      port map(A => \REG_STATE[2]_net_1\, B => N_292, Y => 
        \REG_STATE_ns_i_a4_3_0[3]\);
    
    \ELINK_DINA_2[1]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[1]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_9, E => un1_SM_BANK_SEL_5, Q => 
        \ELINK_DINA_2[1]_net_1\);
    
    \ELINK_ADDRA_11[6]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[6]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_2, E => un1_SM_BANK_SEL_16, Q => 
        \ELINK_ADDRA_11[6]_net_1\);
    
    \RD_USB_ADBUS_RNIRVAJ_1[0]\ : NOR2A
      port map(A => \RD_USB_ADBUS[1]_net_1\, B => 
        \RD_USB_ADBUS[0]_net_1\, Y => N_1352_4);
    
    \ELINKS_STOP_ADDR[3]\ : DFN1E1C0
      port map(D => \ELINKS_STOP_ADDR_T[3]_net_1\, CLK => 
        CLK60MHZ, CLR => P_USB_MASTER_EN_c_14, E => 
        \REG_STATE_d_0[30]\, Q => \ELINKS_STOP_ADDR[3]_net_1\);
    
    \ELINK_DINA_16[2]\ : DFN1E0C0
      port map(D => \N_TFC_DINA[2]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_18, E => N_200, Q => 
        \ELINK_DINA_16[2]_net_1\);
    
    \ELINK_DINA_11[0]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[0]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_11, E => un1_SM_BANK_SEL_16, Q => 
        \ELINK_DINA_11[0]_net_1\);
    
    \TFC_DINA[3]\ : DFN1E0C0
      port map(D => \N_TFC_DINA[3]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_4, E => N_142, Q => \TFC_DINA[3]_net_1\);
    
    U101_PATT_ELINK_BLK : DPRT_512X9_SRAM_1
      port map(ELINK_RWA_0 => \ELINK_RWA[1]_net_1\, 
        ELK_RX_SER_WORD_1(7) => ELK_RX_SER_WORD_1(7), 
        ELK_RX_SER_WORD_1(6) => ELK_RX_SER_WORD_1(6), 
        ELK_RX_SER_WORD_1(5) => ELK_RX_SER_WORD_1(5), 
        ELK_RX_SER_WORD_1(4) => ELK_RX_SER_WORD_1(4), 
        ELK_RX_SER_WORD_1(3) => ELK_RX_SER_WORD_1(3), 
        ELK_RX_SER_WORD_1(2) => ELK_RX_SER_WORD_1(2), 
        ELK_RX_SER_WORD_1(1) => ELK_RX_SER_WORD_1(1), 
        ELK_RX_SER_WORD_1(0) => ELK_RX_SER_WORD_1(0), 
        ELINK_DINA_1(7) => \ELINK_DINA_1[7]_net_1\, 
        ELINK_DINA_1(6) => \ELINK_DINA_1[6]_net_1\, 
        ELINK_DINA_1(5) => \ELINK_DINA_1[5]_net_1\, 
        ELINK_DINA_1(4) => \ELINK_DINA_1[4]_net_1\, 
        ELINK_DINA_1(3) => \ELINK_DINA_1[3]_net_1\, 
        ELINK_DINA_1(2) => \ELINK_DINA_1[2]_net_1\, 
        ELINK_DINA_1(1) => \ELINK_DINA_1[1]_net_1\, 
        ELINK_DINA_1(0) => \ELINK_DINA_1[0]_net_1\, ELINK_BLKA_0
         => \ELINK_BLKA[1]_net_1\, ELKS_ADDRB_0_d0 => 
        ELKS_ADDRB(0), ELKS_ADDRB_1 => ELKS_ADDRB(1), 
        ELKS_ADDRB_3 => ELKS_ADDRB(3), ELKS_ADDRB_5 => 
        ELKS_ADDRB(5), ELKS_ADDRB_7 => ELKS_ADDRB(7), 
        ELKS_ADDRB_0_0 => ELKS_ADDRB_0_0, ELKS_ADDRB_0_2 => 
        ELKS_ADDRB_0_2, ELKS_ADDRB_0_4 => ELKS_ADDRB_0_4, 
        ELINK_ADDRA_1(7) => \ELINK_ADDRA_1[7]_net_1\, 
        ELINK_ADDRA_1(6) => \ELINK_ADDRA_1[6]_net_1\, 
        ELINK_ADDRA_1(5) => \ELINK_ADDRA_1[5]_net_1\, 
        ELINK_ADDRA_1(4) => \ELINK_ADDRA_1[4]_net_1\, 
        ELINK_ADDRA_1(3) => \ELINK_ADDRA_1[3]_net_1\, 
        ELINK_ADDRA_1(2) => \ELINK_ADDRA_1[2]_net_1\, 
        ELINK_ADDRA_1(1) => \ELINK_ADDRA_1[1]_net_1\, 
        ELINK_ADDRA_1(0) => \ELINK_ADDRA_1[0]_net_1\, 
        PATT_ELK_DAT_1(7) => PATT_ELK_DAT_1(7), PATT_ELK_DAT_1(6)
         => PATT_ELK_DAT_1(6), PATT_ELK_DAT_1(5) => 
        PATT_ELK_DAT_1(5), PATT_ELK_DAT_1(4) => PATT_ELK_DAT_1(4), 
        PATT_ELK_DAT_1(3) => PATT_ELK_DAT_1(3), PATT_ELK_DAT_1(2)
         => PATT_ELK_DAT_1(2), PATT_ELK_DAT_1(1) => 
        PATT_ELK_DAT_1(1), PATT_ELK_DAT_1(0) => PATT_ELK_DAT_1(0), 
        ELINK_DOUTA_1(7) => \ELINK_DOUTA_1[7]\, ELINK_DOUTA_1(6)
         => \ELINK_DOUTA_1[6]\, ELINK_DOUTA_1(5) => 
        \ELINK_DOUTA_1[5]\, ELINK_DOUTA_1(4) => 
        \ELINK_DOUTA_1[4]\, ELINK_DOUTA_1(3) => 
        \ELINK_DOUTA_1[3]\, ELINK_DOUTA_1(2) => 
        \ELINK_DOUTA_1[2]\, ELINK_DOUTA_1(1) => 
        \ELINK_DOUTA_1[1]\, ELINK_DOUTA_1(0) => 
        \ELINK_DOUTA_1[0]\, ELKS_RWB => ELKS_RWB, 
        P_USB_MASTER_EN_c_0 => P_USB_MASTER_EN_c_0, CLK_40M_GL
         => CLK_40M_GL, CLK60MHZ => CLK60MHZ, ELKS_RAM_BLKB_EN
         => ELKS_RAM_BLKB_EN);
    
    \ELINK_DINA_13[5]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[5]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_14, E => un1_SM_BANK_SEL_2, Q => 
        \ELINK_DINA_13[5]_net_1\);
    
    \WR_XFER_TYPE_RNO[1]\ : NOR3
      port map(A => N_1819, B => N_1821, C => N_1820, Y => 
        \WR_XFER_TYPE_RNO[1]_net_1\);
    
    \ELINK_RWA_RNO[6]\ : AOI1
      port map(A => \SM_BANK_SEL[13]_net_1\, B => un1_USB_RXF_B_m, 
        C => \ELINK_RWA_i_m[6]\, Y => \N_ELINK_RWA_0_iv[6]\);
    
    \SM_BANK_SEL_RNIL4M41[7]\ : NOR3B
      port map(A => N_469, B => N_477, C => 
        \SM_BANK_SEL[7]_net_1\, Y => 
        \N_ELINK_BLKA_0_iv_0_o2_i_a5_1[11]\);
    
    \ELINK_DINA_19[6]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[6]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_1, E => un1_SM_BANK_SEL_11, Q => 
        \ELINK_DINA_19[6]_net_1\);
    
    \ELINK_BLKA_RNO_0[12]\ : OA1B
      port map(A => N_624_15, B => \N_ELINK_RWA_1[12]\, C => 
        \ELINK_BLKA[12]_net_1\, Y => \ELINK_BLKA_i_m[12]\);
    
    \WR_USB_ADBUS_RNO_25[7]\ : NOR2B
      port map(A => \ELINK_DOUTA_11[7]\, B => un1_SM_BANK_SEL_26, 
        Y => \ELINK_DOUTA_11_m[7]\);
    
    USB_RD_BI_RNO_13 : OR3
      port map(A => N_1864, B => \REG_STATE_0[5]_net_1\, C => 
        N_1359_2, Y => N_USB_RD_BI_i_1);
    
    \WR_USB_ADBUS_RNO_7[4]\ : AO1
      port map(A => \ELINK_DOUTA_4[4]\, B => un1_SM_BANK_SEL_28, 
        C => \ELINK_DOUTA_5_m[4]\, Y => 
        \N_WR_USB_ADBUS_0_iv_7[4]\);
    
    \REG_STATE_RNIVGQN_2[0]\ : OR2
      port map(A => \REG_STATE[0]_net_1\, B => 
        \REG_STATE[3]_net_1\, Y => N_257);
    
    \OP_MODE_T[0]\ : DFN1E1C0
      port map(D => \RD_USB_ADBUS[0]_net_1\, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_17, E => N_OP_MODE_T_0_sqmuxa, Q
         => \OP_MODE_T[0]_net_1\);
    
    \REG_STATE_ns_i_i_a2_0_2[0]\ : AND2
      port map(A => N_414_i, B => \REG_STATE_ns_i_i_a2_0_1[0]\, Y
         => \REG_STATE_ns_i_i_a2_0_2[0]_net_1\);
    
    \RD_XFER_TYPE_RNO_0[2]\ : NOR2A
      port map(A => \RD_USB_ADBUS[2]_net_1\, B => N_1694, Y => 
        N_1798);
    
    \ELINK_DINA_2[3]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[3]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_9, E => un1_SM_BANK_SEL_5, Q => 
        \ELINK_DINA_2[3]_net_1\);
    
    \TFC_DINA[2]\ : DFN1E0C0
      port map(D => \N_TFC_DINA[2]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_4, E => N_142, Q => \TFC_DINA[2]_net_1\);
    
    \SM_BANK_SEL_0[20]\ : DFN1E1C0
      port map(D => un1_N_ELK_N_ACTIVE_2_sqmuxa, CLK => CLK60MHZ, 
        CLR => P_USB_MASTER_EN_c_1_0, E => un1_REG_STATE_30, Q
         => \SM_BANK_SEL_0[20]_net_1\);
    
    \ELINK_DINA_6[4]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[4]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_16, E => un1_SM_BANK_SEL_10, Q => 
        \ELINK_DINA_6[4]_net_1\);
    
    \ELINK_DINA_4[0]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[0]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_12, E => un1_SM_BANK_SEL_8, Q => 
        \ELINK_DINA_4[0]_net_1\);
    
    \WR_USB_ADBUS_RNO_24[5]\ : NOR2B
      port map(A => \ELINK_DOUTA_6[5]\, B => un1_SM_BANK_SEL_30, 
        Y => \ELINK_DOUTA_6_m[5]\);
    
    \SM_BANK_SEL[12]\ : DFN1E1C0
      port map(D => N_1833, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_1_0, E => un1_REG_STATE_30, Q => 
        \SM_BANK_SEL[12]_net_1\);
    
    USB_RD_BI_RNO_2 : OR3
      port map(A => N_1869, B => N_1868, C => N_USB_RD_BI_i_4, Y
         => N_USB_RD_BI_i_5);
    
    \WR_USB_ADBUS_RNO_18[6]\ : NOR2B
      port map(A => \ELINK_DOUTA_4[6]\, B => un1_SM_BANK_SEL_28, 
        Y => \ELINK_DOUTA_4_m[6]\);
    
    U106_PATT_ELINK_BLK : DPRT_512X9_SRAM_6
      port map(ELINK_RWA_0 => \ELINK_RWA[6]_net_1\, 
        ELK_RX_SER_WORD_6(7) => ELK_RX_SER_WORD_6(7), 
        ELK_RX_SER_WORD_6(6) => ELK_RX_SER_WORD_6(6), 
        ELK_RX_SER_WORD_6(5) => ELK_RX_SER_WORD_6(5), 
        ELK_RX_SER_WORD_6(4) => ELK_RX_SER_WORD_6(4), 
        ELK_RX_SER_WORD_6(3) => ELK_RX_SER_WORD_6(3), 
        ELK_RX_SER_WORD_6(2) => ELK_RX_SER_WORD_6(2), 
        ELK_RX_SER_WORD_6(1) => ELK_RX_SER_WORD_6(1), 
        ELK_RX_SER_WORD_6(0) => ELK_RX_SER_WORD_6(0), 
        ELINK_DINA_6(7) => \ELINK_DINA_6[7]_net_1\, 
        ELINK_DINA_6(6) => \ELINK_DINA_6[6]_net_1\, 
        ELINK_DINA_6(5) => \ELINK_DINA_6[5]_net_1\, 
        ELINK_DINA_6(4) => \ELINK_DINA_6[4]_net_1\, 
        ELINK_DINA_6(3) => \ELINK_DINA_6[3]_net_1\, 
        ELINK_DINA_6(2) => \ELINK_DINA_6[2]_net_1\, 
        ELINK_DINA_6(1) => \ELINK_DINA_6[1]_net_1\, 
        ELINK_DINA_6(0) => \ELINK_DINA_6[0]_net_1\, ELINK_BLKA_0
         => \ELINK_BLKA[6]_net_1\, ELKS_ADDRB_0_d0 => 
        ELKS_ADDRB(0), ELKS_ADDRB_1 => ELKS_ADDRB(1), 
        ELKS_ADDRB_3 => ELKS_ADDRB(3), ELKS_ADDRB_5 => 
        ELKS_ADDRB(5), ELKS_ADDRB_7 => ELKS_ADDRB(7), 
        ELKS_ADDRB_0_0 => ELKS_ADDRB_0_0, ELKS_ADDRB_0_2 => 
        ELKS_ADDRB_0_2, ELKS_ADDRB_0_4 => ELKS_ADDRB_0_4, 
        ELINK_ADDRA_6(7) => \ELINK_ADDRA_6[7]_net_1\, 
        ELINK_ADDRA_6(6) => \ELINK_ADDRA_6[6]_net_1\, 
        ELINK_ADDRA_6(5) => \ELINK_ADDRA_6[5]_net_1\, 
        ELINK_ADDRA_6(4) => \ELINK_ADDRA_6[4]_net_1\, 
        ELINK_ADDRA_6(3) => \ELINK_ADDRA_6[3]_net_1\, 
        ELINK_ADDRA_6(2) => \ELINK_ADDRA_6[2]_net_1\, 
        ELINK_ADDRA_6(1) => \ELINK_ADDRA_6[1]_net_1\, 
        ELINK_ADDRA_6(0) => \ELINK_ADDRA_6[0]_net_1\, 
        PATT_ELK_DAT_6(7) => PATT_ELK_DAT_6(7), PATT_ELK_DAT_6(6)
         => PATT_ELK_DAT_6(6), PATT_ELK_DAT_6(5) => 
        PATT_ELK_DAT_6(5), PATT_ELK_DAT_6(4) => PATT_ELK_DAT_6(4), 
        PATT_ELK_DAT_6(3) => PATT_ELK_DAT_6(3), PATT_ELK_DAT_6(2)
         => PATT_ELK_DAT_6(2), PATT_ELK_DAT_6(1) => 
        PATT_ELK_DAT_6(1), PATT_ELK_DAT_6(0) => PATT_ELK_DAT_6(0), 
        ELINK_DOUTA_6(7) => \ELINK_DOUTA_6[7]\, ELINK_DOUTA_6(6)
         => \ELINK_DOUTA_6[6]\, ELINK_DOUTA_6(5) => 
        \ELINK_DOUTA_6[5]\, ELINK_DOUTA_6(4) => 
        \ELINK_DOUTA_6[4]\, ELINK_DOUTA_6(3) => 
        \ELINK_DOUTA_6[3]\, ELINK_DOUTA_6(2) => 
        \ELINK_DOUTA_6[2]\, ELINK_DOUTA_6(1) => 
        \ELINK_DOUTA_6[1]\, ELINK_DOUTA_6(0) => 
        \ELINK_DOUTA_6[0]\, ELKS_RWB => ELKS_RWB, 
        P_USB_MASTER_EN_c_0 => P_USB_MASTER_EN_c_0, CLK_40M_GL
         => CLK_40M_GL, CLK60MHZ => CLK60MHZ, ELKS_RAM_BLKB_EN
         => ELKS_RAM_BLKB_EN);
    
    \ELINK_ADDRA_19[6]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[6]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_13, E => un1_SM_BANK_SEL_11, Q => 
        \ELINK_ADDRA_19[6]_net_1\);
    
    \RD_XFER_TYPE_RNO[3]\ : AO1
      port map(A => \RD_XFER_TYPE[3]_net_1\, B => N_1703, C => 
        N_1800, Y => \RD_XFER_TYPE_RNO[3]_net_1\);
    
    \ELINK_ADDRA_10[4]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[4]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_22, E => un1_SM_BANK_SEL_20, Q => 
        \ELINK_ADDRA_10[4]_net_1\);
    
    \ELINK_DINA_5[2]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[2]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_14, E => un1_SM_BANK_SEL_15, Q => 
        \ELINK_DINA_5[2]_net_1\);
    
    \ELINK_DINA_14[2]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[2]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_16, E => un1_SM_BANK_SEL_1, Q => 
        \ELINK_DINA_14[2]_net_1\);
    
    \REG_STATE_ns_i_8_tz_0_RNO[4]\ : NOR2B
      port map(A => N_1879_1, B => N_287, Y => 
        \REG_STATE_ns_i_a4_2_0[4]\);
    
    \ELINK_RWA[10]\ : DFN1E0P0
      port map(D => \N_ELINK_RWA_0_iv[10]\, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_11, E => \SM_BANK_SEL_0[20]_net_1\, 
        Q => \ELINK_RWA[10]_net_1\);
    
    \OP_MODE[5]\ : DFN1E1C0
      port map(D => \OP_MODE_T[5]_net_1\, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_15, E => \REG_STATE_d[30]\, Q => 
        \OP_MODE[5]_net_1\);
    
    \WR_USB_ADBUS_RNO_12[2]\ : NOR2B
      port map(A => \ELINK_DOUTA_18[2]\, B => un1_SM_BANK_SEL_25, 
        Y => \ELINK_DOUTA_18_m[2]\);
    
    \ELINK_DINA_11[4]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[4]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_11, E => un1_SM_BANK_SEL_16, Q => 
        \ELINK_DINA_11[4]_net_1\);
    
    \ELINK_DINA_15[3]\ : DFN1E0C0
      port map(D => \N_TFC_DINA[3]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_16, E => N_199, Q => 
        \ELINK_DINA_15[3]_net_1\);
    
    \WR_USB_ADBUS_RNO_14[0]\ : NOR2B
      port map(A => \ELINK_DOUTA_13[0]\, B => un1_SM_BANK_SEL_29, 
        Y => \ELINK_DOUTA_13_m[0]\);
    
    \SM_BANK_SEL_RNIHN4B[12]\ : OR2
      port map(A => \SM_BANK_SEL[12]_net_1\, B => 
        \SM_BANK_SEL_0[21]_net_1\, Y => un1_SM_BANK_SEL_12);
    
    \RD_USB_ADBUS_RNI42PD4[4]\ : OR3A
      port map(A => N_290, B => \RD_USB_ADBUS[4]_net_1\, C => 
        N_1717, Y => N_1763);
    
    \SM_BANK_SEL_RNIU5VN[13]\ : OR3A
      port map(A => N_143, B => N_620_10, C => \N_ELINK_RWA_1[5]\, 
        Y => \N_ELINK_RWA_3[5]\);
    
    \ELINK_BLKA[13]\ : DFN1E0P0
      port map(D => N_67, CLK => CLK60MHZ, PRE => 
        P_USB_MASTER_EN_c_20, E => \SM_BANK_SEL[20]_net_1\, Q => 
        \ELINK_BLKA[13]_net_1\);
    
    \ELINK_ADDRA_10[7]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[7]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_22, E => un1_SM_BANK_SEL_20, Q => 
        \ELINK_ADDRA_10[7]_net_1\);
    
    \ELINK_DINA_0[2]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[2]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_5, E => un1_SM_BANK_SEL_6, Q => 
        \ELINK_DINA_0[2]_net_1\);
    
    \N_WR_USB_ADBUS_0_iv_0[4]\ : OR2
      port map(A => \TFC_STOP_ADDR_m[4]\, B => N_1562_i, Y => 
        \N_WR_USB_ADBUS_0_iv_0[4]_net_1\);
    
    \SM_BANK_SEL_RNIMSL6[7]\ : OR2
      port map(A => \SM_BANK_SEL[7]_net_1\, B => 
        \SM_BANK_SEL[21]_net_1\, Y => un1_SM_BANK_SEL_7);
    
    \REG_ADDR_RNIKF203[6]\ : NOR3C
      port map(A => REG_STATE_tr73_7, B => REG_STATE_tr73_6, C
         => N_1421_3, Y => REG_STATE_tr73_9);
    
    \WR_XFER_TYPE_RNI5LLM2_0[0]\ : NOR3C
      port map(A => N_1404_6, B => REG_STATE_tr67_0, C => 
        REG_STATE_tr67_1, Y => REG_STATE_tr67_3);
    
    \REG_STATE_RNIOVPD3[1]\ : NOR2A
      port map(A => N_254, B => \REG_STATE[1]_net_1\, Y => N_1704);
    
    \WR_USB_ADBUS[0]\ : DFN1E0C0
      port map(D => \N_WR_USB_ADBUS[0]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_15, E => un1_REG_STATE_26, Q => 
        \WR_USB_ADBUS[0]_net_1\);
    
    \REG_STATE_RNIVTCJ2[0]\ : MX2
      port map(A => \REG_STATE_ns_i_a4_3_1_0[1]\, B => N_2628, S
         => N_2477_i, Y => N_1275_tz);
    
    \N_TFC_ADDRA_0_a2_2[7]\ : AND2
      port map(A => N_1704, B => N_251, Y => N_429);
    
    \ELINKS_STOP_ADDR_T[7]\ : DFN1E1C0
      port map(D => \RD_USB_ADBUS[7]_net_1\, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_7, E => 
        N_ELINKS_STOP_ADDR_T_0_sqmuxa, Q => 
        \ELINKS_STOP_ADDR_T[7]_net_1\);
    
    U4E_REGCROSS : CLK60M_TO_40M_0
      port map(OP_MODE(7) => \OP_MODE[7]_net_1\, OP_MODE(6) => 
        \OP_MODE[6]_net_1\, OP_MODE(5) => \OP_MODE[5]_net_1\, 
        OP_MODE(4) => \OP_MODE_0[4]\, OP_MODE(3) => 
        \OP_MODE[3]_net_1\, OP_MODE(2) => \OP_MODE[2]_net_1\, 
        OP_MODE(1) => \OP_MODE[1]_net_1\, OP_MODE(0) => 
        \OP_MODE_0[0]\, OP_MODE_0_0 => \OP_MODE[0]_net_1\, 
        OP_MODE_0_4 => \OP_MODE[4]_net_1\, OP_MODE_c_1_d0 => 
        OP_MODE_c_1_d0, OP_MODE_c_5_d0 => OP_MODE_c_5_d0, 
        OP_MODE_c_4_d0 => OP_MODE_c_4_d0, OP_MODE_c_0_d0 => 
        OP_MODE_c_0_d0, OP_MODE_c_0_0 => OP_MODE_c_0_0, 
        OP_MODE_c_1_0 => OP_MODE_c_1_0, OP_MODE_c_2_0 => 
        OP_MODE_c_2_0, OP_MODE_c_3_0 => OP_MODE_c_3_0, 
        OP_MODE_c_4_0 => OP_MODE_c_4_0, OP_MODE_c_5_0 => 
        OP_MODE_c_5_0, OP_MODE_c_6_0 => OP_MODE_c_6_0, 
        P_MASTER_POR_B_c_25 => P_MASTER_POR_B_c_25, 
        P_MASTER_POR_B_c_24 => P_MASTER_POR_B_c_24, 
        P_MASTER_POR_B_c_23 => P_MASTER_POR_B_c_23, 
        P_MASTER_POR_B_c_6 => P_MASTER_POR_B_c_6, 
        P_MASTER_POR_B_c => P_MASTER_POR_B_c, P_MASTER_POR_B_c_1
         => P_MASTER_POR_B_c_1, P_MASTER_POR_B_c_0_0 => 
        P_MASTER_POR_B_c_0_0, CLK_40M_GL => CLK_40M_GL);
    
    \SM_BANK_SEL_RNII64B1[0]\ : NOR3C
      port map(A => N_463, B => N_464, C => N_486, Y => N_503);
    
    \WR_USB_ADBUS_RNO_3[0]\ : AO1
      port map(A => \ELINK_DOUTA_10[0]\, B => un1_SM_BANK_SEL_34, 
        C => \ELINK_DOUTA_11_m[0]\, Y => 
        \N_WR_USB_ADBUS_0_iv_10[0]\);
    
    \WR_USB_ADBUS_RNO_26[3]\ : NOR2B
      port map(A => \ELINK_DOUTA_10[3]\, B => un1_SM_BANK_SEL_34, 
        Y => \ELINK_DOUTA_10_m[3]\);
    
    \REG_STATE_RNIUSCJ2[1]\ : AO1A
      port map(A => N_1352_1, B => N_2526_1, C => N_1745_i, Y => 
        un1_REG_STATE_26_0_1);
    
    \RD_USB_ADBUS_RNINBIK2[2]\ : NOR2A
      port map(A => \RD_USB_ADBUS[2]_net_1\, B => N_206, Y => 
        \N_TFC_DINA[2]\);
    
    \WR_XFER_TYPE[4]\ : DFN1C0
      port map(D => \WR_XFER_TYPE_RNO[4]_net_1\, CLK => CLK60MHZ, 
        CLR => P_USB_MASTER_EN_c, Q => \WR_XFER_TYPE[4]_net_1\);
    
    \ELINKS_STOP_ADDR[0]\ : DFN1E1C0
      port map(D => \ELINKS_STOP_ADDR_T[0]_net_1\, CLK => 
        CLK60MHZ, CLR => P_USB_MASTER_EN_c_14, E => 
        \REG_STATE_d_0[30]\, Q => \ELINKS_STOP_ADDR[0]_net_1\);
    
    \WR_USB_ADBUS_RNO_7[5]\ : NOR2B
      port map(A => \ELINK_DOUTA_14[5]\, B => un1_SM_BANK_SEL_23, 
        Y => \ELINK_DOUTA_14_m[5]\);
    
    \ELINK_ADDRA_1[5]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[5]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_20, E => un1_SM_BANK_SEL_19, Q => 
        \ELINK_ADDRA_1[5]_net_1\);
    
    \SM_BANK_SEL_RNIS3VN[15]\ : OR3A
      port map(A => N_143, B => N_616_11, C => \N_ELINK_RWA_1[3]\, 
        Y => \N_ELINK_RWA_3[3]\);
    
    \WR_USB_ADBUS_RNO_21[6]\ : NOR2B
      port map(A => \ELINK_DOUTA_3[6]\, B => un1_SM_BANK_SEL_43, 
        Y => \ELINK_DOUTA_3_m[6]\);
    
    \RD_XFER_TYPE_RNO_0[1]\ : NOR2A
      port map(A => \RD_USB_ADBUS[1]_net_1\, B => N_1694, Y => 
        N_1796);
    
    U3_USB_DAT_BUS : BIDIR_LVTTL
      port map(WR_USB_ADBUS(7) => \WR_USB_ADBUS[7]_net_1\, 
        WR_USB_ADBUS(6) => \WR_USB_ADBUS[6]_net_1\, 
        WR_USB_ADBUS(5) => \WR_USB_ADBUS[5]_net_1\, 
        WR_USB_ADBUS(4) => \WR_USB_ADBUS[4]_net_1\, 
        WR_USB_ADBUS(3) => \WR_USB_ADBUS[3]_net_1\, 
        WR_USB_ADBUS(2) => \WR_USB_ADBUS[2]_net_1\, 
        WR_USB_ADBUS(1) => \WR_USB_ADBUS[1]_net_1\, 
        WR_USB_ADBUS(0) => \WR_USB_ADBUS[0]_net_1\, 
        N_RD_USB_ADBUS(7) => \N_RD_USB_ADBUS[7]\, 
        N_RD_USB_ADBUS(6) => \N_RD_USB_ADBUS[6]\, 
        N_RD_USB_ADBUS(5) => \N_RD_USB_ADBUS[5]\, 
        N_RD_USB_ADBUS(4) => \N_RD_USB_ADBUS[4]\, 
        N_RD_USB_ADBUS(3) => \N_RD_USB_ADBUS[3]\, 
        N_RD_USB_ADBUS(2) => \N_RD_USB_ADBUS[2]\, 
        N_RD_USB_ADBUS(1) => \N_RD_USB_ADBUS[1]\, 
        N_RD_USB_ADBUS(0) => \N_RD_USB_ADBUS[0]\, 
        BIDIR_USB_ADBUS(7) => BIDIR_USB_ADBUS(7), 
        BIDIR_USB_ADBUS(6) => BIDIR_USB_ADBUS(6), 
        BIDIR_USB_ADBUS(5) => BIDIR_USB_ADBUS(5), 
        BIDIR_USB_ADBUS(4) => BIDIR_USB_ADBUS(4), 
        BIDIR_USB_ADBUS(3) => BIDIR_USB_ADBUS(3), 
        BIDIR_USB_ADBUS(2) => BIDIR_USB_ADBUS(2), 
        BIDIR_USB_ADBUS(1) => BIDIR_USB_ADBUS(1), 
        BIDIR_USB_ADBUS(0) => BIDIR_USB_ADBUS(0), TrienAux => 
        TrienAux);
    
    \REG_STATE_ns_i_i_a2_0_2_RNO[0]\ : OR3C
      port map(A => N_1499_2_i_0, B => \REG_STATE_0[2]_net_1\, C
         => N_414_1, Y => N_414_i);
    
    \WR_USB_ADBUS_RNO_2[3]\ : OR3
      port map(A => \N_WR_USB_ADBUS_0_iv_14[3]\, B => 
        \N_WR_USB_ADBUS_0_iv_13[3]\, C => 
        \N_WR_USB_ADBUS_0_iv_22[3]\, Y => 
        \N_WR_USB_ADBUS_0_iv_25[3]\);
    
    \SM_BANK_SEL[13]\ : DFN1E1C0
      port map(D => N_1844, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_1_0, E => un1_REG_STATE_30, Q => 
        \SM_BANK_SEL[13]_net_1\);
    
    \ELINK_ADDRA_9[7]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[7]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_10, E => un1_SM_BANK_SEL_9, Q => 
        \ELINK_ADDRA_9[7]_net_1\);
    
    \WR_USB_ADBUS_RNO_7[2]\ : NOR2A
      port map(A => \TFC_DOUTA[2]\, B => N_243, Y => 
        \TFC_DOUTA_m[2]\);
    
    \ELINK_DINA_17[4]\ : DFN1E0C0
      port map(D => \N_TFC_DINA[4]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_19, E => N_197, Q => 
        \ELINK_DINA_17[4]_net_1\);
    
    \ELINK_DINA_15[5]\ : DFN1E0C0
      port map(D => \N_TFC_DINA[5]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_16, E => N_199, Q => 
        \ELINK_DINA_15[5]_net_1\);
    
    \WR_USB_ADBUS_RNO_1[5]\ : OR3
      port map(A => \N_WR_USB_ADBUS_0_iv_6[5]\, B => 
        \ELINK_DOUTA_14_m[5]\, C => \N_WR_USB_ADBUS_0_iv_18[5]\, 
        Y => \N_WR_USB_ADBUS_0_iv_23[5]\);
    
    \REG_STATE_RNI4TOT[0]\ : NOR2B
      port map(A => N_2613, B => \REG_STATE[0]_net_1\, Y => 
        N_2617);
    
    \TFC_ADDRA[3]\ : DFN1E0C0
      port map(D => \N_TFC_ADDRA[3]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_9, E => N_142, Q => 
        \TFC_ADDRA[3]_net_1\);
    
    \SM_BANK_SEL_RNI4PV62[19]\ : NOR3A
      port map(A => \SM_BANK_SEL[19]_net_1\, B => N_312_0, C => 
        N_1566_i_i_0, Y => un1_SM_BANK_SEL_31);
    
    \CHKSUM[2]\ : DFN1E1C0
      port map(D => N_234, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_3, E => un1_REG_STATE_22, Q => 
        \CHKSUM[2]_net_1\);
    
    \RD_XFER_TYPE_RNIRNMR[2]\ : OR2
      port map(A => \RD_XFER_TYPE[3]_net_1\, B => 
        \RD_XFER_TYPE[2]_net_1\, Y => N_1367_i_i_o2_0_0);
    
    \ELINK_DINA_0[0]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[0]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_5, E => un1_SM_BANK_SEL_6, Q => 
        \ELINK_DINA_0[0]_net_1\);
    
    \REG_STATE_RNI9K186[1]\ : OR2
      port map(A => N_1905, B => N_1704, Y => X_BLKA_i);
    
    \WR_USB_ADBUS_RNO_7[7]\ : NOR2B
      port map(A => \ELINK_DOUTA_14[7]\, B => un1_SM_BANK_SEL_23, 
        Y => \ELINK_DOUTA_14_m[7]\);
    
    \ELINK_ADDRA_11[0]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[0]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_2, E => un1_SM_BANK_SEL_16, Q => 
        \ELINK_ADDRA_11[0]_net_1\);
    
    USB_RD_BI_RNO_0 : AO1D
      port map(A => un1_REG_STATE_40_i_o2_0, B => N_1756, C => 
        N_1862, Y => N_1675);
    
    \SM_BANK_SEL_RNI9CHH[4]\ : NOR3
      port map(A => \SM_BANK_SEL[6]_net_1\, B => 
        \SM_BANK_SEL[5]_net_1\, C => \SM_BANK_SEL[4]_net_1\, Y
         => \N_ELINK_RWA_i_a2_0_a5_0[16]\);
    
    \SM_BANK_SEL[21]\ : DFN1E1P0
      port map(D => N_1671, CLK => CLK60MHZ, PRE => 
        P_USB_MASTER_EN_c_2, E => un1_REG_STATE_30, Q => 
        \SM_BANK_SEL[21]_net_1\);
    
    \REG_STATE_RNI0IQN[1]\ : NOR2
      port map(A => \REG_STATE[1]_net_1\, B => 
        \REG_STATE[3]_net_1\, Y => N_1690_i);
    
    \WR_USB_ADBUS_RNO_31[0]\ : NOR3B
      port map(A => N_1730_i, B => \ELINKS_STOP_ADDR[0]_net_1\, C
         => N_1726, Y => \ELINKS_STOP_ADDR_m[0]\);
    
    \REG_STATE_ns_i_i_a2_0_RNIIQGG5[0]\ : AO1A
      port map(A => N_244_1, B => 
        \REG_STATE_ns_i_i_a2_0[0]_net_1\, C => N_421, Y => 
        N_511_1);
    
    \RD_XFER_TYPE[2]\ : DFN1C0
      port map(D => \RD_XFER_TYPE_RNO[2]_net_1\, CLK => CLK60MHZ, 
        CLR => P_USB_MASTER_EN_c, Q => \RD_XFER_TYPE[2]_net_1\);
    
    \ELINK_DINA_1[1]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[1]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_7, E => un1_SM_BANK_SEL_19, Q => 
        \ELINK_DINA_1[1]_net_1\);
    
    \WR_USB_ADBUS_RNO[3]\ : OR3
      port map(A => \N_WR_USB_ADBUS_0_iv_24[3]\, B => 
        \N_WR_USB_ADBUS_0_iv_23[3]\, C => 
        \N_WR_USB_ADBUS_0_iv_25[3]\, Y => \N_WR_USB_ADBUS[3]\);
    
    \SM_BANK_SEL_RNI0AK1[10]\ : OR2
      port map(A => \SM_BANK_SEL[10]_net_1\, B => 
        \SM_BANK_SEL[21]_net_1\, Y => un1_SM_BANK_SEL_9);
    
    \SM_BANK_SEL_RNIIO4B[13]\ : OR2
      port map(A => \SM_BANK_SEL[13]_net_1\, B => 
        \SM_BANK_SEL_0[21]_net_1\, Y => un1_SM_BANK_SEL_10);
    
    \RD_USB_ADBUS_RNIP4GES[4]\ : NOR2A
      port map(A => N_1294_tz, B => N_311, Y => 
        \RD_USB_ADBUS_RNIP4GES[4]_net_1\);
    
    \WR_USB_ADBUS_RNO_17[0]\ : NOR2B
      port map(A => \ELINK_DOUTA_7[0]\, B => un1_SM_BANK_SEL_37, 
        Y => \ELINK_DOUTA_7_m[0]\);
    
    \WR_USB_ADBUS_RNO_15[2]\ : NOR2B
      port map(A => \ELINK_DOUTA_4[2]\, B => un1_SM_BANK_SEL_28, 
        Y => \ELINK_DOUTA_4_m[2]\);
    
    \SM_BANK_SEL_RNO[16]\ : NOR3A
      port map(A => N_1882, B => N_1700, C => N_290, Y => N_1835);
    
    \ELINK_RWA_RNO[14]\ : AOI1
      port map(A => \SM_BANK_SEL[5]_net_1\, B => un1_USB_RXF_B_m, 
        C => \ELINK_RWA_i_m[14]\, Y => \N_ELINK_RWA_0_iv[14]\);
    
    \ELINK_DINA_9[6]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[6]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_20, E => un1_SM_BANK_SEL_9, Q => 
        \ELINK_DINA_9[6]_net_1\);
    
    \ELINK_DINA_9[1]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[1]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_19, E => un1_SM_BANK_SEL_9, Q => 
        \ELINK_DINA_9[1]_net_1\);
    
    \RD_USB_ADBUS_RNIPADT2[7]\ : OR2A
      port map(A => \RD_USB_ADBUS[7]_net_1\, B => N_1697, Y => 
        N_1702);
    
    \WR_USB_ADBUS_RNO_11[3]\ : OR3
      port map(A => \ELINK_DOUTA_11_m[3]\, B => 
        \ELINK_DOUTA_10_m[3]\, C => \N_WR_USB_ADBUS_0_iv_16[3]\, 
        Y => \N_WR_USB_ADBUS_0_iv_22[3]\);
    
    \REG_STATE_0_RNIAD3A1_0[0]\ : NOR3A
      port map(A => \REG_STATE_0[0]_net_1\, B => 
        \REG_STATE_0[2]_net_1\, C => \REG_STATE_0[1]_net_1\, Y
         => N_1744_i);
    
    \ELINK_ADDRA_17[7]\ : DFN1E0C0
      port map(D => \N_TFC_ADDRA[7]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_11, E => N_197, Q => 
        \ELINK_ADDRA_17[7]_net_1\);
    
    \WR_USB_ADBUS_RNO[7]\ : OR3
      port map(A => \N_WR_USB_ADBUS_0_iv_24[7]\, B => 
        \N_WR_USB_ADBUS_0_iv_23[7]\, C => 
        \N_WR_USB_ADBUS_0_iv_25[7]\, Y => \N_WR_USB_ADBUS[7]\);
    
    USB_RXF_B_0_RNI27AB1 : OA1C
      port map(A => \REG_STATE_0[3]_net_1\, B => \USB_RXF_B_0\, C
         => \REG_STATE_0[4]_net_1\, Y => 
        un1_REG_STATE_40_i_a2_3_0);
    
    \WR_USB_ADBUS_RNO_30[3]\ : NOR3B
      port map(A => N_1352_1, B => \OP_MODE[3]_net_1\, C => 
        REG_STATE_s20_i_0, Y => \OP_MODE_m[3]\);
    
    \SM_BANK_SEL_RNO[1]\ : NOR3B
      port map(A => un1_N_ELK_N_ACTIVE_0_sqmuxa_15_0_a2_0_0, B
         => N_1352_4, C => N_1697, Y => N_1850);
    
    \REG_STATE_RNI2FIR1[4]\ : NOR2B
      port map(A => N_2537_1, B => N_2497, Y => N_2537);
    
    \N_TFC_ADDRA_0_o2_RNO_3[7]\ : NOR3A
      port map(A => \REG_STATE_0[0]_net_1\, B => 
        \REG_STATE_0[2]_net_1\, C => N_259, Y => N_432);
    
    \WR_USB_ADBUS_RNO_18[7]\ : AO1
      port map(A => \WR_XFER_TYPE[7]_net_1\, B => N_398, C => 
        \N_WR_USB_ADBUS_0_iv_0[7]\, Y => 
        \N_WR_USB_ADBUS_0_iv_2[7]\);
    
    \REG_STATE_0_RNIG1T21[1]\ : OAI1
      port map(A => \REG_STATE_0[2]_net_1\, B => 
        \REG_STATE_0[1]_net_1\, C => \USB_TXE_B\, Y => N_274);
    
    \SM_BANK_SEL_RNIJPL6[4]\ : NOR2
      port map(A => \SM_BANK_SEL[4]_net_1\, B => 
        \SM_BANK_SEL[21]_net_1\, Y => N_199);
    
    \RD_USB_ADBUS_RNI906B1[4]\ : NOR2
      port map(A => \RD_USB_ADBUS[4]_net_1\, B => N_282, Y => 
        \REG_STATE_ns_i_i_a5_1_1_0[2]\);
    
    \ELINK_DINA_6[5]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[5]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_16, E => un1_SM_BANK_SEL_10, Q => 
        \ELINK_DINA_6[5]_net_1\);
    
    \ELINK_ADDRA_9[0]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[0]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_10, E => un1_SM_BANK_SEL_9, Q => 
        \ELINK_ADDRA_9[0]_net_1\);
    
    \ELINK_ADDRA_1[2]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[2]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_20, E => un1_SM_BANK_SEL_19, Q => 
        \ELINK_ADDRA_1[2]_net_1\);
    
    \WR_USB_ADBUS_RNO_9[2]\ : OR3
      port map(A => \ELINK_DOUTA_5_m[2]\, B => 
        \ELINK_DOUTA_4_m[2]\, C => \N_WR_USB_ADBUS_0_iv_8[2]\, Y
         => \N_WR_USB_ADBUS_0_iv_18[2]\);
    
    \WR_USB_ADBUS_RNO_12[4]\ : NOR2B
      port map(A => \ELINK_DOUTA_11[4]\, B => un1_SM_BANK_SEL_26, 
        Y => \ELINK_DOUTA_11_m[4]\);
    
    \ELINK_ADDRA_19[5]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[5]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_13, E => un1_SM_BANK_SEL_11, Q => 
        \ELINK_ADDRA_19[5]_net_1\);
    
    TFC_BLKA : DFN1E0P0
      port map(D => N_TFC_BLKA, CLK => CLK60MHZ, PRE => 
        P_USB_MASTER_EN_c_13, E => N_142, Q => \TFC_BLKA\);
    
    \ELINK_DINA_8[4]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[4]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_18, E => un1_SM_BANK_SEL_21, Q => 
        \ELINK_DINA_8[4]_net_1\);
    
    \REG_STATE_RNI4VN31[4]\ : NOR2B
      port map(A => N_1499_2_i_0, B => \REG_STATE[4]_net_1\, Y
         => N_2537_1);
    
    \REG_ADDR[1]\ : DFN1E1C0
      port map(D => REG_ADDR_n1, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_10, E => REG_ADDRe, Q => 
        \REG_ADDR[1]_net_1\);
    
    \WR_USB_ADBUS[3]\ : DFN1E0C0
      port map(D => \N_WR_USB_ADBUS[3]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_15, E => un1_REG_STATE_26, Q => 
        \WR_USB_ADBUS[3]_net_1\);
    
    USB_TXE_B_RNIVDKA6 : AO1B
      port map(A => \REG_STATE_ns_i_a2_0_0_2[5]\, B => 
        \REG_STATE_ns_i_a2_4_2[5]\, C => N_1404_8, Y => 
        \REG_STATE_ns_i_a2_0_0[5]\);
    
    \REG_STATE_0[2]\ : DFN1C0
      port map(D => \REG_STATE_RNIVPG2K2[2]_net_1\, CLK => 
        CLK60MHZ, CLR => P_USB_MASTER_EN_c_22_0, Q => 
        \REG_STATE_0[2]_net_1\);
    
    \ELINK_DINA_12[7]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[7]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_12, E => un1_SM_BANK_SEL_7, Q => 
        \ELINK_DINA_12[7]_net_1\);
    
    \RD_USB_ADBUS_RNIEQBG1_0[7]\ : NOR3A
      port map(A => N_310, B => N_1700, C => 
        \RD_USB_ADBUS[7]_net_1\, Y => N_489);
    
    \WR_XFER_TYPE_RNI5LLM2[0]\ : NOR3C
      port map(A => N_1404_6, B => REG_STATE_tr72_6_0, C => 
        REG_STATE_tr72_6_1, Y => REG_STATE_tr72_6_3);
    
    \ELINK_ADDRA_9[4]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[4]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_10, E => un1_SM_BANK_SEL_9, Q => 
        \ELINK_ADDRA_9[4]_net_1\);
    
    \REG_ADDR_RNIHKJB1[3]\ : NOR3C
      port map(A => N_1398_i_0_a2_1, B => N_1398_i_0_a2_0, C => 
        N_491, Y => N_1398_i_0_a2_3);
    
    \ELINK_DINA_0[3]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[3]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_5, E => un1_SM_BANK_SEL_6, Q => 
        \ELINK_DINA_0[3]_net_1\);
    
    \ELINK_DINA_13[7]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[7]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_14, E => un1_SM_BANK_SEL_2, Q => 
        \ELINK_DINA_13[7]_net_1\);
    
    \REG_STATE_RNI2KQN_1[1]\ : NOR2
      port map(A => \REG_STATE[1]_net_1\, B => 
        \REG_STATE[5]_net_1\, Y => N_1499_2_i_0);
    
    \ELINK_BLKA[0]\ : DFN1E0P0
      port map(D => \N_ELINK_BLKA_0_iv[0]\, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_19, E => \SM_BANK_SEL_0[20]_net_1\, 
        Q => \ELINK_BLKA[0]_net_1\);
    
    \ELINK_ADDRA_7[1]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[1]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_5, E => un1_SM_BANK_SEL_12, Q => 
        \ELINK_ADDRA_7[1]_net_1\);
    
    \WR_USB_ADBUS_RNO_27[4]\ : NOR2B
      port map(A => \ELINK_DOUTA_19[4]\, B => un1_SM_BANK_SEL_41, 
        Y => \ELINK_DOUTA_19_m[4]\);
    
    \SM_BANK_SEL_RNI8QSA2[21]\ : OR2A
      port map(A => un1_USB_RXF_B_m, B => \SM_BANK_SEL[21]_net_1\, 
        Y => N_206);
    
    \ELINK_ADDRA_10[6]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[6]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_22, E => un1_SM_BANK_SEL_20, Q => 
        \ELINK_ADDRA_10[6]_net_1\);
    
    USB_TXE_B_RNIL2OI : OR2B
      port map(A => \USB_TXE_B\, B => \REG_STATE[4]_net_1\, Y => 
        N_339);
    
    \SM_BANK_SEL_RNIAS63[12]\ : OR3
      port map(A => \SM_BANK_SEL[13]_net_1\, B => 
        \SM_BANK_SEL[12]_net_1\, C => N_622_3, Y => 
        \N_ELINK_RWA_15_1[8]\);
    
    \ELINK_BLKA_RNO_0[3]\ : OA1B
      port map(A => N_616_16, B => \N_ELINK_RWA_3[3]\, C => 
        \ELINK_BLKA[3]_net_1\, Y => \ELINK_BLKA_i_m[3]\);
    
    \WR_USB_ADBUS_RNO_27[2]\ : NOR2B
      port map(A => \ELINK_DOUTA_9[2]\, B => un1_SM_BANK_SEL_42, 
        Y => \ELINK_DOUTA_9_m[2]\);
    
    \WR_USB_ADBUS_RNO_20[7]\ : NOR2A
      port map(A => \TFC_DOUTA[7]\, B => N_243, Y => 
        \TFC_DOUTA_m[7]\);
    
    USB_TXE_B_RNIKJIA1 : OR2B
      port map(A => N_339, B => N_312, Y => 
        \REG_STATE_ns_i_1_tz_1[3]\);
    
    \REG_STATE_RNI59LF1[1]\ : OR2A
      port map(A => N_1499_2_i_0, B => N_1726, Y => 
        REG_STATE_s22_i_0);
    
    \TFC_STRT_ADDR[0]\ : DFN1E1C0
      port map(D => \TFC_STRT_ADDR_T[0]_net_1\, CLK => CLK60MHZ, 
        CLR => P_USB_MASTER_EN_c_13, E => \REG_STATE_d_0[30]\, Q
         => \TFC_STRT_ADDR[0]_net_1\);
    
    \ELINK_BLKA_RNO_0[4]\ : OA1B
      port map(A => N_616_16, B => \N_ELINK_RWA_1[4]\, C => 
        \ELINK_BLKA[4]_net_1\, Y => \ELINK_BLKA_i_m[4]\);
    
    \WR_USB_ADBUS_RNO_22[3]\ : AO1
      port map(A => \ELINK_DOUTA_15[3]\, B => un1_SM_BANK_SEL_24, 
        C => \ELINK_DOUTA_0_m[3]\, Y => 
        \N_WR_USB_ADBUS_0_iv_8[3]\);
    
    \REG_STATE_ns_i_i_o2_1_RNO_1[0]\ : OA1B
      port map(A => N_437, B => N_436, C => 
        \REG_STATE_0[1]_net_1\, Y => N_441);
    
    U114_PATT_ELINK_BLK : DPRT_512X9_SRAM_14
      port map(ELINK_RWA_0 => \ELINK_RWA[14]_net_1\, 
        ELK_RX_SER_WORD_14(7) => ELK_RX_SER_WORD_14(7), 
        ELK_RX_SER_WORD_14(6) => ELK_RX_SER_WORD_14(6), 
        ELK_RX_SER_WORD_14(5) => ELK_RX_SER_WORD_14(5), 
        ELK_RX_SER_WORD_14(4) => ELK_RX_SER_WORD_14(4), 
        ELK_RX_SER_WORD_14(3) => ELK_RX_SER_WORD_14(3), 
        ELK_RX_SER_WORD_14(2) => ELK_RX_SER_WORD_14(2), 
        ELK_RX_SER_WORD_14(1) => ELK_RX_SER_WORD_14(1), 
        ELK_RX_SER_WORD_14(0) => ELK_RX_SER_WORD_14(0), 
        ELINK_DINA_14(7) => \ELINK_DINA_14[7]_net_1\, 
        ELINK_DINA_14(6) => \ELINK_DINA_14[6]_net_1\, 
        ELINK_DINA_14(5) => \ELINK_DINA_14[5]_net_1\, 
        ELINK_DINA_14(4) => \ELINK_DINA_14[4]_net_1\, 
        ELINK_DINA_14(3) => \ELINK_DINA_14[3]_net_1\, 
        ELINK_DINA_14(2) => \ELINK_DINA_14[2]_net_1\, 
        ELINK_DINA_14(1) => \ELINK_DINA_14[1]_net_1\, 
        ELINK_DINA_14(0) => \ELINK_DINA_14[0]_net_1\, 
        ELINK_BLKA_0 => \ELINK_BLKA[14]_net_1\, ELKS_ADDRB_0_d0
         => ELKS_ADDRB(0), ELKS_ADDRB_1 => ELKS_ADDRB(1), 
        ELKS_ADDRB_3 => ELKS_ADDRB(3), ELKS_ADDRB_5 => 
        ELKS_ADDRB(5), ELKS_ADDRB_7 => ELKS_ADDRB(7), 
        ELKS_ADDRB_0_0 => ELKS_ADDRB_0_0, ELKS_ADDRB_0_2 => 
        ELKS_ADDRB_0_2, ELKS_ADDRB_0_4 => ELKS_ADDRB_0_4, 
        ELINK_ADDRA_14(7) => \ELINK_ADDRA_14[7]_net_1\, 
        ELINK_ADDRA_14(6) => \ELINK_ADDRA_14[6]_net_1\, 
        ELINK_ADDRA_14(5) => \ELINK_ADDRA_14[5]_net_1\, 
        ELINK_ADDRA_14(4) => \ELINK_ADDRA_14[4]_net_1\, 
        ELINK_ADDRA_14(3) => \ELINK_ADDRA_14[3]_net_1\, 
        ELINK_ADDRA_14(2) => \ELINK_ADDRA_14[2]_net_1\, 
        ELINK_ADDRA_14(1) => \ELINK_ADDRA_14[1]_net_1\, 
        ELINK_ADDRA_14(0) => \ELINK_ADDRA_14[0]_net_1\, 
        PATT_ELK_DAT_14(7) => PATT_ELK_DAT_14(7), 
        PATT_ELK_DAT_14(6) => PATT_ELK_DAT_14(6), 
        PATT_ELK_DAT_14(5) => PATT_ELK_DAT_14(5), 
        PATT_ELK_DAT_14(4) => PATT_ELK_DAT_14(4), 
        PATT_ELK_DAT_14(3) => PATT_ELK_DAT_14(3), 
        PATT_ELK_DAT_14(2) => PATT_ELK_DAT_14(2), 
        PATT_ELK_DAT_14(1) => PATT_ELK_DAT_14(1), 
        PATT_ELK_DAT_14(0) => PATT_ELK_DAT_14(0), 
        ELINK_DOUTA_14(7) => \ELINK_DOUTA_14[7]\, 
        ELINK_DOUTA_14(6) => \ELINK_DOUTA_14[6]\, 
        ELINK_DOUTA_14(5) => \ELINK_DOUTA_14[5]\, 
        ELINK_DOUTA_14(4) => \ELINK_DOUTA_14[4]\, 
        ELINK_DOUTA_14(3) => \ELINK_DOUTA_14[3]\, 
        ELINK_DOUTA_14(2) => \ELINK_DOUTA_14[2]\, 
        ELINK_DOUTA_14(1) => \ELINK_DOUTA_14[1]\, 
        ELINK_DOUTA_14(0) => \ELINK_DOUTA_14[0]\, ELKS_RWB => 
        ELKS_RWB, P_USB_MASTER_EN_c_0 => P_USB_MASTER_EN_c_0, 
        CLK_40M_GL => CLK_40M_GL, CLK60MHZ => CLK60MHZ, 
        ELKS_RAM_BLKB_EN => ELKS_RAM_BLKB_EN);
    
    \WR_USB_ADBUS_RNO_12[7]\ : NOR2B
      port map(A => \ELINK_DOUTA_2[7]\, B => un1_SM_BANK_SEL_32, 
        Y => \ELINK_DOUTA_2_m[7]\);
    
    REG_STATE_s23_i : OR2
      port map(A => N_1705, B => \REG_STATE_s23_i_2\, Y => N_1501);
    
    \TFC_STRT_ADDR[1]\ : DFN1E1C0
      port map(D => \TFC_STRT_ADDR_T[1]_net_1\, CLK => CLK60MHZ, 
        CLR => P_USB_MASTER_EN_c_13, E => \REG_STATE_d_0[30]\, Q
         => \TFC_STRT_ADDR[1]_net_1\);
    
    \ELINK_ADDRA_10[0]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[0]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_21, E => un1_SM_BANK_SEL_20, Q => 
        \ELINK_ADDRA_10[0]_net_1\);
    
    \SM_BANK_SEL[18]\ : DFN1E1C0
      port map(D => N_1838, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_1_0, E => un1_REG_STATE_30, Q => 
        \SM_BANK_SEL[18]_net_1\);
    
    \WR_USB_ADBUS_RNO_22[0]\ : NOR2B
      port map(A => \ELINK_DOUTA_16[0]\, B => un1_SM_BANK_SEL_39, 
        Y => \ELINK_DOUTA_16_m[0]\);
    
    \ELINK_ADDRA_14[1]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[1]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_5, E => un1_SM_BANK_SEL_1, Q => 
        \ELINK_ADDRA_14[1]_net_1\);
    
    \WR_USB_ADBUS_RNO[0]\ : OR3
      port map(A => \N_WR_USB_ADBUS_0_iv_24[0]\, B => 
        \N_WR_USB_ADBUS_0_iv_23[0]\, C => 
        \N_WR_USB_ADBUS_0_iv_25[0]\, Y => \N_WR_USB_ADBUS[0]\);
    
    \REG_STATE_0_RNI21TJ1[5]\ : AOI1B
      port map(A => N_287, B => \REG_STATE_0[4]_net_1\, C => 
        \REG_STATE_0[5]_net_1\, Y => \REG_STATE_ns_i_a4_0_0[3]\);
    
    \ELINK_ADDRA_19[2]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[2]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_13, E => un1_SM_BANK_SEL_11, Q => 
        \ELINK_ADDRA_19[2]_net_1\);
    
    \REG_ADDR_RNIVAHE[8]\ : NOR2A
      port map(A => \REG_ADDR[7]_net_1\, B => \REG_ADDR[8]_net_1\, 
        Y => N_1398_i_0_a2_0);
    
    \ELINK_RWA_RNO[10]\ : AOI1
      port map(A => \SM_BANK_SEL[9]_net_1\, B => un1_USB_RXF_B_m, 
        C => \ELINK_RWA_i_m[10]\, Y => \N_ELINK_RWA_0_iv[10]\);
    
    \WR_USB_ADBUS_RNO_28[4]\ : AO1
      port map(A => \WR_XFER_TYPE[4]_net_1\, B => N_398, C => 
        \ELINKS_STOP_ADDR_m[4]\, Y => \N_WR_USB_ADBUS_0_iv_3[4]\);
    
    \WR_USB_ADBUS_RNO_15[3]\ : NOR2B
      port map(A => \ELINK_DOUTA_18[3]\, B => un1_SM_BANK_SEL_25, 
        Y => \ELINK_DOUTA_18_m[3]\);
    
    ELK_N_ACTIVE_RNIF389 : OR2A
      port map(A => \ELK_N_ACTIVE\, B => \USB_TXE_B\, Y => 
        \REG_STATE_ns_i_a2_4_0[5]\);
    
    \ELINK_DINA_8[5]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[5]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_18, E => un1_SM_BANK_SEL_21, Q => 
        \ELINK_DINA_8[5]_net_1\);
    
    \REG_STATE_RNI74ED2[2]\ : NOR3B
      port map(A => \REG_STATE_ns_i_a4_7_0[4]\, B => N_1499_2_i_0, 
        C => N_257, Y => N_2570);
    
    \REG_STATE_RNI3UN31_0[3]\ : NOR2A
      port map(A => N_1499_2_i_0, B => \REG_STATE[3]_net_1\, Y
         => N_2622);
    
    \ELINK_RWA_RNO_0[3]\ : OA1B
      port map(A => N_616_16, B => \N_ELINK_RWA_3[3]\, C => 
        \ELINK_RWA[3]_net_1\, Y => \ELINK_RWA_i_m[3]\);
    
    \WR_USB_ADBUS_RNO_30[6]\ : NOR2B
      port map(A => \ELINK_DOUTA_15[6]\, B => un1_SM_BANK_SEL_24, 
        Y => \ELINK_DOUTA_15_m[6]\);
    
    \ELINK_BLKA_RNO[17]\ : OA1C
      port map(A => N_131, B => \ELINK_BLKA[17]_net_1\, C => 
        X_BLKA_i_m_16, Y => \N_ELINK_BLKA_0_iv[17]\);
    
    \ELINK_ADDRA_11[3]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[3]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_2, E => un1_SM_BANK_SEL_16, Q => 
        \ELINK_ADDRA_11[3]_net_1\);
    
    \WR_USB_ADBUS_RNO_31[2]\ : NOR3B
      port map(A => N_1730_i, B => \ELINKS_STOP_ADDR[2]_net_1\, C
         => N_1726, Y => \ELINKS_STOP_ADDR_m[2]\);
    
    \ELINK_DINA_12[5]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[5]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_12, E => un1_SM_BANK_SEL_7, Q => 
        \ELINK_DINA_12[5]_net_1\);
    
    \ELINK_ADDRA_13[7]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[7]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_3, E => un1_SM_BANK_SEL_2, Q => 
        \ELINK_ADDRA_13[7]_net_1\);
    
    \WR_USB_ADBUS_RNO_24[6]\ : NOR2B
      port map(A => \ELINK_DOUTA_14[6]\, B => un1_SM_BANK_SEL_23, 
        Y => \ELINK_DOUTA_14_m[6]\);
    
    \WR_USB_ADBUS_RNO_2[0]\ : OR3
      port map(A => \N_WR_USB_ADBUS_0_iv_14[0]\, B => 
        \N_WR_USB_ADBUS_0_iv_13[0]\, C => 
        \N_WR_USB_ADBUS_0_iv_22[0]\, Y => 
        \N_WR_USB_ADBUS_0_iv_25[0]\);
    
    \SM_BANK_SEL_RNI69HH[5]\ : NOR2A
      port map(A => N_462, B => \SM_BANK_SEL[5]_net_1\, Y => 
        \N_ELINK_RWA_0_iv_0_o2_i_a5_0[13]\);
    
    \RD_USB_ADBUS_RNI91Q57[6]\ : OR3
      port map(A => N_1886, B => N_1887, C => N_1911, Y => N_1756);
    
    \WR_USB_ADBUS_RNO_18[2]\ : AO1A
      port map(A => N_1497, B => \TFC_STRT_ADDR[2]_net_1\, C => 
        \N_WR_USB_ADBUS_0_iv_2[2]\, Y => 
        \N_WR_USB_ADBUS_0_iv_4[2]\);
    
    un1_N_WR_USB_ADBUS_0_sqmuxa_i_0 : OR2A
      port map(A => \SM_BANK_SEL[20]_net_1\, B => \USB_TXE_B\, Y
         => \un1_N_WR_USB_ADBUS_0_sqmuxa_i_0\);
    
    \REG_STATE_ns_i_i_o2_1_RNO_8[0]\ : NOR2B
      port map(A => \REG_STATE[5]_net_1\, B => N_1359_1, Y => 
        \REG_STATE_ns_i_i_a2_9_0[0]\);
    
    \ELINK_DINA_12[0]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[0]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_12, E => un1_SM_BANK_SEL_7, Q => 
        \ELINK_DINA_12[0]_net_1\);
    
    \ELINK_DINA_16[1]\ : DFN1E0C0
      port map(D => \N_TFC_DINA[1]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_18, E => N_200, Q => 
        \ELINK_DINA_16[1]_net_1\);
    
    \ELINK_RWA_RNO[7]\ : AOI1
      port map(A => \SM_BANK_SEL[12]_net_1\, B => un1_USB_RXF_B_m, 
        C => \ELINK_RWA_i_m[7]\, Y => \N_ELINK_RWA_0_iv[7]\);
    
    \WR_USB_ADBUS_RNO_13[5]\ : NOR2B
      port map(A => \ELINK_DOUTA_1[5]\, B => un1_SM_BANK_SEL_36, 
        Y => \ELINK_DOUTA_1_m[5]\);
    
    \ELINK_ADDRA_16[2]\ : DFN1E0C0
      port map(D => \N_TFC_ADDRA[2]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_8, E => N_200, Q => 
        \ELINK_ADDRA_16[2]_net_1\);
    
    \ELINK_BLKA_RNO_0[19]\ : NOR2B
      port map(A => \SM_BANK_SEL[0]_net_1\, B => X_BLKA_i, Y => 
        X_BLKA_i_m_18);
    
    \RD_USB_ADBUS_RNIVNN03[5]\ : OR2
      port map(A => N_1893, B => N_1698, Y => N_1728);
    
    \WR_XFER_TYPE_RNO_0[1]\ : NOR3A
      port map(A => N_1736, B => \RD_USB_ADBUS[1]_net_1\, C => 
        N_1702, Y => N_1819);
    
    \RD_USB_ADBUS_RNISIOG3[4]\ : OR2
      port map(A => N_1702, B => N_293, Y => N_1716);
    
    USB_RXF_B_RNIJ4A61 : NOR2
      port map(A => N_268, B => \USB_RXF_B\, Y => N_446);
    
    \WR_USB_ADBUS_RNO_21[1]\ : NOR2B
      port map(A => \ELINK_DOUTA_19[1]\, B => un1_SM_BANK_SEL_41, 
        Y => \ELINK_DOUTA_19_m[1]\);
    
    \RD_USB_ADBUS_RNIQEIK2[5]\ : NOR2A
      port map(A => \RD_USB_ADBUS[5]_net_1\, B => N_206, Y => 
        \N_TFC_DINA[5]\);
    
    \WR_USB_ADBUS_RNO_13[3]\ : NOR2B
      port map(A => \ELINK_DOUTA_1[3]\, B => un1_SM_BANK_SEL_36, 
        Y => \ELINK_DOUTA_1_m[3]\);
    
    \WR_USB_ADBUS_RNO_23[4]\ : NOR2B
      port map(A => \ELINK_DOUTA_15[4]\, B => un1_SM_BANK_SEL_24, 
        Y => \ELINK_DOUTA_15_m[4]\);
    
    \REG_STATE_RNI4MQN[5]\ : NOR2
      port map(A => \REG_STATE[3]_net_1\, B => 
        \REG_STATE[5]_net_1\, Y => N_2526_1);
    
    \RD_USB_ADBUS_RNIMMEN4[5]\ : OA1B
      port map(A => \RD_USB_ADBUS[5]_net_1\, B => N_1881, C => 
        N_1717, Y => N_1823);
    
    \ELINK_RWA_RNO_0[8]\ : OA1B
      port map(A => N_616_16, B => \N_ELINK_RWA_0[8]\, C => 
        \ELINK_RWA[8]_net_1\, Y => \ELINK_RWA_i_m[8]\);
    
    \SM_BANK_SEL[7]\ : DFN1E1C0
      port map(D => N_1842, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_7, E => un1_REG_STATE_30, Q => 
        \SM_BANK_SEL[7]_net_1\);
    
    \ELINK_BLKA_RNO_0[8]\ : OA1B
      port map(A => N_616_16, B => \N_ELINK_RWA_0[8]\, C => 
        \ELINK_BLKA[8]_net_1\, Y => \ELINK_BLKA_i_m[8]\);
    
    \RD_XFER_TYPE_RNIRON38_0[0]\ : NOR3B
      port map(A => N_480, B => N_1368_i_i_a5_0, C => N_273, Y
         => N_357);
    
    \ELINK_ADDRA_8[0]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[0]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_8, E => un1_SM_BANK_SEL_21, Q => 
        \ELINK_ADDRA_8[0]_net_1\);
    
    \RD_USB_ADBUS_RNIPDIK2[4]\ : NOR2A
      port map(A => \RD_USB_ADBUS[4]_net_1\, B => N_206, Y => 
        \N_TFC_DINA[4]\);
    
    \USB_RD_BI\ : DFN1E0P0
      port map(D => N_1673, CLK => CLK60MHZ, PRE => 
        P_USB_MASTER_EN_c_13, E => N_1675, Q => USB_RD_BI);
    
    un1_REG_STATE_2_i_RNO : OR2
      port map(A => N_1778, B => N_1739, Y => un1_REG_STATE_2_i_0);
    
    U117_PATT_ELINK_BLK : DPRT_512X9_SRAM_17
      port map(ELINK_RWA_0 => \ELINK_RWA[17]_net_1\, 
        ELK_RX_SER_WORD_17(7) => ELK_RX_SER_WORD_17(7), 
        ELK_RX_SER_WORD_17(6) => ELK_RX_SER_WORD_17(6), 
        ELK_RX_SER_WORD_17(5) => ELK_RX_SER_WORD_17(5), 
        ELK_RX_SER_WORD_17(4) => ELK_RX_SER_WORD_17(4), 
        ELK_RX_SER_WORD_17(3) => ELK_RX_SER_WORD_17(3), 
        ELK_RX_SER_WORD_17(2) => ELK_RX_SER_WORD_17(2), 
        ELK_RX_SER_WORD_17(1) => ELK_RX_SER_WORD_17(1), 
        ELK_RX_SER_WORD_17(0) => ELK_RX_SER_WORD_17(0), 
        ELINK_DINA_17(7) => \ELINK_DINA_17[7]_net_1\, 
        ELINK_DINA_17(6) => \ELINK_DINA_17[6]_net_1\, 
        ELINK_DINA_17(5) => \ELINK_DINA_17[5]_net_1\, 
        ELINK_DINA_17(4) => \ELINK_DINA_17[4]_net_1\, 
        ELINK_DINA_17(3) => \ELINK_DINA_17[3]_net_1\, 
        ELINK_DINA_17(2) => \ELINK_DINA_17[2]_net_1\, 
        ELINK_DINA_17(1) => \ELINK_DINA_17[1]_net_1\, 
        ELINK_DINA_17(0) => \ELINK_DINA_17[0]_net_1\, 
        ELINK_BLKA_0 => \ELINK_BLKA[17]_net_1\, ELKS_ADDRB(7) => 
        ELKS_ADDRB(7), ELKS_ADDRB(6) => ELKS_ADDRB(6), 
        ELKS_ADDRB(5) => ELKS_ADDRB(5), ELKS_ADDRB(4) => 
        ELKS_ADDRB(4), ELKS_ADDRB(3) => ELKS_ADDRB(3), 
        ELKS_ADDRB(2) => ELKS_ADDRB(2), ELKS_ADDRB(1) => 
        ELKS_ADDRB(1), ELKS_ADDRB(0) => ELKS_ADDRB(0), 
        ELINK_ADDRA_17(7) => \ELINK_ADDRA_17[7]_net_1\, 
        ELINK_ADDRA_17(6) => \ELINK_ADDRA_17[6]_net_1\, 
        ELINK_ADDRA_17(5) => \ELINK_ADDRA_17[5]_net_1\, 
        ELINK_ADDRA_17(4) => \ELINK_ADDRA_17[4]_net_1\, 
        ELINK_ADDRA_17(3) => \ELINK_ADDRA_17[3]_net_1\, 
        ELINK_ADDRA_17(2) => \ELINK_ADDRA_17[2]_net_1\, 
        ELINK_ADDRA_17(1) => \ELINK_ADDRA_17[1]_net_1\, 
        ELINK_ADDRA_17(0) => \ELINK_ADDRA_17[0]_net_1\, 
        PATT_ELK_DAT_17(7) => PATT_ELK_DAT_17(7), 
        PATT_ELK_DAT_17(6) => PATT_ELK_DAT_17(6), 
        PATT_ELK_DAT_17(5) => PATT_ELK_DAT_17(5), 
        PATT_ELK_DAT_17(4) => PATT_ELK_DAT_17(4), 
        PATT_ELK_DAT_17(3) => PATT_ELK_DAT_17(3), 
        PATT_ELK_DAT_17(2) => PATT_ELK_DAT_17(2), 
        PATT_ELK_DAT_17(1) => PATT_ELK_DAT_17(1), 
        PATT_ELK_DAT_17(0) => PATT_ELK_DAT_17(0), 
        ELINK_DOUTA_17(7) => \ELINK_DOUTA_17[7]\, 
        ELINK_DOUTA_17(6) => \ELINK_DOUTA_17[6]\, 
        ELINK_DOUTA_17(5) => \ELINK_DOUTA_17[5]\, 
        ELINK_DOUTA_17(4) => \ELINK_DOUTA_17[4]\, 
        ELINK_DOUTA_17(3) => \ELINK_DOUTA_17[3]\, 
        ELINK_DOUTA_17(2) => \ELINK_DOUTA_17[2]\, 
        ELINK_DOUTA_17(1) => \ELINK_DOUTA_17[1]\, 
        ELINK_DOUTA_17(0) => \ELINK_DOUTA_17[0]\, ELKS_RWB => 
        ELKS_RWB, P_USB_MASTER_EN_c_0 => P_USB_MASTER_EN_c_0, 
        CLK_40M_GL => CLK_40M_GL, CLK60MHZ => CLK60MHZ, 
        ELKS_RAM_BLKB_EN => ELKS_RAM_BLKB_EN);
    
    \ELINK_DINA_12[2]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[2]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_12, E => un1_SM_BANK_SEL_7, Q => 
        \ELINK_DINA_12[2]_net_1\);
    
    \ELINK_BLKA[11]\ : DFN1E0P0
      port map(D => \N_ELINK_BLKA_0_iv[11]\, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_20, E => \SM_BANK_SEL[20]_net_1\, Q
         => \ELINK_BLKA[11]_net_1\);
    
    \WR_USB_ADBUS_RNO_32[2]\ : NOR3B
      port map(A => N_1352_1, B => \OP_MODE[2]_net_1\, C => 
        REG_STATE_s20_i_0, Y => \OP_MODE_m[2]\);
    
    \CHKSUM_RNO[3]\ : NOR2A
      port map(A => \RD_USB_ADBUS[3]_net_1\, B => N_675, Y => 
        N_1587);
    
    \ELINK_ADDRA_7[5]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[5]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_6, E => un1_SM_BANK_SEL_12, Q => 
        \ELINK_ADDRA_7[5]_net_1\);
    
    \REG_STATE_RNIVGQN_0[0]\ : OR2A
      port map(A => \REG_STATE[0]_net_1\, B => 
        \REG_STATE[3]_net_1\, Y => N_312);
    
    \ELINK_DINA_6[0]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[0]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_16, E => un1_SM_BANK_SEL_10, Q => 
        \ELINK_DINA_6[0]_net_1\);
    
    \WR_USB_ADBUS_RNO_4[6]\ : AO1
      port map(A => \ELINK_DOUTA_7[6]\, B => un1_SM_BANK_SEL_37, 
        C => \ELINK_DOUTA_16_m[6]\, Y => 
        \N_WR_USB_ADBUS_0_iv_8[6]\);
    
    \WR_USB_ADBUS_RNO_26[4]\ : AO1
      port map(A => \ELINK_DOUTA_2[4]\, B => un1_SM_BANK_SEL_32, 
        C => \ELINK_DOUTA_18_m[4]\, Y => 
        \N_WR_USB_ADBUS_0_iv_16[4]\);
    
    USB_WR_BI_RNO : OR3
      port map(A => N_1779, B => un1_REG_STATE_28_0_0, C => N_675, 
        Y => un1_REG_STATE_28);
    
    U4D_REGCROSS : CLK60M_TO_40M_4_2
      port map(ELINKS_STOP_ADDR(7) => \ELINKS_STOP_ADDR[7]_net_1\, 
        ELINKS_STOP_ADDR(6) => \ELINKS_STOP_ADDR[6]_net_1\, 
        ELINKS_STOP_ADDR(5) => \ELINKS_STOP_ADDR[5]_net_1\, 
        ELINKS_STOP_ADDR(4) => \ELINKS_STOP_ADDR[4]_net_1\, 
        ELINKS_STOP_ADDR(3) => \ELINKS_STOP_ADDR[3]_net_1\, 
        ELINKS_STOP_ADDR(2) => \ELINKS_STOP_ADDR[2]_net_1\, 
        ELINKS_STOP_ADDR(1) => \ELINKS_STOP_ADDR[1]_net_1\, 
        ELINKS_STOP_ADDR(0) => \ELINKS_STOP_ADDR[0]_net_1\, 
        ELKS_STOP_ADDR(7) => ELKS_STOP_ADDR(7), ELKS_STOP_ADDR(6)
         => ELKS_STOP_ADDR(6), ELKS_STOP_ADDR(5) => 
        ELKS_STOP_ADDR(5), ELKS_STOP_ADDR(4) => ELKS_STOP_ADDR(4), 
        ELKS_STOP_ADDR(3) => ELKS_STOP_ADDR(3), ELKS_STOP_ADDR(2)
         => ELKS_STOP_ADDR(2), ELKS_STOP_ADDR(1) => 
        ELKS_STOP_ADDR(1), ELKS_STOP_ADDR(0) => ELKS_STOP_ADDR(0), 
        P_MASTER_POR_B_c_26 => P_MASTER_POR_B_c_26, 
        P_MASTER_POR_B_c_30 => P_MASTER_POR_B_c_30, 
        P_MASTER_POR_B_c_3 => P_MASTER_POR_B_c_3, 
        P_MASTER_POR_B_c_25 => P_MASTER_POR_B_c_25, CLK_40M_GL
         => CLK_40M_GL);
    
    \REG_STATE_ns_i_8_tz_1_RNI26A381[4]\ : NOR2B
      port map(A => N_2597, B => \REG_STATE_ns_i_8_tz[4]\, Y => 
        \REG_STATE_ns_i_8[4]\);
    
    \TFC_STRT_ADDR_T[0]\ : DFN1E1C0
      port map(D => \RD_USB_ADBUS[0]_net_1\, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_4, E => N_TFC_STRT_ADDR_T_0_sqmuxa, 
        Q => \TFC_STRT_ADDR_T[0]_net_1\);
    
    \ELINK_DINA_16[0]\ : DFN1E0C0
      port map(D => \N_TFC_DINA[0]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_18, E => N_200, Q => 
        \ELINK_DINA_16[0]_net_1\);
    
    \RD_USB_ADBUS_RNI575O[6]\ : OR2
      port map(A => \RD_USB_ADBUS[6]_net_1\, B => \USB_RXF_B\, Y
         => N_1695);
    
    \ELINK_RWA_RNO_0[9]\ : NOR2B
      port map(A => \SM_BANK_SEL[10]_net_1\, B => un1_USB_RXF_B_m, 
        Y => N_182);
    
    \ELINK_ADDRA_10[2]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[2]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_22, E => un1_SM_BANK_SEL_20, Q => 
        \ELINK_ADDRA_10[2]_net_1\);
    
    \WR_USB_ADBUS_RNO_5[6]\ : OR3
      port map(A => \ELINK_DOUTA_8_m[6]\, B => 
        \ELINK_DOUTA_19_m[6]\, C => \N_WR_USB_ADBUS_0_iv_11[6]\, 
        Y => \N_WR_USB_ADBUS_0_iv_19[6]\);
    
    \WR_USB_ADBUS_RNO_6[5]\ : OR3
      port map(A => \N_WR_USB_ADBUS_0_iv_3[5]\, B => 
        \N_WR_USB_ADBUS_0_iv_2[5]\, C => 
        \N_WR_USB_ADBUS_0_iv_4[5]\, Y => 
        \N_WR_USB_ADBUS_0_iv_6[5]\);
    
    \REG_STATE_ns_i_8_tz_1_RNILKP34[4]\ : OR3
      port map(A => N_457, B => N_456, C => 
        \REG_STATE_ns_i_8_tz_1[4]_net_1\, Y => 
        \REG_STATE_ns_i_8_tz[4]\);
    
    \ELINK_ADDRA_1[7]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[7]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_20, E => un1_SM_BANK_SEL_19, Q => 
        \ELINK_ADDRA_1[7]_net_1\);
    
    \ELINKS_STRT_ADDR[7]\ : DFN1E1C0
      port map(D => \ELINKS_STRT_ADDR_T[7]_net_1\, CLK => 
        CLK60MHZ, CLR => P_USB_MASTER_EN_c_18, E => 
        \REG_STATE_d[30]\, Q => \ELINKS_STRT_ADDR[7]_net_1\);
    
    \CHKSUM_RNO[2]\ : NOR2A
      port map(A => \RD_USB_ADBUS[2]_net_1\, B => N_675, Y => 
        N_234);
    
    \WR_USB_ADBUS_RNO_12[5]\ : NOR2B
      port map(A => \ELINK_DOUTA_2[5]\, B => un1_SM_BANK_SEL_32, 
        Y => \ELINK_DOUTA_2_m[5]\);
    
    USB_TXE_B_RNICNL6Q : OA1
      port map(A => N_1278_tz, B => \REG_STATE_ns_i_a4_8_0[1]\, C
         => N_2587, Y => \REG_STATE_ns_i_3[1]\);
    
    USB_RXF_B_0_RNIGG3L1 : NOR3B
      port map(A => \REG_STATE_0[2]_net_1\, B => N_1690_i, C => 
        \USB_RXF_B_0\, Y => \REG_STATE_ns_i_a4_10_0[1]\);
    
    \REG_STATE_0_RNIICMT1[0]\ : NOR3C
      port map(A => N_292, B => \REG_STATE_0[0]_net_1\, C => 
        N_1499_2_i_0, Y => N_415);
    
    \ELINKS_STOP_ADDR_T[2]\ : DFN1E1C0
      port map(D => \RD_USB_ADBUS[2]_net_1\, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_7, E => 
        N_ELINKS_STOP_ADDR_T_0_sqmuxa, Q => 
        \ELINKS_STOP_ADDR_T[2]_net_1\);
    
    \WR_USB_ADBUS_RNO_16[1]\ : AO1
      port map(A => \ELINK_DOUTA_4[1]\, B => un1_SM_BANK_SEL_28, 
        C => \ELINK_DOUTA_5_m[1]\, Y => 
        \N_WR_USB_ADBUS_0_iv_12[1]\);
    
    \SM_BANK_SEL_RNIH37M1[10]\ : OR3B
      port map(A => N_477, B => N_143, C => \N_ELINK_RWA_0[10]\, 
        Y => \N_ELINK_RWA_2[10]\);
    
    \ELINK_DINA_0[5]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[5]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_5, E => un1_SM_BANK_SEL_6, Q => 
        \ELINK_DINA_0[5]_net_1\);
    
    \SM_BANK_SEL_RNIG11C2[6]\ : NOR3A
      port map(A => \SM_BANK_SEL[6]_net_1\, B => N_312_0, C => 
        N_1566_i_i_0, Y => un1_SM_BANK_SEL_29);
    
    \REG_STATE_ns_i_i_o2_6_1_RNO_0[0]\ : AO1A
      port map(A => N_1359_1, B => \REG_STATE_ns_i_i_a2_5_0[0]\, 
        C => N_452, Y => \REG_STATE_ns_i_i_o2_6_0[0]\);
    
    \SM_BANK_SEL_RNIBDMB[8]\ : NOR2
      port map(A => \SM_BANK_SEL[8]_net_1\, B => 
        \SM_BANK_SEL[7]_net_1\, Y => N_461);
    
    \WR_USB_ADBUS_RNO_5[0]\ : OR3
      port map(A => \ELINK_DOUTA_13_m[0]\, B => 
        \ELINK_DOUTA_12_m[0]\, C => \N_WR_USB_ADBUS_0_iv_12[0]\, 
        Y => \N_WR_USB_ADBUS_0_iv_20[0]\);
    
    \ELINK_DINA_5[5]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[5]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_14, E => un1_SM_BANK_SEL_15, Q => 
        \ELINK_DINA_5[5]_net_1\);
    
    \WR_USB_ADBUS_RNO_8[1]\ : OR3
      port map(A => \TFC_DOUTA_m[1]\, B => \ELINK_DOUTA_19_m[1]\, 
        C => \N_WR_USB_ADBUS_0_iv_8[1]\, Y => 
        \N_WR_USB_ADBUS_0_iv_18[1]\);
    
    \WR_USB_ADBUS_RNO_10[2]\ : OR3
      port map(A => \N_WR_USB_ADBUS_0_iv_5[2]\, B => 
        \N_WR_USB_ADBUS_0_iv_4[2]\, C => \ELINK_DOUTA_3_m[2]\, Y
         => \N_WR_USB_ADBUS_0_iv_17[2]\);
    
    \ELINK_ADDRA_16[3]\ : DFN1E0C0
      port map(D => \N_TFC_ADDRA[3]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_8, E => N_200, Q => 
        \ELINK_ADDRA_16[3]_net_1\);
    
    \WR_XFER_TYPE_RNO_2[1]\ : OA1C
      port map(A => N_1736, B => N_1702, C => 
        \WR_XFER_TYPE[1]_net_1\, Y => N_1820);
    
    \WR_XFER_TYPE_RNO_1[3]\ : NOR2A
      port map(A => N_1716, B => \WR_XFER_TYPE[3]_net_1\, Y => 
        N_1825);
    
    \RD_USB_ADBUS_RNI2CM61[4]\ : NOR3B
      port map(A => \RD_USB_ADBUS[5]_net_1\, B => 
        \RD_USB_ADBUS[4]_net_1\, C => N_1700, Y => 
        un1_N_ELK_N_ACTIVE_0_sqmuxa_15_0_a2_0_0);
    
    \WR_USB_ADBUS_RNO_17[7]\ : AO1A
      port map(A => N_1497, B => \TFC_STRT_ADDR[7]_net_1\, C => 
        \ELINKS_STOP_ADDR_m[7]\, Y => \N_WR_USB_ADBUS_0_iv_3[7]\);
    
    \ELINK_ADDRA_2[0]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[0]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_21, E => un1_SM_BANK_SEL_5, Q => 
        \ELINK_ADDRA_2[0]_net_1\);
    
    \ELINK_DINA_5[7]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[7]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_14, E => un1_SM_BANK_SEL_15, Q => 
        \ELINK_DINA_5[7]_net_1\);
    
    \ELINK_ADDRA_0[4]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[4]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_18, E => un1_SM_BANK_SEL_6, Q => 
        \ELINK_ADDRA_0[4]_net_1\);
    
    \WR_USB_ADBUS_RNO_19[3]\ : OR3A
      port map(A => N_1569, B => \ELINKS_STRT_ADDR_m[3]\, C => 
        \CHKSUM_m[3]\, Y => \N_WR_USB_ADBUS_0_iv_4[3]\);
    
    \ELINK_DINA_16[3]\ : DFN1E0C0
      port map(D => \N_TFC_DINA[3]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_18, E => N_200, Q => 
        \ELINK_DINA_16[3]_net_1\);
    
    \WR_USB_ADBUS_RNO_19[0]\ : AO1
      port map(A => \CHKSUM[0]_net_1\, B => un1_REG_STATE_4, C
         => \N_WR_USB_ADBUS_0_iv_3[0]\, Y => 
        \N_WR_USB_ADBUS_0_iv_5[0]\);
    
    USB_RXF_B_0_RNI0J4O4 : OA1C
      port map(A => N_1351_8, B => N_1398_i_0_0, C => 
        \USB_RXF_B_0\, Y => \REG_STATE_ns_i_i_a2_0[0]_net_1\);
    
    \REG_ADDR_RNIGHPL[1]\ : OR3
      port map(A => \REG_ADDR[1]_net_1\, B => \REG_ADDR[0]_net_1\, 
        C => \REG_ADDR[7]_net_1\, Y => REG_STATE_tr74_tz_tz_tz_4);
    
    \REG_STATE_RNIHK7Q2[0]\ : OA1
      port map(A => N_1713, B => N_1891, C => N_433_1, Y => 
        N_1905);
    
    \REG_STATE_RNI2KQN_0[1]\ : NOR2A
      port map(A => \REG_STATE[5]_net_1\, B => 
        \REG_STATE[1]_net_1\, Y => N_2602);
    
    \REG_ADDR_RNIMRCP[3]\ : NOR3B
      port map(A => N_261, B => \REG_ADDR[3]_net_1\, C => 
        \SM_BANK_SEL_0[21]_net_1\, Y => \N_TFC_ADDRA[3]\);
    
    \REG_STATE_0_RNIGJ3A1[3]\ : OR3C
      port map(A => \REG_STATE_0[2]_net_1\, B => 
        \REG_STATE_0[4]_net_1\, C => \REG_STATE_0[3]_net_1\, Y
         => REG_STATE_s20_i_0);
    
    \N_TFC_ADDRA_0_o2_RNO_4[7]\ : NOR3B
      port map(A => \REG_STATE_0[0]_net_1\, B => N_2600, C => 
        \REG_STATE_0[2]_net_1\, Y => \N_TFC_ADDRA_0_a2_1_1[7]\);
    
    \ELINK_ADDRA_4[7]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[7]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_2_0, E => un1_SM_BANK_SEL_8, Q => 
        \ELINK_ADDRA_4[7]_net_1\);
    
    \REG_STATE_ns_i_8_tz_0_RNO_0[4]\ : NOR3B
      port map(A => \REG_STATE_0[5]_net_1\, B => 
        \REG_STATE_0[3]_net_1\, C => \REG_STATE[2]_net_1\, Y => 
        \REG_STATE_ns_i_a4_5_1[4]\);
    
    USB_RXF_B_RNI1R5C2 : NOR3
      port map(A => N_1751, B => \USB_RXF_B\, C => N_1765, Y => 
        N_OP_MODE_T_0_sqmuxa);
    
    \TFC_STRT_ADDR_T[6]\ : DFN1E1C0
      port map(D => \RD_USB_ADBUS[6]_net_1\, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_5, E => N_TFC_STRT_ADDR_T_0_sqmuxa, 
        Q => \TFC_STRT_ADDR_T[6]_net_1\);
    
    \SM_BANK_SEL_RNO[18]\ : NOR3B
      port map(A => N_1882, B => N_1351_4, C => N_1700, Y => 
        N_1838);
    
    \RD_XFER_TYPE_RNO[4]\ : AO1
      port map(A => \RD_XFER_TYPE[4]_net_1\, B => N_1703, C => 
        N_1802, Y => \RD_XFER_TYPE_RNO[4]_net_1\);
    
    \ELINKS_STRT_ADDR[3]\ : DFN1E1C0
      port map(D => \ELINKS_STRT_ADDR_T[3]_net_1\, CLK => 
        CLK60MHZ, CLR => P_USB_MASTER_EN_c_17, E => 
        \REG_STATE_d[30]\, Q => \ELINKS_STRT_ADDR[3]_net_1\);
    
    \WR_USB_ADBUS_RNO_21[4]\ : NOR2B
      port map(A => \ELINK_DOUTA_3[4]\, B => un1_SM_BANK_SEL_43, 
        Y => \ELINK_DOUTA_3_m[4]\);
    
    USB_RXF_B_0_RNI0N432 : NOR2B
      port map(A => un1_REG_STATE_40_i_a2_3_0, B => N_1710_i_0, Y
         => N_1887);
    
    \SM_BANK_SEL_RNIULLS1[2]\ : OR3B
      port map(A => N_394, B => N_464, C => 
        \SM_BANK_SEL[2]_net_1\, Y => N_130);
    
    \ELINK_ADDRA_12[4]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[4]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_2_0, E => un1_SM_BANK_SEL_7, Q => 
        \ELINK_ADDRA_12[4]_net_1\);
    
    \SM_BANK_SEL_RNIKQL6[5]\ : OR2
      port map(A => \SM_BANK_SEL[5]_net_1\, B => 
        \SM_BANK_SEL[21]_net_1\, Y => un1_SM_BANK_SEL_1);
    
    USB_OE_BI_RNO_1 : NOR3B
      port map(A => N_1879_1, B => \USB_RXF_B\, C => N_1359_2, Y
         => N_1879);
    
    \REG_STATE_0_RNICF3A1[4]\ : NOR2A
      port map(A => N_2462, B => \REG_STATE_0[4]_net_1\, Y => 
        N_414_1);
    
    \SM_BANK_SEL[17]\ : DFN1E1C0
      port map(D => N_1851, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_1_0, E => un1_REG_STATE_30, Q => 
        \SM_BANK_SEL[17]_net_1\);
    
    \SM_BANK_SEL_RNI2NV62[17]\ : NOR3A
      port map(A => \SM_BANK_SEL[17]_net_1\, B => N_312_0, C => 
        N_1566_i_i_0, Y => un1_SM_BANK_SEL_32);
    
    \ELINK_RWA[7]\ : DFN1E0P0
      port map(D => \N_ELINK_RWA_0_iv[7]\, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_6, E => \SM_BANK_SEL_0[20]_net_1\, 
        Q => \ELINK_RWA[7]_net_1\);
    
    \TFC_STRT_ADDR_T[2]\ : DFN1E1C0
      port map(D => \RD_USB_ADBUS[2]_net_1\, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_4, E => N_TFC_STRT_ADDR_T_0_sqmuxa, 
        Q => \TFC_STRT_ADDR_T[2]_net_1\);
    
    \SM_BANK_SEL[11]\ : DFN1E1C0
      port map(D => N_1846, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_1_0, E => un1_REG_STATE_30, Q => 
        \SM_BANK_SEL[11]_net_1\);
    
    \WR_USB_ADBUS_RNO_21[7]\ : NOR2B
      port map(A => \ELINK_DOUTA_19[7]\, B => un1_SM_BANK_SEL_41, 
        Y => \ELINK_DOUTA_19_m[7]\);
    
    \REG_STATE_0_RNIF9MT1[1]\ : OR2
      port map(A => N_1765, B => N_1726, Y => N_1497);
    
    \WR_USB_ADBUS_RNO_15[5]\ : NOR2B
      port map(A => \ELINK_DOUTA_18[5]\, B => un1_SM_BANK_SEL_25, 
        Y => \ELINK_DOUTA_18_m[5]\);
    
    USB_RD_BI_RNO_1 : AO1A
      port map(A => N_1751, B => un1_REG_STATE_40_i_a2_0_0, C => 
        N_1877, Y => un1_REG_STATE_40_i_o2_0);
    
    \REG_STATE_RNIE3U12[5]\ : NOR2B
      port map(A => N_2526_1, B => N_1730_i, Y => N_1917);
    
    USB_TXE_B_RNIMCVT1 : OR3
      port map(A => \REG_STATE_ns_i_a2_0_0_0[5]\, B => 
        \USB_TXE_B\, C => N_252, Y => 
        \REG_STATE_ns_i_a2_0_0_2[5]\);
    
    REG_STATE_s20_i_o2_0_0_o2_0 : OR2B
      port map(A => \REG_STATE[4]_net_1\, B => 
        \REG_STATE[2]_net_1\, Y => N_1705);
    
    \REG_ADDR_RNIVNRI1[2]\ : NOR3C
      port map(A => REG_STATE_tr73_2, B => REG_STATE_tr73_1, C
         => REG_STATE_tr73_4, Y => REG_STATE_tr73_7);
    
    \ELINK_ADDRA_12[3]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[3]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_2_0, E => un1_SM_BANK_SEL_7, Q => 
        \ELINK_ADDRA_12[3]_net_1\);
    
    \WR_USB_ADBUS_RNO_18[5]\ : OR3
      port map(A => \OP_MODE_m[5]\, B => \TFC_STOP_ADDR_m[5]\, C
         => \WR_XFER_TYPE_m[5]\, Y => \N_WR_USB_ADBUS_0_iv_2[5]\);
    
    \WR_USB_ADBUS_RNO_16[6]\ : AO1
      port map(A => \ELINK_DOUTA_9[6]\, B => un1_SM_BANK_SEL_42, 
        C => \ELINK_DOUTA_10_m[6]\, Y => 
        \N_WR_USB_ADBUS_0_iv_11[6]\);
    
    U4B_REGCROSS : CLK60M_TO_40M_4_0
      port map(TFC_STOP_ADDR_0(7) => \TFC_STOP_ADDR[7]_net_1\, 
        TFC_STOP_ADDR_0(6) => \TFC_STOP_ADDR[6]_net_1\, 
        TFC_STOP_ADDR_0(5) => \TFC_STOP_ADDR[5]_net_1\, 
        TFC_STOP_ADDR_0(4) => \TFC_STOP_ADDR[4]_net_1\, 
        TFC_STOP_ADDR_0(3) => \TFC_STOP_ADDR[3]_net_1\, 
        TFC_STOP_ADDR_0(2) => \TFC_STOP_ADDR[2]_net_1\, 
        TFC_STOP_ADDR_0(1) => \TFC_STOP_ADDR[1]_net_1\, 
        TFC_STOP_ADDR_0(0) => \TFC_STOP_ADDR[0]_net_1\, 
        TFC_STOP_ADDR(7) => TFC_STOP_ADDR_0(7), TFC_STOP_ADDR(6)
         => TFC_STOP_ADDR_0(6), TFC_STOP_ADDR(5) => 
        TFC_STOP_ADDR_0(5), TFC_STOP_ADDR(4) => 
        TFC_STOP_ADDR_0(4), TFC_STOP_ADDR(3) => 
        TFC_STOP_ADDR_0(3), TFC_STOP_ADDR(2) => 
        TFC_STOP_ADDR_0(2), TFC_STOP_ADDR(1) => 
        TFC_STOP_ADDR_0(1), TFC_STOP_ADDR(0) => 
        TFC_STOP_ADDR_0(0), P_MASTER_POR_B_c_30 => 
        P_MASTER_POR_B_c_30, P_MASTER_POR_B_c_29 => 
        P_MASTER_POR_B_c_29, P_MASTER_POR_B_c_25 => 
        P_MASTER_POR_B_c_25, P_MASTER_POR_B_c_24_0 => 
        P_MASTER_POR_B_c_24_0, P_MASTER_POR_B_c_19 => 
        P_MASTER_POR_B_c_19, P_MASTER_POR_B_c_23 => 
        P_MASTER_POR_B_c_23, CLK_40M_GL => CLK_40M_GL);
    
    REG_STATE_s23_i_2_RNO_0 : OR2
      port map(A => \REG_STATE[0]_net_1\, B => 
        \REG_STATE[1]_net_1\, Y => REG_STATE_s23_i_0);
    
    \WR_USB_ADBUS_RNO_3[1]\ : AO1
      port map(A => \ELINK_DOUTA_17[1]\, B => un1_SM_BANK_SEL_40, 
        C => \ELINK_DOUTA_2_m[1]\, Y => 
        \N_WR_USB_ADBUS_0_iv_10[1]\);
    
    \ELINK_RWA_RNO_0[16]\ : AOI1
      port map(A => \N_ELINK_RWA_i_a2_0_a5_0[16]\, B => N_503, C
         => \ELINK_RWA[16]_net_1\, Y => \ELINK_RWA_i_m[16]\);
    
    \ELINK_RWA_RNO[8]\ : AOI1
      port map(A => \SM_BANK_SEL[11]_net_1\, B => un1_USB_RXF_B_m, 
        C => \ELINK_RWA_i_m[8]\, Y => \N_ELINK_RWA_0_iv[8]\);
    
    \RD_USB_ADBUS_RNI5LTB4[4]\ : OA1
      port map(A => N_488, B => N_489, C => 
        \REG_STATE_ns_i_i_a5_1_1_0[2]\, Y => 
        \REG_STATE_ns_i_i_a5_1[2]\);
    
    \WR_USB_ADBUS_RNO_31[3]\ : NOR2A
      port map(A => \TFC_STOP_ADDR[3]_net_1\, B => N_1501, Y => 
        \TFC_STOP_ADDR_m[3]\);
    
    \ELINK_ADDRA_19[0]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[0]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_13, E => un1_SM_BANK_SEL_11, Q => 
        \ELINK_ADDRA_19[0]_net_1\);
    
    \TFC_STOP_ADDR[6]\ : DFN1E1C0
      port map(D => \TFC_STOP_ADDR_T[6]_net_1\, CLK => CLK60MHZ, 
        CLR => P_USB_MASTER_EN_c_8, E => \REG_STATE_d_0[30]\, Q
         => \TFC_STOP_ADDR[6]_net_1\);
    
    \WR_USB_ADBUS_RNO_29[7]\ : NOR3B
      port map(A => N_1730_i, B => \ELINKS_STOP_ADDR[7]_net_1\, C
         => N_1726, Y => \ELINKS_STOP_ADDR_m[7]\);
    
    \ELINK_DINA_1[2]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[2]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_7, E => un1_SM_BANK_SEL_19, Q => 
        \ELINK_DINA_1[2]_net_1\);
    
    \ELINK_BLKA_RNO_0[14]\ : OA1B
      port map(A => N_624_15, B => \N_ELINK_RWA_3[14]\, C => 
        \ELINK_BLKA[14]_net_1\, Y => \ELINK_BLKA_i_m[14]\);
    
    \RD_USB_ADBUS[7]\ : DFN1C0
      port map(D => \N_RD_USB_ADBUS[7]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_22_0, Q => \RD_USB_ADBUS[7]_net_1\);
    
    \ELINKS_STRT_ADDR[0]\ : DFN1E1C0
      port map(D => \ELINKS_STRT_ADDR_T[0]_net_1\, CLK => 
        CLK60MHZ, CLR => P_USB_MASTER_EN_c_17, E => 
        \REG_STATE_d[30]\, Q => \ELINKS_STRT_ADDR[0]_net_1\);
    
    \RD_XFER_TYPE_RNITJ4J2[2]\ : OR3
      port map(A => N_1367_i_i_o2_0_1, B => N_1367_i_i_o2_0_0, C
         => N_1367_i_i_o2_0_2, Y => N_273);
    
    \RD_USB_ADBUS_RNIIEKR6[5]\ : AO1A
      port map(A => N_1697, B => 
        un1_N_ELK_N_ACTIVE_2_sqmuxa_0_a2_0_0, C => N_1860, Y => 
        un1_N_ELK_N_ACTIVE_2_sqmuxa);
    
    \WR_USB_ADBUS_RNO_32[4]\ : NOR3B
      port map(A => N_1352_1, B => \OP_MODE[4]_net_1\, C => 
        REG_STATE_s20_i_0, Y => \OP_MODE_m[4]\);
    
    \SM_BANK_SEL[16]\ : DFN1E1C0
      port map(D => N_1835, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_1_0, E => un1_REG_STATE_30, Q => 
        \SM_BANK_SEL[16]_net_1\);
    
    \ELINK_DINA_4[1]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[1]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_12, E => un1_SM_BANK_SEL_8, Q => 
        \ELINK_DINA_4[1]_net_1\);
    
    \ELINKS_STOP_ADDR_T[0]\ : DFN1E1C0
      port map(D => \RD_USB_ADBUS[0]_net_1\, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_7, E => 
        N_ELINKS_STOP_ADDR_T_0_sqmuxa, Q => 
        \ELINKS_STOP_ADDR_T[0]_net_1\);
    
    \ELINK_DINA_4[6]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[6]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_13, E => un1_SM_BANK_SEL_8, Q => 
        \ELINK_DINA_4[6]_net_1\);
    
    \ELINK_DINA_15[0]\ : DFN1E0C0
      port map(D => \N_TFC_DINA[0]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_16, E => N_199, Q => 
        \ELINK_DINA_15[0]_net_1\);
    
    \WR_USB_ADBUS_RNO_26[0]\ : AO1
      port map(A => \ELINK_DOUTA_2[0]\, B => un1_SM_BANK_SEL_32, 
        C => \ELINK_DOUTA_18_m[0]\, Y => 
        \N_WR_USB_ADBUS_0_iv_16[0]\);
    
    \ELINK_ADDRA_14[6]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[6]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_5, E => un1_SM_BANK_SEL_1, Q => 
        \ELINK_ADDRA_14[6]_net_1\);
    
    USB_TXE_B_RNI75TNL2 : NOR3
      port map(A => \REG_STATE_ns_i_3[1]\, B => 
        \REG_STATE_ns_i_2[1]\, C => \REG_STATE_ns_i_4[1]\, Y => 
        \USB_TXE_B_RNI75TNL2\);
    
    \ELINK_DINA_14[6]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[6]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_16, E => un1_SM_BANK_SEL_1, Q => 
        \ELINK_DINA_14[6]_net_1\);
    
    \REG_ADDR_RNIPUCP[6]\ : NOR3B
      port map(A => N_261, B => \REG_ADDR[6]_net_1\, C => 
        \SM_BANK_SEL_0[21]_net_1\, Y => \N_TFC_ADDRA[6]\);
    
    \ELINK_BLKA_RNO_0[10]\ : OA1B
      port map(A => N_624_15, B => \N_ELINK_RWA_2[10]\, C => 
        \ELINK_BLKA[10]_net_1\, Y => \ELINK_BLKA_i_m[10]\);
    
    \WR_USB_ADBUS_RNO_7[6]\ : AO1A
      port map(A => N_243, B => \TFC_DOUTA[6]\, C => 
        \ELINK_DOUTA_4_m[6]\, Y => \N_WR_USB_ADBUS_0_iv_6[6]\);
    
    USB_WR_BI_RNO_1 : AO1B
      port map(A => N_1761_i, B => \REG_STATE_0[5]_net_1\, C => 
        N_1726, Y => un1_REG_STATE_28_0_0);
    
    \REG_ADDR_RNIBCPL[2]\ : NOR3C
      port map(A => \REG_ADDR[0]_net_1\, B => \REG_ADDR[1]_net_1\, 
        C => \REG_ADDR[2]_net_1\, Y => N_474);
    
    \ELINK_DINA_1[4]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[4]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_7, E => un1_SM_BANK_SEL_19, Q => 
        \ELINK_DINA_1[4]_net_1\);
    
    \RD_USB_ADBUS_RNIOCG11[6]\ : OR2A
      port map(A => N_1351_3, B => \RD_USB_ADBUS[6]_net_1\, Y => 
        N_282);
    
    \REG_STATE_RNI3UN31[3]\ : NOR2B
      port map(A => \REG_STATE[3]_net_1\, B => N_2600, Y => 
        \REG_STATE_ns_i_a4_7_0[1]\);
    
    \RD_XFER_TYPE[4]\ : DFN1C0
      port map(D => \RD_XFER_TYPE_RNO[4]_net_1\, CLK => CLK60MHZ, 
        CLR => P_USB_MASTER_EN_c, Q => \RD_XFER_TYPE[4]_net_1\);
    
    \SM_BANK_SEL_RNIIOL6[3]\ : NOR2
      port map(A => \SM_BANK_SEL[3]_net_1\, B => 
        \SM_BANK_SEL[21]_net_1\, Y => N_200);
    
    \ELINK_DINA_8[7]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[7]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_18, E => un1_SM_BANK_SEL_21, Q => 
        \ELINK_DINA_8[7]_net_1\);
    
    \WR_USB_ADBUS_RNO_25[6]\ : NOR2B
      port map(A => \ELINK_DOUTA_1[6]\, B => un1_SM_BANK_SEL_36, 
        Y => \ELINK_DOUTA_1_m[6]\);
    
    \REG_STATE_0_RNIDUOH1[3]\ : NOR2B
      port map(A => N_1352_2, B => N_1359_1, Y => N_1404_8);
    
    \ELINK_DINA_18[2]\ : DFN1E0C0
      port map(D => \N_TFC_DINA[2]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_21, E => N_198, Q => 
        \ELINK_DINA_18[2]_net_1\);
    
    \REG_STATE_0_RNIVN1B5[2]\ : OR2
      port map(A => un1_REG_STATE_18, B => N_675, Y => SI_CNTe);
    
    \N_TFC_ADDRA_0_o2_RNO_5[7]\ : OA1
      port map(A => \SM_BANK_SEL[20]_net_1\, B => \ELK_N_ACTIVE\, 
        C => \REG_STATE_0[4]_net_1\, Y => 
        \N_TFC_ADDRA_0_a2_6_0[7]\);
    
    \RD_XFER_TYPE[7]\ : DFN1C0
      port map(D => \RD_XFER_TYPE_RNO[7]_net_1\, CLK => CLK60MHZ, 
        CLR => P_USB_MASTER_EN_c, Q => \RD_XFER_TYPE[7]_net_1\);
    
    \ELINK_RWA_RNO_0[13]\ : AOI1
      port map(A => \N_ELINK_RWA_0_iv_0_o2_i_a5_0[13]\, B => 
        N_503, C => \ELINK_RWA[13]_net_1\, Y => N_177);
    
    \ELINK_ADDRA_4[2]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[2]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_2, E => un1_SM_BANK_SEL_8, Q => 
        \ELINK_ADDRA_4[2]_net_1\);
    
    \WR_USB_ADBUS_RNO_2[4]\ : OR3
      port map(A => \N_WR_USB_ADBUS_0_iv_14[4]\, B => 
        \N_WR_USB_ADBUS_0_iv_13[4]\, C => 
        \N_WR_USB_ADBUS_0_iv_22[4]\, Y => 
        \N_WR_USB_ADBUS_0_iv_25[4]\);
    
    \ELINKS_STRT_ADDR_T[3]\ : DFN1E1C0
      port map(D => \RD_USB_ADBUS[3]_net_1\, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_21, E => 
        N_ELINKS_STRT_ADDR_T_0_sqmuxa, Q => 
        \ELINKS_STRT_ADDR_T[3]_net_1\);
    
    \WR_USB_ADBUS_RNO_19[6]\ : AO1
      port map(A => \CHKSUM[6]_net_1\, B => un1_REG_STATE_4, C
         => \N_WR_USB_ADBUS_0_iv_2[6]\, Y => 
        \N_WR_USB_ADBUS_0_iv_4[6]\);
    
    \REG_STATE_ns_i_i_o2_1_RNO[0]\ : OA1
      port map(A => N_438, B => N_439, C => 
        \REG_STATE_0[2]_net_1\, Y => N_444);
    
    \SM_BANK_SEL[6]\ : DFN1E1C0
      port map(D => N_1837, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_7, E => un1_REG_STATE_30, Q => 
        \SM_BANK_SEL[6]_net_1\);
    
    \ELINK_BLKA_RNO[18]\ : AOI1B
      port map(A => \SM_BANK_SEL[1]_net_1\, B => X_BLKA_i, C => 
        N_63_tz, Y => N_63);
    
    \WR_USB_ADBUS_RNO_32[7]\ : NOR2B
      port map(A => \ELINK_DOUTA_0[7]\, B => un1_SM_BANK_SEL_31, 
        Y => \ELINK_DOUTA_0_m[7]\);
    
    \ELINK_RWA_RNO[11]\ : OA1B
      port map(A => N_393, B => \ELINK_RWA[11]_net_1\, C => N_180, 
        Y => \N_ELINK_RWA_0_iv[11]\);
    
    U104_PATT_ELINK_BLK : DPRT_512X9_SRAM_4
      port map(ELINK_RWA_0 => \ELINK_RWA[4]_net_1\, 
        ELK_RX_SER_WORD_4(7) => ELK_RX_SER_WORD_4(7), 
        ELK_RX_SER_WORD_4(6) => ELK_RX_SER_WORD_4(6), 
        ELK_RX_SER_WORD_4(5) => ELK_RX_SER_WORD_4(5), 
        ELK_RX_SER_WORD_4(4) => ELK_RX_SER_WORD_4(4), 
        ELK_RX_SER_WORD_4(3) => ELK_RX_SER_WORD_4(3), 
        ELK_RX_SER_WORD_4(2) => ELK_RX_SER_WORD_4(2), 
        ELK_RX_SER_WORD_4(1) => ELK_RX_SER_WORD_4(1), 
        ELK_RX_SER_WORD_4(0) => ELK_RX_SER_WORD_4(0), 
        ELINK_DINA_4(7) => \ELINK_DINA_4[7]_net_1\, 
        ELINK_DINA_4(6) => \ELINK_DINA_4[6]_net_1\, 
        ELINK_DINA_4(5) => \ELINK_DINA_4[5]_net_1\, 
        ELINK_DINA_4(4) => \ELINK_DINA_4[4]_net_1\, 
        ELINK_DINA_4(3) => \ELINK_DINA_4[3]_net_1\, 
        ELINK_DINA_4(2) => \ELINK_DINA_4[2]_net_1\, 
        ELINK_DINA_4(1) => \ELINK_DINA_4[1]_net_1\, 
        ELINK_DINA_4(0) => \ELINK_DINA_4[0]_net_1\, ELINK_BLKA_0
         => \ELINK_BLKA[4]_net_1\, ELKS_ADDRB(7) => ELKS_ADDRB(7), 
        ELKS_ADDRB(6) => ELKS_ADDRB(6), ELKS_ADDRB(5) => 
        ELKS_ADDRB(5), ELKS_ADDRB(4) => ELKS_ADDRB(4), 
        ELKS_ADDRB(3) => ELKS_ADDRB(3), ELKS_ADDRB(2) => 
        ELKS_ADDRB(2), ELKS_ADDRB(1) => ELKS_ADDRB(1), 
        ELKS_ADDRB(0) => ELKS_ADDRB(0), ELINK_ADDRA_4(7) => 
        \ELINK_ADDRA_4[7]_net_1\, ELINK_ADDRA_4(6) => 
        \ELINK_ADDRA_4[6]_net_1\, ELINK_ADDRA_4(5) => 
        \ELINK_ADDRA_4[5]_net_1\, ELINK_ADDRA_4(4) => 
        \ELINK_ADDRA_4[4]_net_1\, ELINK_ADDRA_4(3) => 
        \ELINK_ADDRA_4[3]_net_1\, ELINK_ADDRA_4(2) => 
        \ELINK_ADDRA_4[2]_net_1\, ELINK_ADDRA_4(1) => 
        \ELINK_ADDRA_4[1]_net_1\, ELINK_ADDRA_4(0) => 
        \ELINK_ADDRA_4[0]_net_1\, PATT_ELK_DAT_4(7) => 
        PATT_ELK_DAT_4(7), PATT_ELK_DAT_4(6) => PATT_ELK_DAT_4(6), 
        PATT_ELK_DAT_4(5) => PATT_ELK_DAT_4(5), PATT_ELK_DAT_4(4)
         => PATT_ELK_DAT_4(4), PATT_ELK_DAT_4(3) => 
        PATT_ELK_DAT_4(3), PATT_ELK_DAT_4(2) => PATT_ELK_DAT_4(2), 
        PATT_ELK_DAT_4(1) => PATT_ELK_DAT_4(1), PATT_ELK_DAT_4(0)
         => PATT_ELK_DAT_4(0), ELINK_DOUTA_4(7) => 
        \ELINK_DOUTA_4[7]\, ELINK_DOUTA_4(6) => 
        \ELINK_DOUTA_4[6]\, ELINK_DOUTA_4(5) => 
        \ELINK_DOUTA_4[5]\, ELINK_DOUTA_4(4) => 
        \ELINK_DOUTA_4[4]\, ELINK_DOUTA_4(3) => 
        \ELINK_DOUTA_4[3]\, ELINK_DOUTA_4(2) => 
        \ELINK_DOUTA_4[2]\, ELINK_DOUTA_4(1) => 
        \ELINK_DOUTA_4[1]\, ELINK_DOUTA_4(0) => 
        \ELINK_DOUTA_4[0]\, ELKS_RWB => ELKS_RWB, 
        P_USB_MASTER_EN_c_0 => P_USB_MASTER_EN_c_0, CLK_40M_GL
         => CLK_40M_GL, CLK60MHZ => CLK60MHZ, ELKS_RAM_BLKB_EN
         => ELKS_RAM_BLKB_EN);
    
    \SM_BANK_SEL_RNIN973[19]\ : OR3
      port map(A => \SM_BANK_SEL[17]_net_1\, B => 
        \SM_BANK_SEL[19]_net_1\, C => N_616_2, Y => 
        \N_ELINK_RWA_1[1]\);
    
    \ELINK_ADDRA_2[7]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[7]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_21, E => un1_SM_BANK_SEL_5, Q => 
        \ELINK_ADDRA_2[7]_net_1\);
    
    \WR_USB_ADBUS_RNO_7[0]\ : AO1
      port map(A => \ELINK_DOUTA_4[0]\, B => un1_SM_BANK_SEL_28, 
        C => \ELINK_DOUTA_5_m[0]\, Y => 
        \N_WR_USB_ADBUS_0_iv_7[0]\);
    
    \ELINK_ADDRA_13[5]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[5]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_3, E => un1_SM_BANK_SEL_2, Q => 
        \ELINK_ADDRA_13[5]_net_1\);
    
    \ELINK_ADDRA_8[5]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[5]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_8, E => un1_SM_BANK_SEL_21, Q => 
        \ELINK_ADDRA_8[5]_net_1\);
    
    \OP_MODE[4]\ : DFN1E1C0
      port map(D => \OP_MODE_T[4]_net_1\, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_15, E => \REG_STATE_d[30]\, Q => 
        \OP_MODE[4]_net_1\);
    
    \N_WR_USB_ADBUS_0_iv_0[6]\ : OR2
      port map(A => \TFC_STOP_ADDR_m[6]\, B => N_1562_i, Y => 
        \N_WR_USB_ADBUS_0_iv_0[6]_net_1\);
    
    \ELINK_ADDRA_8[1]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[1]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_8, E => un1_SM_BANK_SEL_21, Q => 
        \ELINK_ADDRA_8[1]_net_1\);
    
    \WR_XFER_TYPE_RNO_0[4]\ : OA1C
      port map(A => \RD_USB_ADBUS[5]_net_1\, B => N_1717, C => 
        \WR_XFER_TYPE[4]_net_1\, Y => N_1827);
    
    U119_PATT_ELINK_BLK : DPRT_512X9_SRAM_19
      port map(ELINK_RWA_0 => \ELINK_RWA[19]_net_1\, 
        ELK_RX_SER_WORD_19(7) => ELK_RX_SER_WORD_19(7), 
        ELK_RX_SER_WORD_19(6) => ELK_RX_SER_WORD_19(6), 
        ELK_RX_SER_WORD_19(5) => ELK_RX_SER_WORD_19(5), 
        ELK_RX_SER_WORD_19(4) => ELK_RX_SER_WORD_19(4), 
        ELK_RX_SER_WORD_19(3) => ELK_RX_SER_WORD_19(3), 
        ELK_RX_SER_WORD_19(2) => ELK_RX_SER_WORD_19(2), 
        ELK_RX_SER_WORD_19(1) => ELK_RX_SER_WORD_19(1), 
        ELK_RX_SER_WORD_19(0) => ELK_RX_SER_WORD_19(0), 
        ELINK_DINA_19(7) => \ELINK_DINA_19[7]_net_1\, 
        ELINK_DINA_19(6) => \ELINK_DINA_19[6]_net_1\, 
        ELINK_DINA_19(5) => \ELINK_DINA_19[5]_net_1\, 
        ELINK_DINA_19(4) => \ELINK_DINA_19[4]_net_1\, 
        ELINK_DINA_19(3) => \ELINK_DINA_19[3]_net_1\, 
        ELINK_DINA_19(2) => \ELINK_DINA_19[2]_net_1\, 
        ELINK_DINA_19(1) => \ELINK_DINA_19[1]_net_1\, 
        ELINK_DINA_19(0) => \ELINK_DINA_19[0]_net_1\, 
        ELINK_BLKA_0 => \ELINK_BLKA[19]_net_1\, ELKS_ADDRB(7) => 
        ELKS_ADDRB(7), ELKS_ADDRB(6) => ELKS_ADDRB(6), 
        ELKS_ADDRB(5) => ELKS_ADDRB(5), ELKS_ADDRB(4) => 
        ELKS_ADDRB(4), ELKS_ADDRB(3) => ELKS_ADDRB(3), 
        ELKS_ADDRB(2) => ELKS_ADDRB(2), ELKS_ADDRB(1) => 
        ELKS_ADDRB(1), ELKS_ADDRB(0) => ELKS_ADDRB(0), 
        ELINK_ADDRA_19(7) => \ELINK_ADDRA_19[7]_net_1\, 
        ELINK_ADDRA_19(6) => \ELINK_ADDRA_19[6]_net_1\, 
        ELINK_ADDRA_19(5) => \ELINK_ADDRA_19[5]_net_1\, 
        ELINK_ADDRA_19(4) => \ELINK_ADDRA_19[4]_net_1\, 
        ELINK_ADDRA_19(3) => \ELINK_ADDRA_19[3]_net_1\, 
        ELINK_ADDRA_19(2) => \ELINK_ADDRA_19[2]_net_1\, 
        ELINK_ADDRA_19(1) => \ELINK_ADDRA_19[1]_net_1\, 
        ELINK_ADDRA_19(0) => \ELINK_ADDRA_19[0]_net_1\, 
        PATT_ELK_DAT_19(7) => PATT_ELK_DAT_19(7), 
        PATT_ELK_DAT_19(6) => PATT_ELK_DAT_19(6), 
        PATT_ELK_DAT_19(5) => PATT_ELK_DAT_19(5), 
        PATT_ELK_DAT_19(4) => PATT_ELK_DAT_19(4), 
        PATT_ELK_DAT_19(3) => PATT_ELK_DAT_19(3), 
        PATT_ELK_DAT_19(2) => PATT_ELK_DAT_19(2), 
        PATT_ELK_DAT_19(1) => PATT_ELK_DAT_19(1), 
        PATT_ELK_DAT_19(0) => PATT_ELK_DAT_19(0), 
        ELINK_DOUTA_19(7) => \ELINK_DOUTA_19[7]\, 
        ELINK_DOUTA_19(6) => \ELINK_DOUTA_19[6]\, 
        ELINK_DOUTA_19(5) => \ELINK_DOUTA_19[5]\, 
        ELINK_DOUTA_19(4) => \ELINK_DOUTA_19[4]\, 
        ELINK_DOUTA_19(3) => \ELINK_DOUTA_19[3]\, 
        ELINK_DOUTA_19(2) => \ELINK_DOUTA_19[2]\, 
        ELINK_DOUTA_19(1) => \ELINK_DOUTA_19[1]\, 
        ELINK_DOUTA_19(0) => \ELINK_DOUTA_19[0]\, ELKS_RWB => 
        ELKS_RWB, P_USB_MASTER_EN_c_0 => P_USB_MASTER_EN_c_0, 
        CLK_40M_GL => CLK_40M_GL, CLK60MHZ => CLK60MHZ, 
        ELKS_RAM_BLKB_EN => ELKS_RAM_BLKB_EN);
    
    \ELINK_BLKA[8]\ : DFN1E0P0
      port map(D => \N_ELINK_BLKA_0_iv[8]\, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_19, E => \SM_BANK_SEL[20]_net_1\, Q
         => \ELINK_BLKA[8]_net_1\);
    
    \SM_BANK_SEL_RNI3OV62[18]\ : NOR3A
      port map(A => \SM_BANK_SEL[18]_net_1\, B => N_312_0, C => 
        N_1566_i_i_0, Y => un1_SM_BANK_SEL_36);
    
    \REG_STATE_0_RNIGPV6T1[0]\ : NOR2
      port map(A => \REG_STATE_ns_i_1_0[3]\, B => 
        \REG_STATE_ns_i_0[3]\, Y => 
        \REG_STATE_0_RNIGPV6T1[0]_net_1\);
    
    \ELINK_BLKA_RNO[2]\ : OA1C
      port map(A => N_618, B => \ELINK_BLKA[2]_net_1\, C => 
        X_BLKA_i_m_1, Y => \N_ELINK_BLKA_0_iv[2]\);
    
    \WR_USB_ADBUS_RNO_0[4]\ : OR3
      port map(A => \N_WR_USB_ADBUS_0_iv_10[4]\, B => 
        \N_WR_USB_ADBUS_0_iv_9[4]\, C => 
        \N_WR_USB_ADBUS_0_iv_20[4]\, Y => 
        \N_WR_USB_ADBUS_0_iv_24[4]\);
    
    \WR_USB_ADBUS_RNO_35[3]\ : NOR2B
      port map(A => \ELINK_DOUTA_0[3]\, B => un1_SM_BANK_SEL_31, 
        Y => \ELINK_DOUTA_0_m[3]\);
    
    \REG_ADDR_RNIM1HE[2]\ : NOR2
      port map(A => \REG_ADDR[4]_net_1\, B => \REG_ADDR[2]_net_1\, 
        Y => REG_STATE_tr73_2);
    
    \ELINK_DINA_9[3]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[3]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_20, E => un1_SM_BANK_SEL_9, Q => 
        \ELINK_DINA_9[3]_net_1\);
    
    \ELINK_ADDRA_16[1]\ : DFN1E0C0
      port map(D => \N_TFC_ADDRA[1]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_8, E => N_200, Q => 
        \ELINK_ADDRA_16[1]_net_1\);
    
    \SM_BANK_SEL_RNIT4VN[14]\ : OR3A
      port map(A => N_143, B => N_616_11, C => N_620_10, Y => 
        \N_ELINK_RWA_1[4]\);
    
    USB_TXE_B_RNI1P4IJ : NOR3B
      port map(A => \REG_STATE_ns_i_a2_0_0[5]\, B => N_2576, C
         => N_1419, Y => N_2581);
    
    \REG_ADDR_RNO[6]\ : XA1B
      port map(A => REG_ADDR_c5, B => \REG_ADDR[6]_net_1\, C => 
        N_675_0, Y => REG_ADDR_n6);
    
    \REG_ADDR_RNO[3]\ : XA1B
      port map(A => N_474, B => \REG_ADDR[3]_net_1\, C => N_675_0, 
        Y => REG_ADDR_n3);
    
    \OP_MODE[3]\ : DFN1E1C0
      port map(D => \OP_MODE_T[3]_net_1\, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_15, E => \REG_STATE_d[30]\, Q => 
        \OP_MODE[3]_net_1\);
    
    \WR_USB_ADBUS_RNO_6[3]\ : OR3
      port map(A => \N_WR_USB_ADBUS_0_iv_3[3]\, B => 
        \N_WR_USB_ADBUS_0_iv_2[3]\, C => 
        \N_WR_USB_ADBUS_0_iv_4[3]\, Y => 
        \N_WR_USB_ADBUS_0_iv_6[3]\);
    
    \WR_USB_ADBUS_RNO_4[5]\ : AO1
      port map(A => \ELINK_DOUTA_16[5]\, B => un1_SM_BANK_SEL_39, 
        C => \ELINK_DOUTA_1_m[5]\, Y => 
        \N_WR_USB_ADBUS_0_iv_9[5]\);
    
    \WR_USB_ADBUS_RNO_11[5]\ : OR3
      port map(A => \ELINK_DOUTA_11_m[5]\, B => 
        \ELINK_DOUTA_10_m[5]\, C => \N_WR_USB_ADBUS_0_iv_16[5]\, 
        Y => \N_WR_USB_ADBUS_0_iv_22[5]\);
    
    \TFC_DINA[1]\ : DFN1E0C0
      port map(D => \N_TFC_DINA[1]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_4, E => N_142, Q => \TFC_DINA[1]_net_1\);
    
    \SM_BANK_SEL_RNI7A6G[9]\ : OR2
      port map(A => \SM_BANK_SEL[9]_net_1\, B => 
        \SM_BANK_SEL_0[21]_net_1\, Y => un1_SM_BANK_SEL_20);
    
    \REG_STATE_RNIP1GM1[2]\ : OR2A
      port map(A => \REG_STATE[2]_net_1\, B => N_256, Y => N_264);
    
    \ELINK_DINA_0[4]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[4]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_5, E => un1_SM_BANK_SEL_6, Q => 
        \ELINK_DINA_0[4]_net_1\);
    
    \REG_STATE_RNIVU1F2[1]\ : NOR2B
      port map(A => N_1745_i, B => N_1907, Y => 
        N_ELINKS_STOP_ADDR_T_0_sqmuxa);
    
    \ELINK_ADDRA_14[0]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[0]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_5, E => un1_SM_BANK_SEL_1, Q => 
        \ELINK_ADDRA_14[0]_net_1\);
    
    \WR_XFER_TYPE_RNI3JSS[3]\ : NOR2
      port map(A => \WR_XFER_TYPE[3]_net_1\, B => 
        \WR_XFER_TYPE[4]_net_1\, Y => N_1404_6);
    
    \SM_BANK_SEL_RNICON91[9]\ : NOR3C
      port map(A => N_461, B => 
        \N_ELINK_BLKA_0_iv_0_o2_i_a5_0[9]\, C => N_477, Y => 
        \N_ELINK_BLKA_0_iv_0_o2_i_a5_2[9]\);
    
    \REG_STATE_RNI3PF72[0]\ : OR2
      port map(A => REG_STATE_s22_i_0, B => N_2497, Y => N_1499);
    
    \REG_STATE_0_RNIAVT12[1]\ : OAI1
      port map(A => \REG_STATE_0[1]_net_1\, B => N_268, C => 
        N_2462, Y => N_2520);
    
    \RD_USB_ADBUS_RNIBNBG1[4]\ : NOR2B
      port map(A => N_1903, B => N_290, Y => N_1893);
    
    \WR_USB_ADBUS_RNO_33[5]\ : NOR2B
      port map(A => \WR_XFER_TYPE[5]_net_1\, B => N_398, Y => 
        \WR_XFER_TYPE_m[5]\);
    
    \ELINK_DINA_5[3]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[3]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_14, E => un1_SM_BANK_SEL_15, Q => 
        \ELINK_DINA_5[3]_net_1\);
    
    \ELINK_DINA_4[7]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[7]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_13, E => un1_SM_BANK_SEL_8, Q => 
        \ELINK_DINA_4[7]_net_1\);
    
    \WR_USB_ADBUS_RNO_15[7]\ : NOR2B
      port map(A => \ELINK_DOUTA_18[7]\, B => un1_SM_BANK_SEL_25, 
        Y => \ELINK_DOUTA_18_m[7]\);
    
    un1_REG_STATE_4_0_a2_RNO : NOR3B
      port map(A => \REG_STATE_0[5]_net_1\, B => 
        \REG_STATE[2]_net_1\, C => \REG_STATE_0[0]_net_1\, Y => 
        un1_REG_STATE_4_0_a2_1);
    
    \SM_BANK_SEL_RNO[17]\ : NOR3B
      port map(A => N_1882, B => N_1352_4, C => N_1700, Y => 
        N_1851);
    
    \CHKSUM[1]\ : DFN1E1C0
      port map(D => N_236, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_3, E => un1_REG_STATE_22, Q => 
        \CHKSUM[1]_net_1\);
    
    \ELINK_ADDRA_18[1]\ : DFN1E0C0
      port map(D => \N_TFC_ADDRA[1]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_12, E => N_198, Q => 
        \ELINK_ADDRA_18[1]_net_1\);
    
    USB_RXF_B_RNIDHGV31 : NOR2B
      port map(A => \REG_STATE_ns_i_a2_1[4]\, B => N_2581, Y => 
        N_2597);
    
    \WR_USB_ADBUS_RNO_14[5]\ : NOR2B
      port map(A => \ELINK_DOUTA_3[5]\, B => un1_SM_BANK_SEL_43, 
        Y => \ELINK_DOUTA_3_m[5]\);
    
    \ELINK_ADDRA_12[0]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[0]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_2_0, E => un1_SM_BANK_SEL_7, Q => 
        \ELINK_ADDRA_12[0]_net_1\);
    
    \WR_USB_ADBUS_RNO_5[3]\ : OR3
      port map(A => \ELINK_DOUTA_3_m[3]\, B => 
        \ELINK_DOUTA_18_m[3]\, C => \N_WR_USB_ADBUS_0_iv_12[3]\, 
        Y => \N_WR_USB_ADBUS_0_iv_20[3]\);
    
    USB_RD_BI_RNO_12 : NOR2A
      port map(A => N_1352_4, B => N_293, Y => 
        N_USB_RD_BI_i_a2_4_3);
    
    \WR_USB_ADBUS_RNO_8[4]\ : OR3
      port map(A => \N_WR_USB_ADBUS_0_iv_5[4]\, B => 
        \N_WR_USB_ADBUS_0_iv_4[4]\, C => \ELINK_DOUTA_3_m[4]\, Y
         => \N_WR_USB_ADBUS_0_iv_17[4]\);
    
    \WR_USB_ADBUS_RNO_33[3]\ : NOR2A
      port map(A => \ELINKS_STRT_ADDR[3]_net_1\, B => N_1499, Y
         => \ELINKS_STRT_ADDR_m[3]\);
    
    \ELINK_DINA_18[0]\ : DFN1E0C0
      port map(D => \N_TFC_DINA[0]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_20, E => N_198, Q => 
        \ELINK_DINA_18[0]_net_1\);
    
    \SI_CNT[1]\ : DFN1E1C0
      port map(D => SI_CNT_n1, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_5, E => SI_CNTe, Q => \SI_CNT[1]_net_1\);
    
    \ELINK_BLKA[3]\ : DFN1E0P0
      port map(D => \N_ELINK_BLKA_0_iv[3]\, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_19, E => \SM_BANK_SEL[20]_net_1\, Q
         => \ELINK_BLKA[3]_net_1\);
    
    \USB_OE_BI\ : DFN1E0P0
      port map(D => N_1679, CLK => CLK60MHZ, PRE => 
        P_USB_MASTER_EN_c_19, E => N_1669, Q => USB_OE_BI);
    
    \WR_XFER_TYPE_RNIDDIL5[5]\ : NOR2B
      port map(A => REG_STATE_tr72_6_5, B => N_1404_8, Y => 
        N_1419);
    
    \WR_USB_ADBUS_RNO_20[1]\ : NOR2A
      port map(A => \TFC_DOUTA[1]\, B => N_243, Y => 
        \TFC_DOUTA_m[1]\);
    
    \ELINKS_STRT_ADDR_T[4]\ : DFN1E1C0
      port map(D => \RD_USB_ADBUS[4]_net_1\, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_21, E => 
        N_ELINKS_STRT_ADDR_T_0_sqmuxa, Q => 
        \ELINKS_STRT_ADDR_T[4]_net_1\);
    
    \SM_BANK_SEL_RNI0LV62[15]\ : NOR3A
      port map(A => \SM_BANK_SEL[15]_net_1\, B => N_312_0, C => 
        N_1566_i_i_0, Y => un1_SM_BANK_SEL_28);
    
    \WR_USB_ADBUS_RNO_8[5]\ : OR3
      port map(A => \TFC_DOUTA_m[5]\, B => \ELINK_DOUTA_19_m[5]\, 
        C => \N_WR_USB_ADBUS_0_iv_8[5]\, Y => 
        \N_WR_USB_ADBUS_0_iv_18[5]\);
    
    \SM_BANK_SEL_RNI27E6[12]\ : OR3
      port map(A => N_622_3, B => N_616_4, C => N_620_10, Y => 
        \N_ELINK_RWA_1[6]\);
    
    \ELINK_ADDRA_8[7]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[7]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_8, E => un1_SM_BANK_SEL_21, Q => 
        \ELINK_ADDRA_8[7]_net_1\);
    
    \ELINK_DINA_5[4]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[4]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_14, E => un1_SM_BANK_SEL_15, Q => 
        \ELINK_DINA_5[4]_net_1\);
    
    \ELINK_ADDRA_14[7]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[7]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_5, E => un1_SM_BANK_SEL_1, Q => 
        \ELINK_ADDRA_14[7]_net_1\);
    
    \WR_USB_ADBUS_RNO_8[3]\ : OR3
      port map(A => \TFC_DOUTA_m[3]\, B => \ELINK_DOUTA_19_m[3]\, 
        C => \N_WR_USB_ADBUS_0_iv_8[3]\, Y => 
        \N_WR_USB_ADBUS_0_iv_18[3]\);
    
    \ELINK_DINA_14[3]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[3]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_16, E => un1_SM_BANK_SEL_1, Q => 
        \ELINK_DINA_14[3]_net_1\);
    
    \ELINK_ADDRA_14[4]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[4]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_5, E => un1_SM_BANK_SEL_1, Q => 
        \ELINK_ADDRA_14[4]_net_1\);
    
    \SM_BANK_SEL_RNIFOJ1[18]\ : OR2
      port map(A => \SM_BANK_SEL[18]_net_1\, B => 
        \SM_BANK_SEL[19]_net_1\, Y => N_618_1);
    
    U107_PATT_ELINK_BLK : DPRT_512X9_SRAM_7
      port map(ELINK_RWA_0 => \ELINK_RWA[7]_net_1\, 
        ELK_RX_SER_WORD_7(7) => ELK_RX_SER_WORD_7(7), 
        ELK_RX_SER_WORD_7(6) => ELK_RX_SER_WORD_7(6), 
        ELK_RX_SER_WORD_7(5) => ELK_RX_SER_WORD_7(5), 
        ELK_RX_SER_WORD_7(4) => ELK_RX_SER_WORD_7(4), 
        ELK_RX_SER_WORD_7(3) => ELK_RX_SER_WORD_7(3), 
        ELK_RX_SER_WORD_7(2) => ELK_RX_SER_WORD_7(2), 
        ELK_RX_SER_WORD_7(1) => ELK_RX_SER_WORD_7(1), 
        ELK_RX_SER_WORD_7(0) => ELK_RX_SER_WORD_7(0), 
        ELINK_DINA_7(7) => \ELINK_DINA_7[7]_net_1\, 
        ELINK_DINA_7(6) => \ELINK_DINA_7[6]_net_1\, 
        ELINK_DINA_7(5) => \ELINK_DINA_7[5]_net_1\, 
        ELINK_DINA_7(4) => \ELINK_DINA_7[4]_net_1\, 
        ELINK_DINA_7(3) => \ELINK_DINA_7[3]_net_1\, 
        ELINK_DINA_7(2) => \ELINK_DINA_7[2]_net_1\, 
        ELINK_DINA_7(1) => \ELINK_DINA_7[1]_net_1\, 
        ELINK_DINA_7(0) => \ELINK_DINA_7[0]_net_1\, ELINK_BLKA_0
         => \ELINK_BLKA[7]_net_1\, ELKS_ADDRB_0_d0 => 
        ELKS_ADDRB(0), ELKS_ADDRB_1 => ELKS_ADDRB(1), 
        ELKS_ADDRB_3 => ELKS_ADDRB(3), ELKS_ADDRB_5 => 
        ELKS_ADDRB(5), ELKS_ADDRB_7 => ELKS_ADDRB(7), 
        ELKS_ADDRB_0_0 => ELKS_ADDRB_0_0, ELKS_ADDRB_0_2 => 
        ELKS_ADDRB_0_2, ELKS_ADDRB_0_4 => ELKS_ADDRB_0_4, 
        ELINK_ADDRA_7(7) => \ELINK_ADDRA_7[7]_net_1\, 
        ELINK_ADDRA_7(6) => \ELINK_ADDRA_7[6]_net_1\, 
        ELINK_ADDRA_7(5) => \ELINK_ADDRA_7[5]_net_1\, 
        ELINK_ADDRA_7(4) => \ELINK_ADDRA_7[4]_net_1\, 
        ELINK_ADDRA_7(3) => \ELINK_ADDRA_7[3]_net_1\, 
        ELINK_ADDRA_7(2) => \ELINK_ADDRA_7[2]_net_1\, 
        ELINK_ADDRA_7(1) => \ELINK_ADDRA_7[1]_net_1\, 
        ELINK_ADDRA_7(0) => \ELINK_ADDRA_7[0]_net_1\, 
        PATT_ELK_DAT_7(7) => PATT_ELK_DAT_7(7), PATT_ELK_DAT_7(6)
         => PATT_ELK_DAT_7(6), PATT_ELK_DAT_7(5) => 
        PATT_ELK_DAT_7(5), PATT_ELK_DAT_7(4) => PATT_ELK_DAT_7(4), 
        PATT_ELK_DAT_7(3) => PATT_ELK_DAT_7(3), PATT_ELK_DAT_7(2)
         => PATT_ELK_DAT_7(2), PATT_ELK_DAT_7(1) => 
        PATT_ELK_DAT_7(1), PATT_ELK_DAT_7(0) => PATT_ELK_DAT_7(0), 
        ELINK_DOUTA_7(7) => \ELINK_DOUTA_7[7]\, ELINK_DOUTA_7(6)
         => \ELINK_DOUTA_7[6]\, ELINK_DOUTA_7(5) => 
        \ELINK_DOUTA_7[5]\, ELINK_DOUTA_7(4) => 
        \ELINK_DOUTA_7[4]\, ELINK_DOUTA_7(3) => 
        \ELINK_DOUTA_7[3]\, ELINK_DOUTA_7(2) => 
        \ELINK_DOUTA_7[2]\, ELINK_DOUTA_7(1) => 
        \ELINK_DOUTA_7[1]\, ELINK_DOUTA_7(0) => 
        \ELINK_DOUTA_7[0]\, ELKS_RWB => ELKS_RWB, 
        P_USB_MASTER_EN_c_0 => P_USB_MASTER_EN_c_0, CLK_40M_GL
         => CLK_40M_GL, CLK60MHZ => CLK60MHZ, ELKS_RAM_BLKB_EN
         => ELKS_RAM_BLKB_EN);
    
    \RD_USB_ADBUS_RNIK0CG1[5]\ : AO1C
      port map(A => N_1700, B => \RD_USB_ADBUS[5]_net_1\, C => 
        N_293, Y => N_1698);
    
    \WR_USB_ADBUS_RNO_3[7]\ : AO1
      port map(A => \ELINK_DOUTA_17[7]\, B => un1_SM_BANK_SEL_40, 
        C => \ELINK_DOUTA_2_m[7]\, Y => 
        \N_WR_USB_ADBUS_0_iv_10[7]\);
    
    \ELINK_DINA_18[5]\ : DFN1E0C0
      port map(D => \N_TFC_DINA[5]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_21, E => N_198, Q => 
        \ELINK_DINA_18[5]_net_1\);
    
    \ELINK_BLKA_RNO[0]\ : AOI1
      port map(A => \SM_BANK_SEL[19]_net_1\, B => X_BLKA_i, C => 
        \ELINK_BLKA_i_m[0]\, Y => \N_ELINK_BLKA_0_iv[0]\);
    
    \ELINK_ADDRA_8[3]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[3]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_8, E => un1_SM_BANK_SEL_21, Q => 
        \ELINK_ADDRA_8[3]_net_1\);
    
    \WR_USB_ADBUS_RNO_0[1]\ : OR3
      port map(A => \N_WR_USB_ADBUS_0_iv_10[1]\, B => 
        \N_WR_USB_ADBUS_0_iv_9[1]\, C => 
        \N_WR_USB_ADBUS_0_iv_20[1]\, Y => 
        \N_WR_USB_ADBUS_0_iv_24[1]\);
    
    \ELINKS_STOP_ADDR[2]\ : DFN1E1C0
      port map(D => \ELINKS_STOP_ADDR_T[2]_net_1\, CLK => 
        CLK60MHZ, CLR => P_USB_MASTER_EN_c_14, E => 
        \REG_STATE_d_0[30]\, Q => \ELINKS_STOP_ADDR[2]_net_1\);
    
    \WR_USB_ADBUS_RNO_6[6]\ : AO1
      port map(A => \ELINK_DOUTA_5[6]\, B => un1_SM_BANK_SEL_35, 
        C => \ELINK_DOUTA_6_m[6]\, Y => 
        \N_WR_USB_ADBUS_0_iv_7[6]\);
    
    \SM_BANK_SEL_RNO[11]\ : NOR3B
      port map(A => N_1892, B => N_1902, C => 
        \RD_USB_ADBUS[2]_net_1\, Y => N_1846);
    
    \ELINK_ADDRA_15[0]\ : DFN1E0C0
      port map(D => \N_TFC_ADDRA[0]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_6, E => N_199, Q => 
        \ELINK_ADDRA_15[0]_net_1\);
    
    \SM_BANK_SEL[15]\ : DFN1E1C0
      port map(D => N_1843, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_1_0, E => un1_REG_STATE_30, Q => 
        \SM_BANK_SEL[15]_net_1\);
    
    \ELINK_DINA_18[4]\ : DFN1E0C0
      port map(D => \N_TFC_DINA[4]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_21, E => N_198, Q => 
        \ELINK_DINA_18[4]_net_1\);
    
    \SM_BANK_SEL_RNIC2P72[0]\ : NOR3A
      port map(A => \SM_BANK_SEL[0]_net_1\, B => N_312, C => 
        N_1566_i_i_0, Y => un1_SM_BANK_SEL_41);
    
    \ELINK_DINA_4[4]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[4]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_13, E => un1_SM_BANK_SEL_8, Q => 
        \ELINK_DINA_4[4]_net_1\);
    
    \WR_USB_ADBUS_RNO_16[3]\ : AO1
      port map(A => \ELINK_DOUTA_4[3]\, B => un1_SM_BANK_SEL_28, 
        C => \ELINK_DOUTA_5_m[3]\, Y => 
        \N_WR_USB_ADBUS_0_iv_12[3]\);
    
    \ELINK_DINA_7[0]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[0]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_17, E => un1_SM_BANK_SEL_12, Q => 
        \ELINK_DINA_7[0]_net_1\);
    
    \ELINK_DINA_17[1]\ : DFN1E0C0
      port map(D => \N_TFC_DINA[1]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_19, E => N_197, Q => 
        \ELINK_DINA_17[1]_net_1\);
    
    \REG_STATE_0_RNIBRL53[2]\ : MX2
      port map(A => N_346, B => N_2616, S => 
        \REG_STATE_0[2]_net_1\, Y => N_349);
    
    \WR_XFER_TYPE[1]\ : DFN1C0
      port map(D => \WR_XFER_TYPE_RNO[1]_net_1\, CLK => CLK60MHZ, 
        CLR => P_USB_MASTER_EN_c, Q => \WR_XFER_TYPE[1]_net_1\);
    
    \WR_USB_ADBUS_RNO_24[4]\ : NOR2B
      port map(A => \ELINK_DOUTA_17[4]\, B => un1_SM_BANK_SEL_40, 
        Y => \ELINK_DOUTA_17_m[4]\);
    
    \REG_STATE_0_RNIO8J481[1]\ : OA1
      port map(A => \REG_STATE_ns_i_a4_0[4]\, B => 
        \REG_STATE_ns_i_a4_9_1[4]\, C => N_2597, Y => 
        \REG_STATE_ns_i_4[4]\);
    
    \WR_USB_ADBUS_RNO_32[5]\ : NOR2A
      port map(A => \TFC_STOP_ADDR[5]_net_1\, B => N_1501, Y => 
        \TFC_STOP_ADDR_m[5]\);
    
    \WR_USB_ADBUS_RNO_23[7]\ : NOR2B
      port map(A => \ELINK_DOUTA_9[7]\, B => un1_SM_BANK_SEL_42, 
        Y => \ELINK_DOUTA_9_m[7]\);
    
    \WR_USB_ADBUS_RNO_11[6]\ : OR3
      port map(A => \ELINK_DOUTA_14_m[6]\, B => 
        \ELINK_DOUTA_1_m[6]\, C => \N_WR_USB_ADBUS_0_iv_15[6]\, Y
         => \N_WR_USB_ADBUS_0_iv_21[6]\);
    
    \N_WR_USB_ADBUS_0_iv_0_RNO[2]\ : NOR2A
      port map(A => \TFC_STOP_ADDR[2]_net_1\, B => N_1501, Y => 
        \TFC_STOP_ADDR_m[2]\);
    
    \WR_USB_ADBUS_RNO_36[1]\ : NOR2B
      port map(A => \ELINK_DOUTA_13[1]\, B => un1_SM_BANK_SEL_29, 
        Y => \ELINK_DOUTA_13_m[1]\);
    
    \WR_USB_ADBUS_RNO_0[7]\ : OR3
      port map(A => \N_WR_USB_ADBUS_0_iv_10[7]\, B => 
        \N_WR_USB_ADBUS_0_iv_9[7]\, C => 
        \N_WR_USB_ADBUS_0_iv_20[7]\, Y => 
        \N_WR_USB_ADBUS_0_iv_24[7]\);
    
    \REG_STATE_ns_i_i_o2_1_RNO_7[0]\ : NOR3
      port map(A => \REG_STATE_0[2]_net_1\, B => \USB_TXE_B\, C
         => N_312, Y => N_436);
    
    \ELINKS_STOP_ADDR_T[5]\ : DFN1E1C0
      port map(D => \RD_USB_ADBUS[5]_net_1\, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_7, E => 
        N_ELINKS_STOP_ADDR_T_0_sqmuxa, Q => 
        \ELINKS_STOP_ADDR_T[5]_net_1\);
    
    \RD_XFER_TYPE[6]\ : DFN1C0
      port map(D => \RD_XFER_TYPE_RNO[6]_net_1\, CLK => CLK60MHZ, 
        CLR => P_USB_MASTER_EN_c, Q => \RD_XFER_TYPE[6]_net_1\);
    
    \WR_USB_ADBUS_RNO_30[2]\ : AO1
      port map(A => \ELINK_DOUTA_14[2]\, B => un1_SM_BANK_SEL_23, 
        C => \ELINK_DOUTA_19_m[2]\, Y => 
        \N_WR_USB_ADBUS_0_iv_12[2]\);
    
    \WR_USB_ADBUS_RNO_26[2]\ : NOR2B
      port map(A => \ELINK_DOUTA_11[2]\, B => un1_SM_BANK_SEL_26, 
        Y => \ELINK_DOUTA_11_m[2]\);
    
    \TFC_STRT_ADDR_T[5]\ : DFN1E1C0
      port map(D => \RD_USB_ADBUS[5]_net_1\, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_4, E => N_TFC_STRT_ADDR_T_0_sqmuxa, 
        Q => \TFC_STRT_ADDR_T[5]_net_1\);
    
    \REG_ADDR[8]\ : DFN1E1C0
      port map(D => REG_ADDR_n8, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_10, E => REG_ADDRe, Q => 
        \REG_ADDR[8]_net_1\);
    
    USB_TXE_B_RNIOELU : NOR2A
      port map(A => N_1421_3, B => \USB_TXE_B\, Y => 
        REG_STATE_tr74_0);
    
    un1_REG_STATE_4_0 : OR2
      port map(A => N_1782, B => N_1781, Y => un1_REG_STATE_4);
    
    \WR_USB_ADBUS_RNO_20[4]\ : AO1A
      port map(A => N_1497, B => \TFC_STRT_ADDR[4]_net_1\, C => 
        \N_WR_USB_ADBUS_0_iv_2[4]\, Y => 
        \N_WR_USB_ADBUS_0_iv_4[4]\);
    
    \ELINK_ADDRA_6[0]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[0]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_4, E => un1_SM_BANK_SEL_10, Q => 
        \ELINK_ADDRA_6[0]_net_1\);
    
    \WR_USB_ADBUS_RNO_25[4]\ : NOR2B
      port map(A => \ELINK_DOUTA_1[4]\, B => un1_SM_BANK_SEL_36, 
        Y => \ELINK_DOUTA_1_m[4]\);
    
    \WR_USB_ADBUS_RNO_20[0]\ : AO1A
      port map(A => N_1497, B => \TFC_STRT_ADDR[0]_net_1\, C => 
        \N_WR_USB_ADBUS_0_iv_2[0]\, Y => 
        \N_WR_USB_ADBUS_0_iv_4[0]\);
    
    U4A_REGCROSS : CLK60M_TO_40M_4
      port map(TFC_STRT_ADDR_0(7) => \TFC_STRT_ADDR[7]_net_1\, 
        TFC_STRT_ADDR_0(6) => \TFC_STRT_ADDR[6]_net_1\, 
        TFC_STRT_ADDR_0(5) => \TFC_STRT_ADDR[5]_net_1\, 
        TFC_STRT_ADDR_0(4) => \TFC_STRT_ADDR[4]_net_1\, 
        TFC_STRT_ADDR_0(3) => \TFC_STRT_ADDR[3]_net_1\, 
        TFC_STRT_ADDR_0(2) => \TFC_STRT_ADDR[2]_net_1\, 
        TFC_STRT_ADDR_0(1) => \TFC_STRT_ADDR[1]_net_1\, 
        TFC_STRT_ADDR_0(0) => \TFC_STRT_ADDR[0]_net_1\, 
        TFC_STRT_ADDR(7) => TFC_STRT_ADDR_0(7), TFC_STRT_ADDR(6)
         => TFC_STRT_ADDR_0(6), TFC_STRT_ADDR(5) => 
        TFC_STRT_ADDR_0(5), TFC_STRT_ADDR(4) => 
        TFC_STRT_ADDR_0(4), TFC_STRT_ADDR(3) => 
        TFC_STRT_ADDR_0(3), TFC_STRT_ADDR(2) => 
        TFC_STRT_ADDR_0(2), TFC_STRT_ADDR(1) => 
        TFC_STRT_ADDR_0(1), TFC_STRT_ADDR(0) => 
        TFC_STRT_ADDR_0(0), P_MASTER_POR_B_c_22 => 
        P_MASTER_POR_B_c_22, P_MASTER_POR_B_c_21 => 
        P_MASTER_POR_B_c_21, P_MASTER_POR_B_c_32_0 => 
        P_MASTER_POR_B_c_32_0, P_MASTER_POR_B_c_32 => 
        P_MASTER_POR_B_c_32, P_MASTER_POR_B_c_17 => 
        P_MASTER_POR_B_c_17, P_MASTER_POR_B_c_27 => 
        P_MASTER_POR_B_c_27, CLK_40M_GL => CLK_40M_GL);
    
    un1_N_WR_USB_ADBUS_0_sqmuxa_i_RNO : OR2
      port map(A => N_312, B => N_1566_i_i_0, Y => N_78);
    
    \REG_ADDR_RNO[7]\ : XA1B
      port map(A => REG_ADDR_c6, B => \REG_ADDR[7]_net_1\, C => 
        N_675_0, Y => REG_ADDR_n7);
    
    \WR_USB_ADBUS_RNO_26[7]\ : NOR2B
      port map(A => \ELINK_DOUTA_10[7]\, B => un1_SM_BANK_SEL_34, 
        Y => \ELINK_DOUTA_10_m[7]\);
    
    \REG_STATE_0[5]\ : DFN1C0
      port map(D => \USB_TXE_B_RNIV2O4Q\, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_22_0, Q => \REG_STATE_0[5]_net_1\);
    
    \N_TFC_ADDRA_0_o2_RNO_1[7]\ : NOR3B
      port map(A => N_257, B => \N_TFC_ADDRA_0_a2_1_1[7]\, C => 
        \USB_TXE_B\, Y => N_428);
    
    \WR_USB_ADBUS_RNO_8[7]\ : OR3
      port map(A => \TFC_DOUTA_m[7]\, B => \ELINK_DOUTA_19_m[7]\, 
        C => \N_WR_USB_ADBUS_0_iv_8[7]\, Y => 
        \N_WR_USB_ADBUS_0_iv_18[7]\);
    
    \ELINK_DINA_19[1]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[1]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_0, E => un1_SM_BANK_SEL_11, Q => 
        \ELINK_DINA_19[1]_net_1\);
    
    \SM_BANK_SEL_RNIJ41C2[9]\ : NOR3A
      port map(A => \SM_BANK_SEL[9]_net_1\, B => N_312_0, C => 
        N_1566_i_i_0, Y => un1_SM_BANK_SEL_34);
    
    \RD_USB_ADBUS_RNI4J1Q1[7]\ : OR3
      port map(A => N_459, B => \RD_USB_ADBUS[7]_net_1\, C => 
        N_356, Y => N_1387_i_0_1);
    
    \ELINK_DINA_6[1]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[1]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_16, E => un1_SM_BANK_SEL_10, Q => 
        \ELINK_DINA_6[1]_net_1\);
    
    \CHKSUM_RNO[4]\ : NOR2A
      port map(A => \RD_USB_ADBUS[4]_net_1\, B => N_675, Y => 
        N_232);
    
    USB_RXF_B_RNIJV1A2 : NOR2A
      port map(A => un1_REG_STATE_40_i_a2_2_0, B => N_1713, Y => 
        N_1886);
    
    USB_WR_BI_RNO_2 : XOR2
      port map(A => \REG_STATE[1]_net_1\, B => 
        \REG_STATE[2]_net_1\, Y => N_1761_i);
    
    \SM_BANK_SEL_RNO[9]\ : NOR3B
      port map(A => N_1892, B => N_1352_4, C => 
        \RD_USB_ADBUS[2]_net_1\, Y => N_1847);
    
    \SM_BANK_SEL_RNI9R63[13]\ : OR3
      port map(A => \SM_BANK_SEL[13]_net_1\, B => 
        \SM_BANK_SEL[11]_net_1\, C => N_622_3, Y => 
        \N_ELINK_RWA_1[7]\);
    
    \ELINK_DINA_17[3]\ : DFN1E0C0
      port map(D => \N_TFC_DINA[3]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_19, E => N_197, Q => 
        \ELINK_DINA_17[3]_net_1\);
    
    \OP_MODE_T[6]\ : DFN1E1C0
      port map(D => \RD_USB_ADBUS[6]_net_1\, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_17, E => N_OP_MODE_T_0_sqmuxa, Q
         => \OP_MODE_T[6]_net_1\);
    
    \SI_CNT_RNO[2]\ : XA1B
      port map(A => \SI_CNT[2]_net_1\, B => N_2607, C => N_678, Y
         => N_44);
    
    \RD_USB_ADBUS_RNICJ0T[4]\ : NOR2A
      port map(A => N_290, B => \RD_USB_ADBUS[4]_net_1\, Y => 
        N_1881);
    
    \SM_BANK_SEL_RNI9JK1[19]\ : OR2
      port map(A => \SM_BANK_SEL[19]_net_1\, B => 
        \SM_BANK_SEL[21]_net_1\, Y => un1_SM_BANK_SEL_6);
    
    \REG_STATE_0_RNI7DRP1[5]\ : OA1A
      port map(A => \REG_STATE_0[4]_net_1\, B => N_2617, C => 
        \REG_STATE_0[5]_net_1\, Y => \REG_STATE_ns_i_a4_0[1]\);
    
    \WR_USB_ADBUS_RNO_35[5]\ : NOR2B
      port map(A => \CHKSUM[5]_net_1\, B => un1_REG_STATE_4, Y
         => \CHKSUM_m[5]\);
    
    \REG_STATE_RNI1JQN_0[3]\ : NOR2B
      port map(A => \REG_STATE[3]_net_1\, B => 
        \REG_STATE[2]_net_1\, Y => N_1359_2);
    
    \ELINK_ADDRA_18[0]\ : DFN1E0C0
      port map(D => \N_TFC_ADDRA[0]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_12, E => N_198, Q => 
        \ELINK_ADDRA_18[0]_net_1\);
    
    \SM_BANK_SEL[14]\ : DFN1E1C0
      port map(D => N_1841, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_1_0, E => un1_REG_STATE_30, Q => 
        \SM_BANK_SEL[14]_net_1\);
    
    \ELINK_BLKA[15]\ : DFN1E0P0
      port map(D => N_65, CLK => CLK60MHZ, PRE => 
        P_USB_MASTER_EN_c_20, E => \SM_BANK_SEL[20]_net_1\, Q => 
        \ELINK_BLKA[15]_net_1\);
    
    \CHKSUM[3]\ : DFN1E1C0
      port map(D => N_1587, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_3, E => un1_REG_STATE_22, Q => 
        \CHKSUM[3]_net_1\);
    
    un1_REG_STATE_2_i : NOR2
      port map(A => un1_REG_STATE_2_i_0, B => N_1726, Y => 
        N_1562_i);
    
    \REG_ADDR_RNIP4HE[4]\ : NOR2B
      port map(A => \REG_ADDR[5]_net_1\, B => \REG_ADDR[4]_net_1\, 
        Y => N_491);
    
    \ELINK_ADDRA_11[1]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[1]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_2, E => un1_SM_BANK_SEL_16, Q => 
        \ELINK_ADDRA_11[1]_net_1\);
    
    \SM_BANK_SEL_0[21]\ : DFN1E1P0
      port map(D => N_1671, CLK => CLK60MHZ, PRE => 
        P_USB_MASTER_EN_c_2_0, E => un1_REG_STATE_30, Q => 
        \SM_BANK_SEL_0[21]_net_1\);
    
    \N_WR_USB_ADBUS_0_iv_0_RNO[4]\ : NOR2A
      port map(A => \TFC_STOP_ADDR[4]_net_1\, B => N_1501, Y => 
        \TFC_STOP_ADDR_m[4]\);
    
    USB_RXF_B_RNI21E81 : OA1C
      port map(A => \REG_STATE[2]_net_1\, B => \USB_RXF_B\, C => 
        \REG_STATE_0[3]_net_1\, Y => \REG_STATE_ns_i_a4_1_1_0[1]\);
    
    \WR_USB_ADBUS_RNO_24[1]\ : NOR2B
      port map(A => \ELINK_DOUTA_8[1]\, B => un1_SM_BANK_SEL_38, 
        Y => \ELINK_DOUTA_8_m[1]\);
    
    \REG_ADDR_RNO[4]\ : XA1B
      port map(A => \REG_ADDR[4]_net_1\, B => REG_ADDR_c3, C => 
        N_675_0, Y => REG_ADDR_n4);
    
    \WR_USB_ADBUS_RNO_4[7]\ : AO1
      port map(A => \ELINK_DOUTA_16[7]\, B => un1_SM_BANK_SEL_39, 
        C => \ELINK_DOUTA_1_m[7]\, Y => 
        \N_WR_USB_ADBUS_0_iv_9[7]\);
    
    \ELINK_DINA_2[2]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[2]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_9, E => un1_SM_BANK_SEL_5, Q => 
        \ELINK_DINA_2[2]_net_1\);
    
    USB_RXF_B_RNIKSCQ_0 : NOR2
      port map(A => \USB_RXF_B\, B => \REG_STATE[4]_net_1\, Y => 
        N_TFC_STRT_ADDR_T_0_sqmuxa_0_a2_0);
    
    \N_TFC_ADDRA_0_o2_RNO[7]\ : AO1
      port map(A => N_433_1, B => N_260, C => N_428, Y => 
        \N_TFC_ADDRA_0_o2_0[7]\);
    
    \REG_STATE_RNIVGQN[0]\ : XOR2
      port map(A => \REG_STATE[3]_net_1\, B => 
        \REG_STATE[0]_net_1\, Y => N_2628);
    
    \ELINK_DINA_0[6]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[6]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_5, E => un1_SM_BANK_SEL_6, Q => 
        \ELINK_DINA_0[6]_net_1\);
    
    USB_TXE_B_RNILBLU : NOR2B
      port map(A => N_2602, B => \USB_TXE_B\, Y => N_2606);
    
    \ELINK_BLKA_RNO_0[18]\ : AO1D
      port map(A => \N_ELINK_RWA_0_iv_0_o2_0[18]\, B => N_624_15, 
        C => \ELINK_BLKA[18]_net_1\, Y => N_63_tz);
    
    \SM_BANK_SEL_RNINT4B[18]\ : OR2
      port map(A => \SM_BANK_SEL[18]_net_1\, B => 
        \SM_BANK_SEL_0[21]_net_1\, Y => un1_SM_BANK_SEL_19);
    
    \N_WR_USB_ADBUS_0_iv_0_RNO[0]\ : NOR2A
      port map(A => \TFC_STOP_ADDR[0]_net_1\, B => N_1501, Y => 
        \TFC_STOP_ADDR_m[0]\);
    
    \TFC_STOP_ADDR_T[2]\ : DFN1E1C0
      port map(D => \RD_USB_ADBUS[2]_net_1\, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_15, E => N_TFC_STOP_ADDR_T_0_sqmuxa, 
        Q => \TFC_STOP_ADDR_T[2]_net_1\);
    
    \SM_BANK_SEL_RNI7HK1[17]\ : OR2
      port map(A => \SM_BANK_SEL[17]_net_1\, B => 
        \SM_BANK_SEL[21]_net_1\, Y => un1_SM_BANK_SEL_5);
    
    \WR_USB_ADBUS_RNO_1[4]\ : OR3
      port map(A => \N_WR_USB_ADBUS_0_iv_8[4]\, B => 
        \N_WR_USB_ADBUS_0_iv_7[4]\, C => 
        \N_WR_USB_ADBUS_0_iv_17[4]\, Y => 
        \N_WR_USB_ADBUS_0_iv_23[4]\);
    
    \SM_BANK_SEL[20]\ : DFN1E1C0
      port map(D => un1_N_ELK_N_ACTIVE_2_sqmuxa, CLK => CLK60MHZ, 
        CLR => P_USB_MASTER_EN_c_1_0, E => un1_REG_STATE_30, Q
         => \SM_BANK_SEL[20]_net_1\);
    
    \REG_STATE_RNI1SN31[5]\ : NOR2B
      port map(A => N_1710_i_0, B => \REG_STATE[5]_net_1\, Y => 
        N_427);
    
    \WR_USB_ADBUS_RNO_17[4]\ : NOR2B
      port map(A => \ELINK_DOUTA_7[4]\, B => un1_SM_BANK_SEL_37, 
        Y => \ELINK_DOUTA_7_m[4]\);
    
    \WR_USB_ADBUS_RNO_3[3]\ : AO1
      port map(A => \ELINK_DOUTA_17[3]\, B => un1_SM_BANK_SEL_40, 
        C => \ELINK_DOUTA_2_m[3]\, Y => 
        \N_WR_USB_ADBUS_0_iv_10[3]\);
    
    \WR_USB_ADBUS_RNO_23[2]\ : NOR2B
      port map(A => \ELINK_DOUTA_7[2]\, B => un1_SM_BANK_SEL_37, 
        Y => \ELINK_DOUTA_7_m[2]\);
    
    \WR_USB_ADBUS_RNO_17[2]\ : AO1
      port map(A => \CHKSUM[2]_net_1\, B => un1_REG_STATE_4, C
         => \N_WR_USB_ADBUS_0_iv_3[2]\, Y => 
        \N_WR_USB_ADBUS_0_iv_5[2]\);
    
    \WR_USB_ADBUS_RNO_10[7]\ : AO1
      port map(A => \ELINK_DOUTA_6[7]\, B => un1_SM_BANK_SEL_30, 
        C => \ELINK_DOUTA_8_m[7]\, Y => 
        \N_WR_USB_ADBUS_0_iv_13[7]\);
    
    \WR_USB_ADBUS_RNO_12[3]\ : NOR2B
      port map(A => \ELINK_DOUTA_2[3]\, B => un1_SM_BANK_SEL_32, 
        Y => \ELINK_DOUTA_2_m[3]\);
    
    \REG_STATE_0_RNIIQR51[3]\ : NOR2B
      port map(A => N_2477_i, B => \REG_STATE_0[3]_net_1\, Y => 
        N_417);
    
    \SM_BANK_SEL_RNI696G[8]\ : OR2
      port map(A => \SM_BANK_SEL[8]_net_1\, B => 
        \SM_BANK_SEL_0[21]_net_1\, Y => un1_SM_BANK_SEL_16);
    
    \SM_BANK_SEL_RNI1AJ1[12]\ : OR2
      port map(A => \SM_BANK_SEL[12]_net_1\, B => 
        \SM_BANK_SEL[11]_net_1\, Y => N_616_4);
    
    \ELINK_DINA_16[4]\ : DFN1E0C0
      port map(D => \N_TFC_DINA[4]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_18, E => N_200, Q => 
        \ELINK_DINA_16[4]_net_1\);
    
    \REG_STATE_ns_i_i_o2_1_RNO_0[0]\ : OA1
      port map(A => N_441, B => N_440, C => 
        \REG_STATE_ns_i_i_a2_1_0[0]\, Y => N_443);
    
    \REG_STATE_RNISQSJ1[1]\ : OR2
      port map(A => N_1879_1, B => N_2462, Y => N_346);
    
    \SM_BANK_SEL_RNIH21C2[7]\ : NOR3A
      port map(A => \SM_BANK_SEL[7]_net_1\, B => N_312_0, C => 
        N_1566_i_i_0, Y => un1_SM_BANK_SEL_33);
    
    USB_RD_BI_RNO_10 : XA1A
      port map(A => \REG_STATE_0[3]_net_1\, B => \USB_RXF_B_0\, C
         => \REG_STATE_0[1]_net_1\, Y => un1_REG_STATE_40_i_a2_0);
    
    \REG_STATE_0_RNI149EV[0]\ : AO1
      port map(A => N_2592, B => \REG_STATE_ns_i_1_tz[3]\, C => 
        N_2561, Y => \REG_STATE_ns_i_0[3]\);
    
    \ELINK_ADDRA_8[2]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[2]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_8, E => un1_SM_BANK_SEL_21, Q => 
        \ELINK_ADDRA_8[2]_net_1\);
    
    \WR_USB_ADBUS_RNO_12[0]\ : NOR2B
      port map(A => \ELINK_DOUTA_11[0]\, B => un1_SM_BANK_SEL_26, 
        Y => \ELINK_DOUTA_11_m[0]\);
    
    \WR_USB_ADBUS_RNO[4]\ : OR3
      port map(A => \N_WR_USB_ADBUS_0_iv_24[4]\, B => 
        \N_WR_USB_ADBUS_0_iv_23[4]\, C => 
        \N_WR_USB_ADBUS_0_iv_25[4]\, Y => \N_WR_USB_ADBUS[4]\);
    
    \REG_STATE_0_RNIO7N96[0]\ : OR3
      port map(A => N_415, B => N_418, C => 
        \REG_STATE_ns_i_i_o2_10_0[2]\, Y => 
        \REG_STATE_ns_i_i_o2_10_2[2]\);
    
    \RD_XFER_TYPE_RNINJMR_0[0]\ : NOR2A
      port map(A => \RD_XFER_TYPE[1]_net_1\, B => 
        \RD_XFER_TYPE[0]_net_1\, Y => N_1368_i_i_a5_0);
    
    \OP_MODE_T[4]\ : DFN1E1C0
      port map(D => \RD_USB_ADBUS[4]_net_1\, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_17, E => N_OP_MODE_T_0_sqmuxa, Q
         => \OP_MODE_T[4]_net_1\);
    
    \WR_USB_ADBUS_RNO_4[3]\ : AO1
      port map(A => \ELINK_DOUTA_16[3]\, B => un1_SM_BANK_SEL_39, 
        C => \ELINK_DOUTA_1_m[3]\, Y => 
        \N_WR_USB_ADBUS_0_iv_9[3]\);
    
    \WR_USB_ADBUS_RNO_18[4]\ : NOR2B
      port map(A => \ELINK_DOUTA_5[4]\, B => un1_SM_BANK_SEL_35, 
        Y => \ELINK_DOUTA_5_m[4]\);
    
    \ELINK_ADDRA_5[6]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[6]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_3, E => un1_SM_BANK_SEL_15, Q => 
        \ELINK_ADDRA_5[6]_net_1\);
    
    \TFC_STOP_ADDR_T[7]\ : DFN1E1C0
      port map(D => \RD_USB_ADBUS[7]_net_1\, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_15, E => N_TFC_STOP_ADDR_T_0_sqmuxa, 
        Q => \TFC_STOP_ADDR_T[7]_net_1\);
    
    U109_PATT_ELINK_BLK : DPRT_512X9_SRAM_9
      port map(ELINK_RWA_0 => \ELINK_RWA[9]_net_1\, 
        ELK_RX_SER_WORD_9(7) => ELK_RX_SER_WORD_9(7), 
        ELK_RX_SER_WORD_9(6) => ELK_RX_SER_WORD_9(6), 
        ELK_RX_SER_WORD_9(5) => ELK_RX_SER_WORD_9(5), 
        ELK_RX_SER_WORD_9(4) => ELK_RX_SER_WORD_9(4), 
        ELK_RX_SER_WORD_9(3) => ELK_RX_SER_WORD_9(3), 
        ELK_RX_SER_WORD_9(2) => ELK_RX_SER_WORD_9(2), 
        ELK_RX_SER_WORD_9(1) => ELK_RX_SER_WORD_9(1), 
        ELK_RX_SER_WORD_9(0) => ELK_RX_SER_WORD_9(0), 
        ELINK_DINA_9(7) => \ELINK_DINA_9[7]_net_1\, 
        ELINK_DINA_9(6) => \ELINK_DINA_9[6]_net_1\, 
        ELINK_DINA_9(5) => \ELINK_DINA_9[5]_net_1\, 
        ELINK_DINA_9(4) => \ELINK_DINA_9[4]_net_1\, 
        ELINK_DINA_9(3) => \ELINK_DINA_9[3]_net_1\, 
        ELINK_DINA_9(2) => \ELINK_DINA_9[2]_net_1\, 
        ELINK_DINA_9(1) => \ELINK_DINA_9[1]_net_1\, 
        ELINK_DINA_9(0) => \ELINK_DINA_9[0]_net_1\, ELINK_BLKA_0
         => \ELINK_BLKA[9]_net_1\, ELKS_ADDRB(7) => ELKS_ADDRB(7), 
        ELKS_ADDRB(6) => ELKS_ADDRB(6), ELKS_ADDRB(5) => 
        ELKS_ADDRB(5), ELKS_ADDRB(4) => ELKS_ADDRB(4), 
        ELKS_ADDRB(3) => ELKS_ADDRB(3), ELKS_ADDRB(2) => 
        ELKS_ADDRB(2), ELKS_ADDRB(1) => ELKS_ADDRB(1), 
        ELKS_ADDRB(0) => ELKS_ADDRB(0), ELINK_ADDRA_9(7) => 
        \ELINK_ADDRA_9[7]_net_1\, ELINK_ADDRA_9(6) => 
        \ELINK_ADDRA_9[6]_net_1\, ELINK_ADDRA_9(5) => 
        \ELINK_ADDRA_9[5]_net_1\, ELINK_ADDRA_9(4) => 
        \ELINK_ADDRA_9[4]_net_1\, ELINK_ADDRA_9(3) => 
        \ELINK_ADDRA_9[3]_net_1\, ELINK_ADDRA_9(2) => 
        \ELINK_ADDRA_9[2]_net_1\, ELINK_ADDRA_9(1) => 
        \ELINK_ADDRA_9[1]_net_1\, ELINK_ADDRA_9(0) => 
        \ELINK_ADDRA_9[0]_net_1\, PATT_ELK_DAT_9(7) => 
        PATT_ELK_DAT_9(7), PATT_ELK_DAT_9(6) => PATT_ELK_DAT_9(6), 
        PATT_ELK_DAT_9(5) => PATT_ELK_DAT_9(5), PATT_ELK_DAT_9(4)
         => PATT_ELK_DAT_9(4), PATT_ELK_DAT_9(3) => 
        PATT_ELK_DAT_9(3), PATT_ELK_DAT_9(2) => PATT_ELK_DAT_9(2), 
        PATT_ELK_DAT_9(1) => PATT_ELK_DAT_9(1), PATT_ELK_DAT_9(0)
         => PATT_ELK_DAT_9(0), ELINK_DOUTA_9(7) => 
        \ELINK_DOUTA_9[7]\, ELINK_DOUTA_9(6) => 
        \ELINK_DOUTA_9[6]\, ELINK_DOUTA_9(5) => 
        \ELINK_DOUTA_9[5]\, ELINK_DOUTA_9(4) => 
        \ELINK_DOUTA_9[4]\, ELINK_DOUTA_9(3) => 
        \ELINK_DOUTA_9[3]\, ELINK_DOUTA_9(2) => 
        \ELINK_DOUTA_9[2]\, ELINK_DOUTA_9(1) => 
        \ELINK_DOUTA_9[1]\, ELINK_DOUTA_9(0) => 
        \ELINK_DOUTA_9[0]\, ELKS_RWB => ELKS_RWB, 
        P_USB_MASTER_EN_c_0 => P_USB_MASTER_EN_c_0, CLK_40M_GL
         => CLK_40M_GL, CLK60MHZ => CLK60MHZ, ELKS_RAM_BLKB_EN
         => ELKS_RAM_BLKB_EN);
    
    \WR_USB_ADBUS_RNO_0[5]\ : OR3
      port map(A => \N_WR_USB_ADBUS_0_iv_10[5]\, B => 
        \N_WR_USB_ADBUS_0_iv_9[5]\, C => 
        \N_WR_USB_ADBUS_0_iv_20[5]\, Y => 
        \N_WR_USB_ADBUS_0_iv_24[5]\);
    
    \ELINK_ADDRA_17[6]\ : DFN1E0C0
      port map(D => \N_TFC_ADDRA[6]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_11, E => N_197, Q => 
        \ELINK_ADDRA_17[6]_net_1\);
    
    \WR_USB_ADBUS_RNO_3[6]\ : AO1
      port map(A => \ELINK_DOUTA_17[6]\, B => un1_SM_BANK_SEL_40, 
        C => \ELINK_DOUTA_18_m[6]\, Y => 
        \N_WR_USB_ADBUS_0_iv_9[6]\);
    
    \REG_ADDR[5]\ : DFN1E1C0
      port map(D => REG_ADDR_n5, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_10, E => REG_ADDRe, Q => 
        \REG_ADDR[5]_net_1\);
    
    \RD_USB_ADBUS_RNIOEOG3[7]\ : OR2
      port map(A => N_1702, B => N_1700, Y => N_1717);
    
    \REG_STATE_ns_i_i_a2_0[0]\ : NOR2A
      port map(A => \REG_STATE_ns_i_i_a2_0_2[0]_net_1\, B => 
        N_275, Y => N_421);
    
    \WR_USB_ADBUS_RNO_14[6]\ : NOR2B
      port map(A => \ELINK_DOUTA_8[6]\, B => un1_SM_BANK_SEL_38, 
        Y => \ELINK_DOUTA_8_m[6]\);
    
    \RD_USB_ADBUS_RNIL9IK2[0]\ : NOR2A
      port map(A => \RD_USB_ADBUS[0]_net_1\, B => N_206, Y => 
        \N_TFC_DINA[0]\);
    
    \ELINK_BLKA_RNO_0[7]\ : OA1B
      port map(A => N_616_16, B => \N_ELINK_RWA_3[7]\, C => 
        \ELINK_BLKA[7]_net_1\, Y => \ELINK_BLKA_i_m[7]\);
    
    \WR_USB_ADBUS_RNO_29[5]\ : NOR2B
      port map(A => \ELINK_DOUTA_5[5]\, B => un1_SM_BANK_SEL_35, 
        Y => \ELINK_DOUTA_5_m[5]\);
    
    \SM_BANK_SEL_RNI35MB[3]\ : NOR2
      port map(A => \SM_BANK_SEL[3]_net_1\, B => 
        \SM_BANK_SEL[4]_net_1\, Y => N_462);
    
    \OP_MODE[7]\ : DFN1E1C0
      port map(D => \OP_MODE_T[7]_net_1\, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_15, E => \REG_STATE_d[30]\, Q => 
        \OP_MODE[7]_net_1\);
    
    \WR_USB_ADBUS_RNO_31[5]\ : NOR3B
      port map(A => N_1352_1, B => \OP_MODE[5]_net_1\, C => 
        REG_STATE_s20_i_0, Y => \OP_MODE_m[5]\);
    
    \WR_USB_ADBUS_RNO_5[5]\ : OR3
      port map(A => \ELINK_DOUTA_3_m[5]\, B => 
        \ELINK_DOUTA_18_m[5]\, C => \N_WR_USB_ADBUS_0_iv_12[5]\, 
        Y => \N_WR_USB_ADBUS_0_iv_20[5]\);
    
    \RD_USB_ADBUS_RNI38BJ[4]\ : OR2A
      port map(A => \RD_USB_ADBUS[5]_net_1\, B => 
        \RD_USB_ADBUS[4]_net_1\, Y => N_293);
    
    \REG_STATE_0_RNISQSJ1[1]\ : NOR3A
      port map(A => \REG_STATE_0[1]_net_1\, B => 
        \REG_STATE_0[2]_net_1\, C => N_312, Y => 
        \REG_STATE_ns_i_a4_9_1[4]\);
    
    \RD_USB_ADBUS_RNIV3BJ[3]\ : OR2
      port map(A => \RD_USB_ADBUS[3]_net_1\, B => 
        \RD_USB_ADBUS[2]_net_1\, Y => N_1700);
    
    \ELINK_RWA[1]\ : DFN1E0P0
      port map(D => \N_ELINK_RWA_0_iv[1]\, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_6, E => \SM_BANK_SEL_0[20]_net_1\, 
        Q => \ELINK_RWA[1]_net_1\);
    
    \CHKSUM_RNO[1]\ : NOR2A
      port map(A => \RD_USB_ADBUS[1]_net_1\, B => N_675, Y => 
        N_236);
    
    \ELINK_DINA_17[6]\ : DFN1E0C0
      port map(D => \N_TFC_DINA[6]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_19, E => N_197, Q => 
        \ELINK_DINA_17[6]_net_1\);
    
    \WR_USB_ADBUS_RNO_3[5]\ : AO1
      port map(A => \ELINK_DOUTA_17[5]\, B => un1_SM_BANK_SEL_40, 
        C => \ELINK_DOUTA_2_m[5]\, Y => 
        \N_WR_USB_ADBUS_0_iv_10[5]\);
    
    \WR_XFER_TYPE[7]\ : DFN1C0
      port map(D => \WR_XFER_TYPE_RNO[7]_net_1\, CLK => CLK60MHZ, 
        CLR => P_USB_MASTER_EN_c, Q => \WR_XFER_TYPE[7]_net_1\);
    
    \SM_BANK_SEL_RNITMN22[10]\ : NOR3A
      port map(A => \SM_BANK_SEL[10]_net_1\, B => N_312, C => 
        N_1566_i_i_0, Y => un1_SM_BANK_SEL_42);
    
    \N_WR_USB_ADBUS_0_iv_0[0]\ : OR2
      port map(A => \TFC_STOP_ADDR_m[0]\, B => N_1562_i, Y => 
        \N_WR_USB_ADBUS_0_iv_0[0]_net_1\);
    
    \ELINK_DINA_2[0]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[0]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_9, E => un1_SM_BANK_SEL_5, Q => 
        \ELINK_DINA_2[0]_net_1\);
    
    \REG_STATE_0_RNICKR51[1]\ : OR2A
      port map(A => \REG_STATE_0[1]_net_1\, B => N_2497, Y => 
        N_1765);
    
    \ELINK_ADDRA_10[1]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[1]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_22, E => un1_SM_BANK_SEL_20, Q => 
        \ELINK_ADDRA_10[1]_net_1\);
    
    \SM_BANK_SEL_RNIHT4J[10]\ : NOR2B
      port map(A => N_469, B => N_461, Y => N_486);
    
    \ELINK_DINA_11[2]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[2]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_11, E => un1_SM_BANK_SEL_16, Q => 
        \ELINK_DINA_11[2]_net_1\);
    
    \WR_USB_ADBUS_RNO_27[5]\ : NOR2B
      port map(A => \ELINK_DOUTA_10[5]\, B => un1_SM_BANK_SEL_34, 
        Y => \ELINK_DOUTA_10_m[5]\);
    
    USB_TXE_B_RNIJIIA1 : NOR2B
      port map(A => \USB_TXE_B\, B => N_2616, Y => 
        \REG_STATE_ns_i_a4_8_0[1]\);
    
    \REG_STATE_ns_i_i_o2_1[0]\ : OR2
      port map(A => N_444, B => N_443, Y => N_275);
    
    \WR_USB_ADBUS_RNO_11[1]\ : OR3
      port map(A => \ELINK_DOUTA_11_m[1]\, B => 
        \ELINK_DOUTA_10_m[1]\, C => \N_WR_USB_ADBUS_0_iv_16[1]\, 
        Y => \N_WR_USB_ADBUS_0_iv_22[1]\);
    
    \RD_XFER_TYPE_RNI30NR[6]\ : OR2
      port map(A => \RD_XFER_TYPE[7]_net_1\, B => 
        \RD_XFER_TYPE[6]_net_1\, Y => N_1367_i_i_o2_0_1);
    
    USB_RD_BI_RNO_11 : NOR3C
      port map(A => \REG_STATE_0[1]_net_1\, B => 
        \RD_USB_ADBUS[7]_net_1\, C => N_1352_5, Y => 
        N_USB_RD_BI_i_a2_4_1);
    
    \ELINK_ADDRA_2[4]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[4]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_21, E => un1_SM_BANK_SEL_5, Q => 
        \ELINK_ADDRA_2[4]_net_1\);
    
    \RD_USB_ADBUS_RNIRVAJ_2[0]\ : NOR2A
      port map(A => \RD_USB_ADBUS[0]_net_1\, B => 
        \RD_USB_ADBUS[1]_net_1\, Y => N_1351_4);
    
    \ELINK_RWA[17]\ : DFN1E0P0
      port map(D => \N_ELINK_RWA_0_iv[17]\, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_12, E => \SM_BANK_SEL_0[20]_net_1\, 
        Q => \ELINK_RWA[17]_net_1\);
    
    \WR_USB_ADBUS_RNO_24[2]\ : AO1
      port map(A => \WR_XFER_TYPE[2]_net_1\, B => N_398, C => 
        \ELINKS_STOP_ADDR_m[2]\, Y => \N_WR_USB_ADBUS_0_iv_3[2]\);
    
    \ELINK_RWA_RNO_0[14]\ : OA1B
      port map(A => N_624_15, B => \N_ELINK_RWA_3[14]\, C => 
        \ELINK_RWA[14]_net_1\, Y => \ELINK_RWA_i_m[14]\);
    
    \WR_USB_ADBUS_RNO_13[4]\ : NOR2B
      port map(A => \ELINK_DOUTA_9[4]\, B => un1_SM_BANK_SEL_42, 
        Y => \ELINK_DOUTA_9_m[4]\);
    
    U118_PATT_ELINK_BLK : DPRT_512X9_SRAM_18
      port map(ELINK_RWA_0 => \ELINK_RWA[18]_net_1\, 
        ELK_RX_SER_WORD_18(7) => ELK_RX_SER_WORD_18(7), 
        ELK_RX_SER_WORD_18(6) => ELK_RX_SER_WORD_18(6), 
        ELK_RX_SER_WORD_18(5) => ELK_RX_SER_WORD_18(5), 
        ELK_RX_SER_WORD_18(4) => ELK_RX_SER_WORD_18(4), 
        ELK_RX_SER_WORD_18(3) => ELK_RX_SER_WORD_18(3), 
        ELK_RX_SER_WORD_18(2) => ELK_RX_SER_WORD_18(2), 
        ELK_RX_SER_WORD_18(1) => ELK_RX_SER_WORD_18(1), 
        ELK_RX_SER_WORD_18(0) => ELK_RX_SER_WORD_18(0), 
        ELINK_DINA_18(7) => \ELINK_DINA_18[7]_net_1\, 
        ELINK_DINA_18(6) => \ELINK_DINA_18[6]_net_1\, 
        ELINK_DINA_18(5) => \ELINK_DINA_18[5]_net_1\, 
        ELINK_DINA_18(4) => \ELINK_DINA_18[4]_net_1\, 
        ELINK_DINA_18(3) => \ELINK_DINA_18[3]_net_1\, 
        ELINK_DINA_18(2) => \ELINK_DINA_18[2]_net_1\, 
        ELINK_DINA_18(1) => \ELINK_DINA_18[1]_net_1\, 
        ELINK_DINA_18(0) => \ELINK_DINA_18[0]_net_1\, 
        ELINK_BLKA_0 => \ELINK_BLKA[18]_net_1\, ELKS_ADDRB_0_d0
         => ELKS_ADDRB(0), ELKS_ADDRB_1 => ELKS_ADDRB(1), 
        ELKS_ADDRB_3 => ELKS_ADDRB(3), ELKS_ADDRB_5 => 
        ELKS_ADDRB(5), ELKS_ADDRB_7 => ELKS_ADDRB(7), 
        ELKS_ADDRB_0_0 => ELKS_ADDRB_0_0, ELKS_ADDRB_0_2 => 
        ELKS_ADDRB_0_2, ELKS_ADDRB_0_4 => ELKS_ADDRB_0_4, 
        ELINK_ADDRA_18(7) => \ELINK_ADDRA_18[7]_net_1\, 
        ELINK_ADDRA_18(6) => \ELINK_ADDRA_18[6]_net_1\, 
        ELINK_ADDRA_18(5) => \ELINK_ADDRA_18[5]_net_1\, 
        ELINK_ADDRA_18(4) => \ELINK_ADDRA_18[4]_net_1\, 
        ELINK_ADDRA_18(3) => \ELINK_ADDRA_18[3]_net_1\, 
        ELINK_ADDRA_18(2) => \ELINK_ADDRA_18[2]_net_1\, 
        ELINK_ADDRA_18(1) => \ELINK_ADDRA_18[1]_net_1\, 
        ELINK_ADDRA_18(0) => \ELINK_ADDRA_18[0]_net_1\, 
        PATT_ELK_DAT_18(7) => PATT_ELK_DAT_18(7), 
        PATT_ELK_DAT_18(6) => PATT_ELK_DAT_18(6), 
        PATT_ELK_DAT_18(5) => PATT_ELK_DAT_18(5), 
        PATT_ELK_DAT_18(4) => PATT_ELK_DAT_18(4), 
        PATT_ELK_DAT_18(3) => PATT_ELK_DAT_18(3), 
        PATT_ELK_DAT_18(2) => PATT_ELK_DAT_18(2), 
        PATT_ELK_DAT_18(1) => PATT_ELK_DAT_18(1), 
        PATT_ELK_DAT_18(0) => PATT_ELK_DAT_18(0), 
        ELINK_DOUTA_18(7) => \ELINK_DOUTA_18[7]\, 
        ELINK_DOUTA_18(6) => \ELINK_DOUTA_18[6]\, 
        ELINK_DOUTA_18(5) => \ELINK_DOUTA_18[5]\, 
        ELINK_DOUTA_18(4) => \ELINK_DOUTA_18[4]\, 
        ELINK_DOUTA_18(3) => \ELINK_DOUTA_18[3]\, 
        ELINK_DOUTA_18(2) => \ELINK_DOUTA_18[2]\, 
        ELINK_DOUTA_18(1) => \ELINK_DOUTA_18[1]\, 
        ELINK_DOUTA_18(0) => \ELINK_DOUTA_18[0]\, ELKS_RWB => 
        ELKS_RWB, P_USB_MASTER_EN_c_0 => P_USB_MASTER_EN_c_0, 
        CLK_40M_GL => CLK_40M_GL, CLK60MHZ => CLK60MHZ, 
        ELKS_RAM_BLKB_EN => ELKS_RAM_BLKB_EN);
    
    \REG_STATE_RNIB6E34[2]\ : OR3
      port map(A => \REG_STATE_ns_i_a4_3_0[3]\, B => 
        \REG_STATE_ns_i_1_tz_0[3]\, C => 
        \REG_STATE_ns_i_1_tz_1[3]\, Y => \REG_STATE_ns_i_1_tz[3]\);
    
    \ELINKS_STRT_ADDR[5]\ : DFN1E1C0
      port map(D => \ELINKS_STRT_ADDR_T[5]_net_1\, CLK => 
        CLK60MHZ, CLR => P_USB_MASTER_EN_c_17, E => 
        \REG_STATE_d[30]\, Q => \ELINKS_STRT_ADDR[5]_net_1\);
    
    \RD_XFER_TYPE_RNO_0[6]\ : NOR2A
      port map(A => \RD_USB_ADBUS[6]_net_1\, B => N_1694, Y => 
        N_1806);
    
    \ELINK_ADDRA_15[7]\ : DFN1E0C0
      port map(D => \N_TFC_ADDRA[7]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_6, E => N_199, Q => 
        \ELINK_ADDRA_15[7]_net_1\);
    
    \REG_STATE_ns_i_i_o2_6_1_RNO_4[0]\ : NOR3A
      port map(A => N_2462, B => N_252, C => N_268, Y => N_452);
    
    \ELINK_DINA_2[7]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[7]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_9, E => un1_SM_BANK_SEL_5, Q => 
        \ELINK_DINA_2[7]_net_1\);
    
    \WR_USB_ADBUS_RNO_34[5]\ : NOR2A
      port map(A => \ELINKS_STRT_ADDR[5]_net_1\, B => N_1499, Y
         => \ELINKS_STRT_ADDR_m[5]\);
    
    USB_RXF_B_RNIJ4CL3 : AO1
      port map(A => \REG_STATE_ns_i_a4_1_1_0[1]\, B => N_1879_1, 
        C => \REG_STATE_ns_i_a4_10_0[1]\, Y => 
        REG_STATE_ns_i_245_tz_0);
    
    \ELINK_DINA_9[7]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[7]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_20, E => un1_SM_BANK_SEL_9, Q => 
        \ELINK_DINA_9[7]_net_1\);
    
    \WR_USB_ADBUS_RNO_29[2]\ : NOR2B
      port map(A => \ELINK_DOUTA_12[2]\, B => un1_SM_BANK_SEL_33, 
        Y => \ELINK_DOUTA_12_m[2]\);
    
    \REG_STATE_0_RNIDLR51[3]\ : OR2
      port map(A => N_1359_1, B => \REG_STATE_0[3]_net_1\, Y => 
        N_2515);
    
    \WR_XFER_TYPE_RNIUDSS[0]\ : NOR2A
      port map(A => \WR_XFER_TYPE[0]_net_1\, B => 
        \WR_XFER_TYPE[2]_net_1\, Y => REG_STATE_tr67_0);
    
    \REG_STATE_0_RNI8PBS2[4]\ : AO1C
      port map(A => \REG_STATE_0[4]_net_1\, B => N_470, C => 
        N_256, Y => \REG_STATE_ns_i_i_o2_10_3[2]\);
    
    \ELINK_RWA_RNO_0[5]\ : OA1B
      port map(A => N_616_16, B => \N_ELINK_RWA_3[5]\, C => 
        \ELINK_RWA[5]_net_1\, Y => N_183);
    
    \ELINK_DINA_18[7]\ : DFN1E0C0
      port map(D => \N_TFC_DINA[7]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_21, E => N_198, Q => 
        \ELINK_DINA_18[7]_net_1\);
    
    \ELINK_DINA_14[7]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[7]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_16, E => un1_SM_BANK_SEL_1, Q => 
        \ELINK_DINA_14[7]_net_1\);
    
    \WR_USB_ADBUS_RNO_20[5]\ : NOR2A
      port map(A => \TFC_DOUTA[5]\, B => N_243, Y => 
        \TFC_DOUTA_m[5]\);
    
    \REG_ADDR_RNILQCP[2]\ : NOR3B
      port map(A => N_261, B => \REG_ADDR[2]_net_1\, C => 
        \SM_BANK_SEL_0[21]_net_1\, Y => \N_TFC_ADDRA[2]\);
    
    \SM_BANK_SEL[2]\ : DFN1E1C0
      port map(D => N_1840, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_7, E => un1_REG_STATE_30, Q => 
        \SM_BANK_SEL[2]_net_1\);
    
    \ELINK_DINA_10[6]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[6]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_9, E => un1_SM_BANK_SEL_20, Q => 
        \ELINK_DINA_10[6]_net_1\);
    
    \SM_BANK_SEL_RNIPB73[15]\ : OR3
      port map(A => \SM_BANK_SEL[15]_net_1\, B => 
        \SM_BANK_SEL[17]_net_1\, C => N_618_1, Y => 
        \N_ELINK_RWA_1[3]\);
    
    \REG_STATE_RNI2KQN[4]\ : NOR2A
      port map(A => \REG_STATE[4]_net_1\, B => 
        \REG_STATE[2]_net_1\, Y => N_2477_i);
    
    \WR_USB_ADBUS_RNO_28[3]\ : NOR2B
      port map(A => \ELINK_DOUTA_5[3]\, B => un1_SM_BANK_SEL_35, 
        Y => \ELINK_DOUTA_5_m[3]\);
    
    \REG_STATE_RNIVGQN_3[0]\ : NOR2B
      port map(A => \REG_STATE[0]_net_1\, B => 
        \REG_STATE[3]_net_1\, Y => N_2571_1);
    
    \REG_ADDR_RNO_0[8]\ : NOR2B
      port map(A => \REG_ADDR[7]_net_1\, B => REG_ADDR_c6, Y => 
        REG_ADDR_75_0);
    
    \ELINK_ADDRA_13[1]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[1]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_3, E => un1_SM_BANK_SEL_2, Q => 
        \ELINK_ADDRA_13[1]_net_1\);
    
    USB_TXE_B : DFN1P0
      port map(D => P_USB_TXE_B_c, CLK => CLK60MHZ, PRE => 
        P_USB_MASTER_EN_c_22, Q => \USB_TXE_B\);
    
    U115_PATT_ELINK_BLK : DPRT_512X9_SRAM_15
      port map(ELINK_RWA_0 => \ELINK_RWA[15]_net_1\, 
        ELK_RX_SER_WORD_15(7) => ELK_RX_SER_WORD_15(7), 
        ELK_RX_SER_WORD_15(6) => ELK_RX_SER_WORD_15(6), 
        ELK_RX_SER_WORD_15(5) => ELK_RX_SER_WORD_15(5), 
        ELK_RX_SER_WORD_15(4) => ELK_RX_SER_WORD_15(4), 
        ELK_RX_SER_WORD_15(3) => ELK_RX_SER_WORD_15(3), 
        ELK_RX_SER_WORD_15(2) => ELK_RX_SER_WORD_15(2), 
        ELK_RX_SER_WORD_15(1) => ELK_RX_SER_WORD_15(1), 
        ELK_RX_SER_WORD_15(0) => ELK_RX_SER_WORD_15(0), 
        ELINK_DINA_15(7) => \ELINK_DINA_15[7]_net_1\, 
        ELINK_DINA_15(6) => \ELINK_DINA_15[6]_net_1\, 
        ELINK_DINA_15(5) => \ELINK_DINA_15[5]_net_1\, 
        ELINK_DINA_15(4) => \ELINK_DINA_15[4]_net_1\, 
        ELINK_DINA_15(3) => \ELINK_DINA_15[3]_net_1\, 
        ELINK_DINA_15(2) => \ELINK_DINA_15[2]_net_1\, 
        ELINK_DINA_15(1) => \ELINK_DINA_15[1]_net_1\, 
        ELINK_DINA_15(0) => \ELINK_DINA_15[0]_net_1\, 
        ELINK_BLKA_0 => \ELINK_BLKA[15]_net_1\, ELKS_ADDRB(7) => 
        ELKS_ADDRB(7), ELKS_ADDRB(6) => ELKS_ADDRB(6), 
        ELKS_ADDRB(5) => ELKS_ADDRB(5), ELKS_ADDRB(4) => 
        ELKS_ADDRB(4), ELKS_ADDRB(3) => ELKS_ADDRB(3), 
        ELKS_ADDRB(2) => ELKS_ADDRB(2), ELKS_ADDRB(1) => 
        ELKS_ADDRB(1), ELKS_ADDRB(0) => ELKS_ADDRB(0), 
        ELINK_ADDRA_15(7) => \ELINK_ADDRA_15[7]_net_1\, 
        ELINK_ADDRA_15(6) => \ELINK_ADDRA_15[6]_net_1\, 
        ELINK_ADDRA_15(5) => \ELINK_ADDRA_15[5]_net_1\, 
        ELINK_ADDRA_15(4) => \ELINK_ADDRA_15[4]_net_1\, 
        ELINK_ADDRA_15(3) => \ELINK_ADDRA_15[3]_net_1\, 
        ELINK_ADDRA_15(2) => \ELINK_ADDRA_15[2]_net_1\, 
        ELINK_ADDRA_15(1) => \ELINK_ADDRA_15[1]_net_1\, 
        ELINK_ADDRA_15(0) => \ELINK_ADDRA_15[0]_net_1\, 
        PATT_ELK_DAT_15(7) => PATT_ELK_DAT_15(7), 
        PATT_ELK_DAT_15(6) => PATT_ELK_DAT_15(6), 
        PATT_ELK_DAT_15(5) => PATT_ELK_DAT_15(5), 
        PATT_ELK_DAT_15(4) => PATT_ELK_DAT_15(4), 
        PATT_ELK_DAT_15(3) => PATT_ELK_DAT_15(3), 
        PATT_ELK_DAT_15(2) => PATT_ELK_DAT_15(2), 
        PATT_ELK_DAT_15(1) => PATT_ELK_DAT_15(1), 
        PATT_ELK_DAT_15(0) => PATT_ELK_DAT_15(0), 
        ELINK_DOUTA_15(7) => \ELINK_DOUTA_15[7]\, 
        ELINK_DOUTA_15(6) => \ELINK_DOUTA_15[6]\, 
        ELINK_DOUTA_15(5) => \ELINK_DOUTA_15[5]\, 
        ELINK_DOUTA_15(4) => \ELINK_DOUTA_15[4]\, 
        ELINK_DOUTA_15(3) => \ELINK_DOUTA_15[3]\, 
        ELINK_DOUTA_15(2) => \ELINK_DOUTA_15[2]\, 
        ELINK_DOUTA_15(1) => \ELINK_DOUTA_15[1]\, 
        ELINK_DOUTA_15(0) => \ELINK_DOUTA_15[0]\, ELKS_RWB => 
        ELKS_RWB, P_USB_MASTER_EN_c_0 => P_USB_MASTER_EN_c_0, 
        CLK_40M_GL => CLK_40M_GL, CLK60MHZ => CLK60MHZ, 
        ELKS_RAM_BLKB_EN => ELKS_RAM_BLKB_EN);
    
    \ELINK_DINA_7[7]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[7]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_17, E => un1_SM_BANK_SEL_12, Q => 
        \ELINK_DINA_7[7]_net_1\);
    
    \REG_STATE_0_RNIF9MT1[4]\ : OR3B
      port map(A => \REG_STATE_0[4]_net_1\, B => N_470, C => 
        \REG_STATE[2]_net_1\, Y => N_1569);
    
    \REG_STATE_0_RNIHK3A1[3]\ : OA1C
      port map(A => \REG_STATE_0[3]_net_1\, B => 
        \REG_STATE_0[5]_net_1\, C => \REG_STATE_0[2]_net_1\, Y
         => \REG_STATE_ns_i_a4_1_0[3]\);
    
    \ELINK_DINA_3[6]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[6]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_11, E => un1_SM_BANK_SEL_4, Q => 
        \ELINK_DINA_3[6]_net_1\);
    
    \REG_ADDR_RNIJOCP[0]\ : NOR3B
      port map(A => N_261, B => \REG_ADDR[0]_net_1\, C => 
        \SM_BANK_SEL_0[21]_net_1\, Y => \N_TFC_ADDRA[0]\);
    
    \WR_USB_ADBUS_RNO_16[4]\ : AO1
      port map(A => \ELINK_DOUTA_14[4]\, B => un1_SM_BANK_SEL_23, 
        C => \ELINK_DOUTA_19_m[4]\, Y => 
        \N_WR_USB_ADBUS_0_iv_12[4]\);
    
    \ELINK_RWA_RNO[1]\ : AOI1
      port map(A => \SM_BANK_SEL[18]_net_1\, B => un1_USB_RXF_B_m, 
        C => N_185, Y => \N_ELINK_RWA_0_iv[1]\);
    
    \WR_USB_ADBUS[2]\ : DFN1E0C0
      port map(D => \N_WR_USB_ADBUS[2]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_15, E => un1_REG_STATE_26, Q => 
        \WR_USB_ADBUS[2]_net_1\);
    
    \RD_XFER_TYPE_RNO_0[5]\ : NOR2A
      port map(A => \RD_USB_ADBUS[5]_net_1\, B => N_1694, Y => 
        N_1804);
    
    \ELINK_ADDRA_2[2]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[2]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_21, E => un1_SM_BANK_SEL_5, Q => 
        \ELINK_ADDRA_2[2]_net_1\);
    
    \REG_STATE_0_RNIU5QV1[4]\ : NOR3C
      port map(A => \REG_STATE_0[2]_net_1\, B => 
        \REG_STATE_0[4]_net_1\, C => N_470, Y => N_398);
    
    \CHKSUM_RNO[7]\ : NOR2A
      port map(A => \RD_USB_ADBUS[7]_net_1\, B => N_675, Y => 
        N_226);
    
    \RD_USB_ADBUS_RNIJUIL[6]\ : NOR2A
      port map(A => \REG_STATE[2]_net_1\, B => 
        \RD_USB_ADBUS[6]_net_1\, Y => un1_REG_STATE_35_i_a2_0);
    
    \ELINK_ADDRA_15[3]\ : DFN1E0C0
      port map(D => \N_TFC_ADDRA[3]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_6, E => N_199, Q => 
        \ELINK_ADDRA_15[3]_net_1\);
    
    \SM_BANK_SEL_RNIRBHA1[5]\ : NOR2B
      port map(A => N_486, B => N_477, Y => N_394);
    
    \REG_STATE_RNI0DIR1_1[4]\ : NOR2A
      port map(A => N_1710_i_0, B => N_1691, Y => N_675);
    
    ELK_N_ACTIVE_RNIS2SQ2 : OR3
      port map(A => \REG_STATE_ns_i_a2_4_0[5]\, B => 
        \REG_STATE_ns_i_a2_4_tz_tz_tz_tz[5]\, C => N_252, Y => 
        \REG_STATE_ns_i_a2_4_2[5]\);
    
    \TFC_STOP_ADDR_T[5]\ : DFN1E1C0
      port map(D => \RD_USB_ADBUS[5]_net_1\, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_15, E => N_TFC_STOP_ADDR_T_0_sqmuxa, 
        Q => \TFC_STOP_ADDR_T[5]_net_1\);
    
    \REG_STATE_0_RNI269CG[5]\ : OR3
      port map(A => N_457, B => N_456, C => 
        \REG_STATE_ns_i_i_o2_10_5[2]\, Y => N_510);
    
    \WR_USB_ADBUS_RNO_36[3]\ : NOR2B
      port map(A => \ELINK_DOUTA_13[3]\, B => un1_SM_BANK_SEL_29, 
        Y => \ELINK_DOUTA_13_m[3]\);
    
    \SI_CNT[2]\ : DFN1E1C0
      port map(D => N_44, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_5, E => SI_CNTe, Q => \SI_CNT[2]_net_1\);
    
    \SM_BANK_SEL_RNO[8]\ : NOR3A
      port map(A => N_1892, B => \RD_USB_ADBUS[2]_net_1\, C => 
        N_290, Y => N_1836);
    
    \WR_USB_ADBUS_RNO_2[5]\ : OR3
      port map(A => \N_WR_USB_ADBUS_0_iv_14[5]\, B => 
        \N_WR_USB_ADBUS_0_iv_13[5]\, C => 
        \N_WR_USB_ADBUS_0_iv_22[5]\, Y => 
        \N_WR_USB_ADBUS_0_iv_25[5]\);
    
    \RD_USB_ADBUS_RNI2CM61_0[4]\ : AOI1B
      port map(A => N_1700, B => \RD_USB_ADBUS[4]_net_1\, C => 
        \RD_USB_ADBUS[5]_net_1\, Y => 
        \REG_STATE_ns_i_i_a5_0_1_0[2]\);
    
    \ELINK_DINA_13[6]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[6]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_14, E => un1_SM_BANK_SEL_2, Q => 
        \ELINK_DINA_13[6]_net_1\);
    
    \WR_USB_ADBUS_RNO_25[1]\ : NOR2B
      port map(A => \ELINK_DOUTA_11[1]\, B => un1_SM_BANK_SEL_26, 
        Y => \ELINK_DOUTA_11_m[1]\);
    
    \ELINK_DINA_7[4]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[4]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_17, E => un1_SM_BANK_SEL_12, Q => 
        \ELINK_DINA_7[4]_net_1\);
    
    \ELINK_BLKA_RNO[10]\ : AOI1
      port map(A => \SM_BANK_SEL[9]_net_1\, B => X_BLKA_i, C => 
        \ELINK_BLKA_i_m[10]\, Y => \N_ELINK_BLKA_0_iv[10]\);
    
    \ELINK_BLKA[1]\ : DFN1E0P0
      port map(D => \N_ELINK_BLKA_0_iv[1]\, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_19, E => \SM_BANK_SEL_0[20]_net_1\, 
        Q => \ELINK_BLKA[1]_net_1\);
    
    \ELINK_DINA_14[1]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[1]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_16, E => un1_SM_BANK_SEL_1, Q => 
        \ELINK_DINA_14[1]_net_1\);
    
    \ELINK_DINA_6[7]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[7]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_16, E => un1_SM_BANK_SEL_10, Q => 
        \ELINK_DINA_6[7]_net_1\);
    
    \ELINK_ADDRA_3[1]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[1]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_1, E => un1_SM_BANK_SEL_4, Q => 
        \ELINK_ADDRA_3[1]_net_1\);
    
    \WR_USB_ADBUS_RNO_31[6]\ : NOR3B
      port map(A => N_1352_1, B => \OP_MODE[6]_net_1\, C => 
        REG_STATE_s20_i_0, Y => \OP_MODE_m[6]\);
    
    USB_OE_BI_RNO_2 : NOR3B
      port map(A => N_1352_4, B => N_1710_i_0, C => N_1695, Y => 
        N_USB_OE_BI_iv_0_i_a2_0_5);
    
    \ELINK_BLKA_RNO[14]\ : AOI1
      port map(A => \SM_BANK_SEL[5]_net_1\, B => X_BLKA_i, C => 
        \ELINK_BLKA_i_m[14]\, Y => \N_ELINK_BLKA_0_iv[14]\);
    
    USB_RD_BI_RNO_3 : NOR2B
      port map(A => N_1713, B => \REG_STATE[4]_net_1\, Y => 
        N_1867);
    
    \OP_MODE_T[5]\ : DFN1E1C0
      port map(D => \RD_USB_ADBUS[5]_net_1\, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_17, E => N_OP_MODE_T_0_sqmuxa, Q
         => \OP_MODE_T[5]_net_1\);
    
    \ELINK_DINA_7[6]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[6]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_17, E => un1_SM_BANK_SEL_12, Q => 
        \ELINK_DINA_7[6]_net_1\);
    
    USB_RXF_B_RNIKSCQ : NOR2B
      port map(A => \USB_RXF_B\, B => \REG_STATE[4]_net_1\, Y => 
        \REG_STATE_ns_i_a4_3_0[4]\);
    
    ELK_N_ACTIVE_RNO : AO1A
      port map(A => N_1697, B => N_1698, C => N_1873, Y => 
        \ELK_N_ACTIVE_RNO\);
    
    \ELINK_ADDRA_0[5]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[5]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_18, E => un1_SM_BANK_SEL_6, Q => 
        \ELINK_ADDRA_0[5]_net_1\);
    
    \WR_USB_ADBUS_RNO_24[3]\ : NOR2B
      port map(A => \ELINK_DOUTA_8[3]\, B => un1_SM_BANK_SEL_38, 
        Y => \ELINK_DOUTA_8_m[3]\);
    
    USB_RXF_B_RNIM7A61 : NOR2B
      port map(A => \USB_RXF_B\, B => N_2526_1, Y => 
        un1_REG_STATE_40_i_a2_2_0);
    
    \SM_BANK_SEL_RNICGCN[7]\ : OR3A
      port map(A => N_462, B => \SM_BANK_SEL[7]_net_1\, C => 
        \SM_BANK_SEL[6]_net_1\, Y => \N_ELINK_RWA_1[14]\);
    
    \WR_XFER_TYPE_RNO[7]\ : AO1A
      port map(A => N_1702, B => N_1728, C => 
        \WR_XFER_TYPE[7]_net_1\, Y => \WR_XFER_TYPE_RNO[7]_net_1\);
    
    \ELINK_ADDRA_0[6]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[6]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_18, E => un1_SM_BANK_SEL_6, Q => 
        \ELINK_ADDRA_0[6]_net_1\);
    
    \ELINK_ADDRA_3[5]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[5]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_1, E => un1_SM_BANK_SEL_4, Q => 
        \ELINK_ADDRA_3[5]_net_1\);
    
    USB_RD_BI_RNO_14 : NOR3B
      port map(A => \REG_STATE_0[2]_net_1\, B => N_1739, C => 
        \USB_RXF_B_0\, Y => N_1865);
    
    \WR_XFER_TYPE_RNI88PP1[2]\ : NOR3B
      port map(A => \WR_XFER_TYPE[7]_net_1\, B => N_1404_6, C => 
        \WR_XFER_TYPE[2]_net_1\, Y => 
        \REG_STATE_ns_i_a2_4_tz_tz_tz_tz[5]\);
    
    \ELINK_ADDRA_15[1]\ : DFN1E0C0
      port map(D => \N_TFC_ADDRA[1]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_6, E => N_199, Q => 
        \ELINK_ADDRA_15[1]_net_1\);
    
    \WR_USB_ADBUS_RNO_5[4]\ : OR3
      port map(A => \ELINK_DOUTA_13_m[4]\, B => 
        \ELINK_DOUTA_12_m[4]\, C => \N_WR_USB_ADBUS_0_iv_12[4]\, 
        Y => \N_WR_USB_ADBUS_0_iv_20[4]\);
    
    \REG_STATE_RNITNN31[2]\ : OR2A
      port map(A => \REG_STATE[2]_net_1\, B => N_1352_1, Y => 
        N_1713);
    
    \ELINKS_STRT_ADDR[1]\ : DFN1E1C0
      port map(D => \ELINKS_STRT_ADDR_T[1]_net_1\, CLK => 
        CLK60MHZ, CLR => P_USB_MASTER_EN_c_17, E => 
        \REG_STATE_d[30]\, Q => \ELINKS_STRT_ADDR[1]_net_1\);
    
    \TFC_STOP_ADDR[0]\ : DFN1E1C0
      port map(D => \TFC_STOP_ADDR_T[0]_net_1\, CLK => CLK60MHZ, 
        CLR => P_USB_MASTER_EN_c_8, E => \REG_STATE_d_0[30]\, Q
         => \TFC_STOP_ADDR[0]_net_1\);
    
    \ELINK_RWA_RNO_0[6]\ : NOR2A
      port map(A => N_622, B => \ELINK_RWA[6]_net_1\, Y => 
        \ELINK_RWA_i_m[6]\);
    
    \ELINK_DINA_9[5]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[5]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_20, E => un1_SM_BANK_SEL_9, Q => 
        \ELINK_DINA_9[5]_net_1\);
    
    \WR_USB_ADBUS_RNO_29[1]\ : NOR3B
      port map(A => N_1730_i, B => \ELINKS_STOP_ADDR[1]_net_1\, C
         => N_1726, Y => \ELINKS_STOP_ADDR_m[1]\);
    
    \ELINK_ADDRA_12[1]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[1]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_2_0, E => un1_SM_BANK_SEL_7, Q => 
        \ELINK_ADDRA_12[1]_net_1\);
    
    \SM_BANK_SEL_RNIJP4B[14]\ : OR2
      port map(A => \SM_BANK_SEL[14]_net_1\, B => 
        \SM_BANK_SEL_0[21]_net_1\, Y => un1_SM_BANK_SEL_15);
    
    \ELINK_RWA_RNO[17]\ : OA1C
      port map(A => N_131, B => \ELINK_RWA[17]_net_1\, C => N_174, 
        Y => \N_ELINK_RWA_0_iv[17]\);
    
    \ELINK_DINA_4[3]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[3]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_13, E => un1_SM_BANK_SEL_8, Q => 
        \ELINK_DINA_4[3]_net_1\);
    
    \ELINK_ADDRA_11[2]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[2]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_2, E => un1_SM_BANK_SEL_16, Q => 
        \ELINK_ADDRA_11[2]_net_1\);
    
    \SM_BANK_SEL_RNI7GJ1[14]\ : OR2
      port map(A => \SM_BANK_SEL[14]_net_1\, B => 
        \SM_BANK_SEL[15]_net_1\, Y => N_622_3);
    
    \REG_STATE_ns_i_i_o2_1_RNO_5[0]\ : NOR3B
      port map(A => \REG_STATE_0[4]_net_1\, B => 
        \REG_STATE_0[5]_net_1\, C => N_2577, Y => 
        \REG_STATE_ns_i_i_a2_1_0[0]\);
    
    \WR_USB_ADBUS_RNO_11[4]\ : OR3
      port map(A => \ELINK_DOUTA_17_m[4]\, B => 
        \ELINK_DOUTA_1_m[4]\, C => \N_WR_USB_ADBUS_0_iv_16[4]\, Y
         => \N_WR_USB_ADBUS_0_iv_22[4]\);
    
    \SM_BANK_SEL_RNIMDLS1[7]\ : NOR3C
      port map(A => N_463, B => N_464, C => 
        \N_ELINK_BLKA_0_iv_0_o2_i_a5_1[11]\, Y => N_393);
    
    \ELINK_BLKA_RNO_0[13]\ : AO1
      port map(A => \N_ELINK_RWA_0_iv_0_o2_i_a5_0[13]\, B => 
        N_503, C => \ELINK_BLKA[13]_net_1\, Y => N_67_tz);
    
    \ELINK_ADDRA_6[1]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[1]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_4, E => un1_SM_BANK_SEL_10, Q => 
        \ELINK_ADDRA_6[1]_net_1\);
    
    USB_OE_BI_RNO : AOI1
      port map(A => N_USB_OE_BI_iv_0_i_a2_0_5, B => 
        N_USB_OE_BI_iv_0_i_a2_0_4, C => N_1871, Y => N_1679);
    
    \REG_STATE_RNIF0PH1[5]\ : NOR2A
      port map(A => \REG_STATE[5]_net_1\, B => N_1765, Y => 
        N_1784);
    
    \ELINK_RWA[18]\ : DFN1E0P0
      port map(D => \N_ELINK_RWA_0_iv[18]\, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_12, E => \SM_BANK_SEL_0[20]_net_1\, 
        Q => \ELINK_RWA[18]_net_1\);
    
    \ELINK_DINA_19[0]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[0]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_0, E => un1_SM_BANK_SEL_11, Q => 
        \ELINK_DINA_19[0]_net_1\);
    
    \REG_STATE_RNIUON31[1]\ : NOR2B
      port map(A => \REG_STATE[1]_net_1\, B => N_2571_1, Y => 
        \REG_STATE_ns_i_a4_3_1_0[1]\);
    
    \ELINK_ADDRA_19[3]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[3]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_13, E => un1_SM_BANK_SEL_11, Q => 
        \ELINK_ADDRA_19[3]_net_1\);
    
    \WR_USB_ADBUS_RNO_1[3]\ : OR3
      port map(A => \N_WR_USB_ADBUS_0_iv_6[3]\, B => 
        \ELINK_DOUTA_14_m[3]\, C => \N_WR_USB_ADBUS_0_iv_18[3]\, 
        Y => \N_WR_USB_ADBUS_0_iv_23[3]\);
    
    \ELINK_RWA_RNO_0[10]\ : OA1B
      port map(A => N_624_15, B => \N_ELINK_RWA_2[10]\, C => 
        \ELINK_RWA[10]_net_1\, Y => \ELINK_RWA_i_m[10]\);
    
    \RD_USB_ADBUS_RNI8S273[4]\ : NOR2
      port map(A => N_1697, B => N_293, Y => N_1882);
    
    \ELINK_RWA_RNO[9]\ : OA1B
      port map(A => N_392, B => \ELINK_RWA[9]_net_1\, C => N_182, 
        Y => \N_ELINK_RWA_0_iv[9]\);
    
    \ELINK_RWA[15]\ : DFN1E0P0
      port map(D => \N_ELINK_RWA_0_iv[15]\, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_12, E => \SM_BANK_SEL_0[20]_net_1\, 
        Q => \ELINK_RWA[15]_net_1\);
    
    \REG_STATE_0_RNIJPPT5[5]\ : OR3
      port map(A => un1_REG_STATE_26_0_1, B => 
        un1_REG_STATE_26_0_0, C => N_1784, Y => un1_REG_STATE_26);
    
    \SM_BANK_SEL_RNO[0]\ : NOR3A
      port map(A => un1_N_ELK_N_ACTIVE_0_sqmuxa_15_0_a2_0_0, B
         => N_1697, C => N_290, Y => N_1834);
    
    \SM_BANK_SEL_RNI6QM12[1]\ : OR3A
      port map(A => N_143, B => \N_ELINK_RWA_1[2]\, C => N_616_16, 
        Y => N_618);
    
    USB_RXF_B_RNICOBDG : OA1
      port map(A => N_285, B => N_1398_i_0_0, C => 
        \REG_STATE_ns_i_a2_0[4]\, Y => \REG_STATE_ns_i_a2_1[4]\);
    
    \TFC_STOP_ADDR[4]\ : DFN1E1C0
      port map(D => \TFC_STOP_ADDR_T[4]_net_1\, CLK => CLK60MHZ, 
        CLR => P_USB_MASTER_EN_c_8, E => \REG_STATE_d_0[30]\, Q
         => \TFC_STOP_ADDR[4]_net_1\);
    
    \SM_BANK_SEL_RNO[12]\ : NOR3B
      port map(A => N_1882, B => N_1359_6, C => N_290, Y => 
        N_1833);
    
    \WR_USB_ADBUS_RNO_27[6]\ : NOR2B
      port map(A => \ELINK_DOUTA_10[6]\, B => un1_SM_BANK_SEL_34, 
        Y => \ELINK_DOUTA_10_m[6]\);
    
    \RD_USB_ADBUS_RNIEVC06[7]\ : OR3
      port map(A => N_1387_i_0_2, B => N_1387_i_0_1, C => N_285, 
        Y => N_1387_i);
    
    \ELINK_RWA_RNO_0[11]\ : NOR2B
      port map(A => \SM_BANK_SEL[8]_net_1\, B => un1_USB_RXF_B_m, 
        Y => N_180);
    
    \WR_USB_ADBUS_RNO_22[1]\ : AO1
      port map(A => \ELINK_DOUTA_15[1]\, B => un1_SM_BANK_SEL_24, 
        C => \ELINK_DOUTA_0_m[1]\, Y => 
        \N_WR_USB_ADBUS_0_iv_8[1]\);
    
    \WR_USB_ADBUS_RNO_11[7]\ : OR3
      port map(A => \ELINK_DOUTA_11_m[7]\, B => 
        \ELINK_DOUTA_10_m[7]\, C => \N_WR_USB_ADBUS_0_iv_16[7]\, 
        Y => \N_WR_USB_ADBUS_0_iv_22[7]\);
    
    \WR_USB_ADBUS_RNO_0[2]\ : OR3
      port map(A => \ELINK_DOUTA_17_m[2]\, B => 
        \ELINK_DOUTA_1_m[2]\, C => \N_WR_USB_ADBUS_0_iv_16[2]\, Y
         => \N_WR_USB_ADBUS_0_iv_22[2]\);
    
    \REG_ADDR_RNO[1]\ : XA1B
      port map(A => \REG_ADDR[1]_net_1\, B => \REG_ADDR[0]_net_1\, 
        C => N_675_0, Y => REG_ADDR_n1);
    
    \RD_USB_ADBUS_RNIV3BJ_0[3]\ : NOR2A
      port map(A => \RD_USB_ADBUS[2]_net_1\, B => 
        \RD_USB_ADBUS[3]_net_1\, Y => N_1359_6);
    
    \ELINK_ADDRA_5[7]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[7]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_3, E => un1_SM_BANK_SEL_15, Q => 
        \ELINK_ADDRA_5[7]_net_1\);
    
    \WR_USB_ADBUS_RNO_23[0]\ : NOR2B
      port map(A => \ELINK_DOUTA_15[0]\, B => un1_SM_BANK_SEL_24, 
        Y => \ELINK_DOUTA_15_m[0]\);
    
    \ELINK_BLKA_RNO_0[2]\ : NOR2B
      port map(A => \SM_BANK_SEL[17]_net_1\, B => X_BLKA_i, Y => 
        X_BLKA_i_m_1);
    
    \REG_ADDR[7]\ : DFN1E1C0
      port map(D => REG_ADDR_n7, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_10, E => REG_ADDRe, Q => 
        \REG_ADDR[7]_net_1\);
    
    \REG_ADDR_RNIJA2T[8]\ : OR3A
      port map(A => \REG_ADDR[8]_net_1\, B => \REG_ADDR[4]_net_1\, 
        C => REG_STATE_tr74_tz_tz_tz_2, Y => 
        REG_STATE_tr74_tz_tz_tz_5);
    
    \N_TFC_ADDRA_0_o2_RNO_6[7]\ : NOR2
      port map(A => N_2497, B => \REG_STATE[1]_net_1\, Y => N_424);
    
    USB_OE_BI_RNO_4 : NOR2A
      port map(A => N_675, B => \USB_RXF_B\, Y => N_1871);
    
    \WR_USB_ADBUS_RNO[5]\ : OR3
      port map(A => \N_WR_USB_ADBUS_0_iv_24[5]\, B => 
        \N_WR_USB_ADBUS_0_iv_23[5]\, C => 
        \N_WR_USB_ADBUS_0_iv_25[5]\, Y => \N_WR_USB_ADBUS[5]\);
    
    \SM_BANK_SEL_RNIUVLB[0]\ : NOR2
      port map(A => \SM_BANK_SEL[0]_net_1\, B => 
        \SM_BANK_SEL[2]_net_1\, Y => N_463);
    
    \WR_USB_ADBUS_RNO_22[6]\ : NOR2B
      port map(A => \ELINK_DOUTA_13[6]\, B => un1_SM_BANK_SEL_29, 
        Y => \ELINK_DOUTA_13_m[6]\);
    
    \SM_BANK_SEL_RNIAUM12[1]\ : OR3A
      port map(A => N_143, B => \N_ELINK_RWA_1[6]\, C => N_616_16, 
        Y => N_622);
    
    \SI_CNT_RNO_0[3]\ : OR2B
      port map(A => N_2607, B => \SI_CNT[2]_net_1\, Y => N_1630);
    
    \ELINK_ADDRA_13[2]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[2]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_3, E => un1_SM_BANK_SEL_2, Q => 
        \ELINK_ADDRA_13[2]_net_1\);
    
    \WR_XFER_TYPE_RNO[5]\ : AO1
      port map(A => N_1763, B => \WR_XFER_TYPE[5]_net_1\, C => 
        N_1829, Y => \WR_XFER_TYPE_RNO[5]_net_1\);
    
    \REG_STATE_RNIOS8OT[0]\ : AO1
      port map(A => N_2587, B => N_1275_tz, C => 
        \REG_STATE_ns_i_1[1]\, Y => \REG_STATE_ns_i_2[1]\);
    
    \ELINK_DINA_13[1]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[1]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_14, E => un1_SM_BANK_SEL_2, Q => 
        \ELINK_DINA_13[1]_net_1\);
    
    \WR_USB_ADBUS_RNO_19[7]\ : AO1
      port map(A => \CHKSUM[7]_net_1\, B => un1_REG_STATE_4, C
         => \N_WR_USB_ADBUS_0_iv_1[7]\, Y => 
        \N_WR_USB_ADBUS_0_iv_4[7]\);
    
    \REG_STATE_0_RNIR72S[0]\ : XNOR2
      port map(A => \REG_STATE_0[1]_net_1\, B => 
        \REG_STATE_0[0]_net_1\, Y => N_2462);
    
    \ELINK_BLKA[17]\ : DFN1E0P0
      port map(D => \N_ELINK_BLKA_0_iv[17]\, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_20, E => \SM_BANK_SEL[20]_net_1\, Q
         => \ELINK_BLKA[17]_net_1\);
    
    USB_RXF_B : DFN1P0
      port map(D => P_USB_RXF_B_c, CLK => CLK60MHZ, PRE => 
        P_USB_MASTER_EN_c, Q => \USB_RXF_B\);
    
    \WR_USB_ADBUS_RNO_9[4]\ : AO1
      port map(A => \ELINK_DOUTA_0[4]\, B => un1_SM_BANK_SEL_31, 
        C => \ELINK_DOUTA_16_m[4]\, Y => 
        \N_WR_USB_ADBUS_0_iv_14[4]\);
    
    \ELINKS_STRT_ADDR[2]\ : DFN1E1C0
      port map(D => \ELINKS_STRT_ADDR_T[2]_net_1\, CLK => 
        CLK60MHZ, CLR => P_USB_MASTER_EN_c_17, E => 
        \REG_STATE_d[30]\, Q => \ELINKS_STRT_ADDR[2]_net_1\);
    
    \ELINK_ADDRA_9[2]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[2]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_10, E => un1_SM_BANK_SEL_9, Q => 
        \ELINK_ADDRA_9[2]_net_1\);
    
    \WR_USB_ADBUS_RNO_24[7]\ : NOR2B
      port map(A => \ELINK_DOUTA_8[7]\, B => un1_SM_BANK_SEL_38, 
        Y => \ELINK_DOUTA_8_m[7]\);
    
    \RD_USB_ADBUS_RNITB1Q1[5]\ : NOR3B
      port map(A => N_1352_4, B => N_1903, C => 
        \RD_USB_ADBUS[5]_net_1\, Y => 
        un1_N_ELK_N_ACTIVE_2_sqmuxa_0_a2_0_0);
    
    \ELINK_BLKA[2]\ : DFN1E0P0
      port map(D => \N_ELINK_BLKA_0_iv[2]\, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_19, E => \SM_BANK_SEL[20]_net_1\, Q
         => \ELINK_BLKA[2]_net_1\);
    
    \ELINK_ADDRA_4[6]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[6]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_2_0, E => un1_SM_BANK_SEL_8, Q => 
        \ELINK_ADDRA_4[6]_net_1\);
    
    \REG_STATE_0_RNIJDMT1[5]\ : AO1D
      port map(A => N_312, B => \REG_STATE_0[5]_net_1\, C => 
        N_1877_1, Y => N_2467);
    
    \ELINK_DINA_11[7]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[7]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_11, E => un1_SM_BANK_SEL_16, Q => 
        \ELINK_DINA_11[7]_net_1\);
    
    \SM_BANK_SEL_RNII31C2[8]\ : NOR3A
      port map(A => \SM_BANK_SEL[8]_net_1\, B => N_312_0, C => 
        N_1566_i_i_0, Y => un1_SM_BANK_SEL_26);
    
    \REG_ADDR_RNI6T1T[3]\ : NOR2B
      port map(A => N_474, B => \REG_ADDR[3]_net_1\, Y => 
        REG_ADDR_c3);
    
    ELK_N_ACTIVE_RNI3GEF9 : AOI1
      port map(A => N_480, B => \ELK_N_ACTIVE\, C => N_1374, Y
         => \REG_STATE_ns_i_a2_0[3]\);
    
    \REG_ADDR_RNO[0]\ : NOR2
      port map(A => \REG_ADDR[0]_net_1\, B => N_675, Y => N_2624);
    
    \ELINK_RWA_RNO_0[12]\ : OA1B
      port map(A => N_624_15, B => \N_ELINK_RWA_1[12]\, C => 
        \ELINK_RWA[12]_net_1\, Y => \ELINK_RWA_i_m[12]\);
    
    \ELINKS_STRT_ADDR_T[7]\ : DFN1E1C0
      port map(D => \RD_USB_ADBUS[7]_net_1\, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_21, E => 
        N_ELINKS_STRT_ADDR_T_0_sqmuxa, Q => 
        \ELINKS_STRT_ADDR_T[7]_net_1\);
    
    \WR_USB_ADBUS_RNO_25[0]\ : NOR2B
      port map(A => \ELINK_DOUTA_1[0]\, B => un1_SM_BANK_SEL_36, 
        Y => \ELINK_DOUTA_1_m[0]\);
    
    \WR_USB_ADBUS_RNO_16[0]\ : AO1
      port map(A => \ELINK_DOUTA_14[0]\, B => un1_SM_BANK_SEL_23, 
        C => \ELINK_DOUTA_19_m[0]\, Y => 
        \N_WR_USB_ADBUS_0_iv_12[0]\);
    
    \RD_USB_ADBUS_RNIMAJO2[6]\ : NOR2A
      port map(A => N_1729, B => N_1694, Y => N_1911);
    
    \ELINK_RWA_RNO[19]\ : OA1C
      port map(A => N_130, B => \ELINK_RWA[19]_net_1\, C => N_170, 
        Y => \N_ELINK_RWA_0_iv[19]\);
    
    \ELINK_ADDRA_1[6]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[6]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_20, E => un1_SM_BANK_SEL_19, Q => 
        \ELINK_ADDRA_1[6]_net_1\);
    
    \WR_USB_ADBUS_RNO_26[5]\ : NOR2B
      port map(A => \ELINK_DOUTA_11[5]\, B => un1_SM_BANK_SEL_26, 
        Y => \ELINK_DOUTA_11_m[5]\);
    
    \RD_USB_ADBUS_RNIRVAJ[0]\ : XOR2
      port map(A => \RD_USB_ADBUS[1]_net_1\, B => 
        \RD_USB_ADBUS[0]_net_1\, Y => N_310);
    
    \ELINK_BLKA_RNO_0[16]\ : AOI1
      port map(A => \N_ELINK_RWA_i_a2_0_a5_0[16]\, B => N_503, C
         => \ELINK_BLKA[16]_net_1\, Y => \ELINK_BLKA_i_m[16]\);
    
    \TFC_STRT_ADDR_T[7]\ : DFN1E1C0
      port map(D => \RD_USB_ADBUS[7]_net_1\, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_5, E => N_TFC_STRT_ADDR_T_0_sqmuxa, 
        Q => \TFC_STRT_ADDR_T[7]_net_1\);
    
    TFC_RWA : DFN1E0P0
      port map(D => N_206, CLK => CLK60MHZ, PRE => 
        P_USB_MASTER_EN_c_3, E => N_142, Q => \TFC_RWA\);
    
    USB_RXF_B_0_RNIU2AB1 : MX2
      port map(A => \REG_STATE_0[2]_net_1\, B => \USB_RXF_B_0\, S
         => \REG_STATE_0[1]_net_1\, Y => N_2498);
    
    \REG_STATE_RNIUFQN[0]\ : OR2B
      port map(A => \REG_STATE[0]_net_1\, B => 
        \REG_STATE[2]_net_1\, Y => N_2497);
    
    \ELINK_BLKA[10]\ : DFN1E0P0
      port map(D => \N_ELINK_BLKA_0_iv[10]\, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_20, E => \SM_BANK_SEL[20]_net_1\, Q
         => \ELINK_BLKA[10]_net_1\);
    
    \ELINK_ADDRA_2[1]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[1]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_21, E => un1_SM_BANK_SEL_5, Q => 
        \ELINK_ADDRA_2[1]_net_1\);
    
    \WR_USB_ADBUS_RNO_15[6]\ : NOR2B
      port map(A => \ELINK_DOUTA_19[6]\, B => un1_SM_BANK_SEL_41, 
        Y => \ELINK_DOUTA_19_m[6]\);
    
    TFC_BLKA_RNO : OR2A
      port map(A => X_BLKA_i, B => \SM_BANK_SEL[21]_net_1\, Y => 
        N_TFC_BLKA);
    
    \REG_STATE_0_RNIGFUP[3]\ : NOR2
      port map(A => \REG_STATE_0[3]_net_1\, B => 
        \REG_STATE[2]_net_1\, Y => N_1352_2);
    
    \SM_BANK_SEL_RNO[13]\ : NOR3C
      port map(A => N_1882, B => N_1359_6, C => N_1352_4, Y => 
        N_1844);
    
    USB_OE_BI_RNO_3 : NOR3A
      port map(A => N_USB_OE_BI_iv_0_i_a2_0_1, B => N_1751, C => 
        N_293, Y => N_USB_OE_BI_iv_0_i_a2_0_4);
    
    \WR_USB_ADBUS_RNO_30[7]\ : AO1A
      port map(A => N_1501, B => \TFC_STOP_ADDR[7]_net_1\, C => 
        \OP_MODE_m[7]\, Y => \N_WR_USB_ADBUS_0_iv_0[7]\);
    
    \REG_STATE_RNIP2V25[4]\ : AO1
      port map(A => N_2613, B => N_350, C => N_675_0, Y => N_678);
    
    un1_REG_STATE_4_0_a2_0 : NOR2A
      port map(A => N_1782_1, B => N_1726, Y => N_1782);
    
    \SM_BANK_SEL[3]\ : DFN1E1C0
      port map(D => N_1849, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_7, E => un1_REG_STATE_30, Q => 
        \SM_BANK_SEL[3]_net_1\);
    
    \SM_BANK_SEL[10]\ : DFN1E1C0
      port map(D => N_1839, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_1_0, E => un1_REG_STATE_30, Q => 
        \SM_BANK_SEL[10]_net_1\);
    
    \WR_USB_ADBUS_RNO_32[3]\ : NOR2B
      port map(A => \WR_XFER_TYPE[3]_net_1\, B => N_398, Y => 
        \WR_XFER_TYPE_m[3]\);
    
    \ELINK_ADDRA_18[5]\ : DFN1E0C0
      port map(D => \N_TFC_ADDRA[5]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_12, E => N_198, Q => 
        \ELINK_ADDRA_18[5]_net_1\);
    
    \ELINK_DINA_1[5]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[5]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_7, E => un1_SM_BANK_SEL_19, Q => 
        \ELINK_DINA_1[5]_net_1\);
    
    \ELINK_DINA_19[4]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[4]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_1, E => un1_SM_BANK_SEL_11, Q => 
        \ELINK_DINA_19[4]_net_1\);
    
    \SM_BANK_SEL_RNI9IJ1[16]\ : OR2
      port map(A => \SM_BANK_SEL[16]_net_1\, B => 
        \SM_BANK_SEL[15]_net_1\, Y => N_616_2);
    
    USB_TXE_B_RNIB8SV6 : OR3
      port map(A => N_1704, B => N_396, C => N_675_0, Y => 
        REG_ADDRe);
    
    \REG_STATE_RNIGERD2[4]\ : NOR2B
      port map(A => N_1917, B => \REG_STATE[4]_net_1\, Y => 
        N_1860);
    
    \ELINK_BLKA[19]\ : DFN1E0P0
      port map(D => \N_ELINK_BLKA_0_iv[19]\, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_20, E => \SM_BANK_SEL[20]_net_1\, Q
         => \ELINK_BLKA[19]_net_1\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    USB_TXE_B_RNIJRFM1 : NOR3B
      port map(A => N_2600, B => N_2497, C => \USB_TXE_B\, Y => 
        N_396);
    
    \WR_USB_ADBUS_RNO_32[0]\ : NOR3B
      port map(A => N_1352_1, B => \OP_MODE[0]_net_1\, C => 
        REG_STATE_s20_i_0, Y => \OP_MODE_m[0]\);
    
    \SM_BANK_SEL_RNI19VN[1]\ : OR2A
      port map(A => N_143, B => N_624_15, Y => \N_ELINK_RWA_0[8]\);
    
    \WR_USB_ADBUS_RNO_27[1]\ : AO1
      port map(A => \ELINK_DOUTA_12[1]\, B => un1_SM_BANK_SEL_33, 
        C => \ELINK_DOUTA_13_m[1]\, Y => 
        \N_WR_USB_ADBUS_0_iv_16[1]\);
    
    \REG_STATE_RNIPNS13[5]\ : AO1A
      port map(A => N_252, B => N_446, C => N_427, Y => N_254);
    
    \ELINK_DINA_15[6]\ : DFN1E0C0
      port map(D => \N_TFC_DINA[6]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_16, E => N_199, Q => 
        \ELINK_DINA_15[6]_net_1\);
    
    U0_PATT_TFC_BLK : DPRT_512X9_SRAM
      port map(TFC_RX_SER_WORD(7) => TFC_RX_SER_WORD(7), 
        TFC_RX_SER_WORD(6) => TFC_RX_SER_WORD(6), 
        TFC_RX_SER_WORD(5) => TFC_RX_SER_WORD(5), 
        TFC_RX_SER_WORD(4) => TFC_RX_SER_WORD(4), 
        TFC_RX_SER_WORD(3) => TFC_RX_SER_WORD(3), 
        TFC_RX_SER_WORD(2) => TFC_RX_SER_WORD(2), 
        TFC_RX_SER_WORD(1) => TFC_RX_SER_WORD(1), 
        TFC_RX_SER_WORD(0) => TFC_RX_SER_WORD(0), TFC_DINA(7) => 
        \TFC_DINA[7]_net_1\, TFC_DINA(6) => \TFC_DINA[6]_net_1\, 
        TFC_DINA(5) => \TFC_DINA[5]_net_1\, TFC_DINA(4) => 
        \TFC_DINA[4]_net_1\, TFC_DINA(3) => \TFC_DINA[3]_net_1\, 
        TFC_DINA(2) => \TFC_DINA[2]_net_1\, TFC_DINA(1) => 
        \TFC_DINA[1]_net_1\, TFC_DINA(0) => \TFC_DINA[0]_net_1\, 
        TFC_ADDRB(7) => TFC_ADDRB(7), TFC_ADDRB(6) => 
        TFC_ADDRB(6), TFC_ADDRB(5) => TFC_ADDRB(5), TFC_ADDRB(4)
         => TFC_ADDRB(4), TFC_ADDRB(3) => TFC_ADDRB(3), 
        TFC_ADDRB(2) => TFC_ADDRB(2), TFC_ADDRB(1) => 
        TFC_ADDRB(1), TFC_ADDRB(0) => TFC_ADDRB(0), TFC_ADDRA(7)
         => \TFC_ADDRA[7]_net_1\, TFC_ADDRA(6) => 
        \TFC_ADDRA[6]_net_1\, TFC_ADDRA(5) => 
        \TFC_ADDRA[5]_net_1\, TFC_ADDRA(4) => 
        \TFC_ADDRA[4]_net_1\, TFC_ADDRA(3) => 
        \TFC_ADDRA[3]_net_1\, TFC_ADDRA(2) => 
        \TFC_ADDRA[2]_net_1\, TFC_ADDRA(1) => 
        \TFC_ADDRA[1]_net_1\, TFC_ADDRA(0) => 
        \TFC_ADDRA[0]_net_1\, PATT_TFC_DAT(7) => PATT_TFC_DAT(7), 
        PATT_TFC_DAT(6) => PATT_TFC_DAT(6), PATT_TFC_DAT(5) => 
        PATT_TFC_DAT(5), PATT_TFC_DAT(4) => PATT_TFC_DAT(4), 
        PATT_TFC_DAT(3) => PATT_TFC_DAT(3), PATT_TFC_DAT(2) => 
        PATT_TFC_DAT(2), PATT_TFC_DAT(1) => PATT_TFC_DAT(1), 
        PATT_TFC_DAT(0) => PATT_TFC_DAT(0), TFC_DOUTA(7) => 
        \TFC_DOUTA[7]\, TFC_DOUTA(6) => \TFC_DOUTA[6]\, 
        TFC_DOUTA(5) => \TFC_DOUTA[5]\, TFC_DOUTA(4) => 
        \TFC_DOUTA[4]\, TFC_DOUTA(3) => \TFC_DOUTA[3]\, 
        TFC_DOUTA(2) => \TFC_DOUTA[2]\, TFC_DOUTA(1) => 
        \TFC_DOUTA[1]\, TFC_DOUTA(0) => \TFC_DOUTA[0]\, TFC_RWB
         => TFC_RWB, TFC_RWA => \TFC_RWA\, P_USB_MASTER_EN_c_0
         => P_USB_MASTER_EN_c_0, CLK_40M_GL => CLK_40M_GL, 
        CLK60MHZ => CLK60MHZ, TFC_RAM_BLKB_EN => TFC_RAM_BLKB_EN, 
        TFC_BLKA => \TFC_BLKA\);
    
    \REG_STATE_RNIUON31_0[1]\ : NOR2A
      port map(A => \REG_STATE[1]_net_1\, B => N_257, Y => N_470);
    
    \RD_XFER_TYPE[1]\ : DFN1C0
      port map(D => \RD_XFER_TYPE_RNO[1]_net_1\, CLK => CLK60MHZ, 
        CLR => P_USB_MASTER_EN_c, Q => \RD_XFER_TYPE[1]_net_1\);
    
    \REG_STATE_RNIUFQN_0[0]\ : NOR2
      port map(A => \REG_STATE[0]_net_1\, B => 
        \REG_STATE[2]_net_1\, Y => N_1710_i_0);
    
    \ELINK_BLKA_RNO[13]\ : AOI1B
      port map(A => \SM_BANK_SEL[6]_net_1\, B => X_BLKA_i, C => 
        N_67_tz, Y => N_67);
    
    \ELINK_BLKA_RNO[7]\ : AOI1
      port map(A => \SM_BANK_SEL[12]_net_1\, B => X_BLKA_i, C => 
        \ELINK_BLKA_i_m[7]\, Y => \N_ELINK_BLKA_0_iv[7]\);
    
    \SM_BANK_SEL_RNI7P63[13]\ : OR3
      port map(A => \SM_BANK_SEL[15]_net_1\, B => 
        \SM_BANK_SEL[13]_net_1\, C => N_616_4, Y => 
        \N_ELINK_RWA_1[5]\);
    
    \SM_BANK_SEL_RNIUIV62[13]\ : NOR3A
      port map(A => \SM_BANK_SEL[13]_net_1\, B => N_312_0, C => 
        N_1566_i_i_0, Y => un1_SM_BANK_SEL_30);
    
    \RD_XFER_TYPE_RNI9C6HP[0]\ : OR3
      port map(A => N_358, B => N_357, C => 
        \REG_STATE_ns_i_i_0[0]\, Y => \REG_STATE_ns_i_i_2[0]\);
    
    \RD_USB_ADBUS_RNIJ9NS7[6]\ : AOI1B
      port map(A => un1_REG_STATE_35_i_a2_0, B => N_1772, C => 
        N_1737, Y => N_1671);
    
    \SM_BANK_SEL_RNIHNL6[2]\ : NOR2
      port map(A => \SM_BANK_SEL[2]_net_1\, B => 
        \SM_BANK_SEL[21]_net_1\, Y => N_197);
    
    \REG_STATE_ns_i_i_o2_1_RNO_2[0]\ : NOR3B
      port map(A => \REG_STATE_0[4]_net_1\, B => 
        \REG_STATE_ns_i_i_a2_9_0[0]\, C => N_2577, Y => N_438);
    
    \ELINK_ADDRA_13[3]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[3]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_3, E => un1_SM_BANK_SEL_2, Q => 
        \ELINK_ADDRA_13[3]_net_1\);
    
    \ELINK_DINA_8[2]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[2]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_18, E => un1_SM_BANK_SEL_21, Q => 
        \ELINK_DINA_8[2]_net_1\);
    
    \ELINK_DINA_17[0]\ : DFN1E0C0
      port map(D => \N_TFC_DINA[0]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_19, E => N_197, Q => 
        \ELINK_DINA_17[0]_net_1\);
    
    \WR_USB_ADBUS_RNO_29[4]\ : OR3
      port map(A => \N_WR_USB_ADBUS_0_iv_0[4]_net_1\, B => 
        \OP_MODE_m[4]\, C => \ELINKS_STRT_ADDR_m[4]\, Y => 
        \N_WR_USB_ADBUS_0_iv_2[4]\);
    
    \ELINK_BLKA[5]\ : DFN1E0P0
      port map(D => \N_ELINK_BLKA_0_iv[5]\, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_19, E => \SM_BANK_SEL[20]_net_1\, Q
         => \ELINK_BLKA[5]_net_1\);
    
    \WR_USB_ADBUS_RNO_8[0]\ : OR3
      port map(A => \N_WR_USB_ADBUS_0_iv_5[0]\, B => 
        \N_WR_USB_ADBUS_0_iv_4[0]\, C => \ELINK_DOUTA_3_m[0]\, Y
         => \N_WR_USB_ADBUS_0_iv_17[0]\);
    
    \REG_STATE_ns_i_i_o2_1_RNO_3[0]\ : NOR3A
      port map(A => \REG_STATE_0[2]_net_1\, B => 
        \REG_STATE_0[0]_net_1\, C => \USB_TXE_B\, Y => N_440);
    
    \WR_USB_ADBUS_RNO_0[3]\ : OR3
      port map(A => \N_WR_USB_ADBUS_0_iv_10[3]\, B => 
        \N_WR_USB_ADBUS_0_iv_9[3]\, C => 
        \N_WR_USB_ADBUS_0_iv_20[3]\, Y => 
        \N_WR_USB_ADBUS_0_iv_24[3]\);
    
    \ELINK_DINA_10[5]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[5]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_9, E => un1_SM_BANK_SEL_20, Q => 
        \ELINK_DINA_10[5]_net_1\);
    
    \WR_USB_ADBUS_RNO_8[6]\ : OR3
      port map(A => \N_WR_USB_ADBUS_0_iv_4[6]\, B => 
        \N_WR_USB_ADBUS_0_iv_3[6]\, C => \ELINK_DOUTA_3_m[6]\, Y
         => \N_WR_USB_ADBUS_0_iv_16[6]\);
    
    USB_TXE_B_RNIL2OI_0 : OR2A
      port map(A => \REG_STATE[4]_net_1\, B => \USB_TXE_B\, Y => 
        N_1749);
    
    U110_PATT_ELINK_BLK : DPRT_512X9_SRAM_10
      port map(ELINK_RWA_0 => \ELINK_RWA[10]_net_1\, 
        ELK_RX_SER_WORD_10(7) => ELK_RX_SER_WORD_10(7), 
        ELK_RX_SER_WORD_10(6) => ELK_RX_SER_WORD_10(6), 
        ELK_RX_SER_WORD_10(5) => ELK_RX_SER_WORD_10(5), 
        ELK_RX_SER_WORD_10(4) => ELK_RX_SER_WORD_10(4), 
        ELK_RX_SER_WORD_10(3) => ELK_RX_SER_WORD_10(3), 
        ELK_RX_SER_WORD_10(2) => ELK_RX_SER_WORD_10(2), 
        ELK_RX_SER_WORD_10(1) => ELK_RX_SER_WORD_10(1), 
        ELK_RX_SER_WORD_10(0) => ELK_RX_SER_WORD_10(0), 
        ELINK_DINA_10(7) => \ELINK_DINA_10[7]_net_1\, 
        ELINK_DINA_10(6) => \ELINK_DINA_10[6]_net_1\, 
        ELINK_DINA_10(5) => \ELINK_DINA_10[5]_net_1\, 
        ELINK_DINA_10(4) => \ELINK_DINA_10[4]_net_1\, 
        ELINK_DINA_10(3) => \ELINK_DINA_10[3]_net_1\, 
        ELINK_DINA_10(2) => \ELINK_DINA_10[2]_net_1\, 
        ELINK_DINA_10(1) => \ELINK_DINA_10[1]_net_1\, 
        ELINK_DINA_10(0) => \ELINK_DINA_10[0]_net_1\, 
        ELINK_BLKA_0 => \ELINK_BLKA[10]_net_1\, ELKS_ADDRB_0_d0
         => ELKS_ADDRB(0), ELKS_ADDRB_1 => ELKS_ADDRB(1), 
        ELKS_ADDRB_3 => ELKS_ADDRB(3), ELKS_ADDRB_5 => 
        ELKS_ADDRB(5), ELKS_ADDRB_7 => ELKS_ADDRB(7), 
        ELKS_ADDRB_0_0 => ELKS_ADDRB_0_0, ELKS_ADDRB_0_2 => 
        ELKS_ADDRB_0_2, ELKS_ADDRB_0_4 => ELKS_ADDRB_0_4, 
        ELINK_ADDRA_10(7) => \ELINK_ADDRA_10[7]_net_1\, 
        ELINK_ADDRA_10(6) => \ELINK_ADDRA_10[6]_net_1\, 
        ELINK_ADDRA_10(5) => \ELINK_ADDRA_10[5]_net_1\, 
        ELINK_ADDRA_10(4) => \ELINK_ADDRA_10[4]_net_1\, 
        ELINK_ADDRA_10(3) => \ELINK_ADDRA_10[3]_net_1\, 
        ELINK_ADDRA_10(2) => \ELINK_ADDRA_10[2]_net_1\, 
        ELINK_ADDRA_10(1) => \ELINK_ADDRA_10[1]_net_1\, 
        ELINK_ADDRA_10(0) => \ELINK_ADDRA_10[0]_net_1\, 
        PATT_ELK_DAT_10(7) => PATT_ELK_DAT_10(7), 
        PATT_ELK_DAT_10(6) => PATT_ELK_DAT_10(6), 
        PATT_ELK_DAT_10(5) => PATT_ELK_DAT_10(5), 
        PATT_ELK_DAT_10(4) => PATT_ELK_DAT_10(4), 
        PATT_ELK_DAT_10(3) => PATT_ELK_DAT_10(3), 
        PATT_ELK_DAT_10(2) => PATT_ELK_DAT_10(2), 
        PATT_ELK_DAT_10(1) => PATT_ELK_DAT_10(1), 
        PATT_ELK_DAT_10(0) => PATT_ELK_DAT_10(0), 
        ELINK_DOUTA_10(7) => \ELINK_DOUTA_10[7]\, 
        ELINK_DOUTA_10(6) => \ELINK_DOUTA_10[6]\, 
        ELINK_DOUTA_10(5) => \ELINK_DOUTA_10[5]\, 
        ELINK_DOUTA_10(4) => \ELINK_DOUTA_10[4]\, 
        ELINK_DOUTA_10(3) => \ELINK_DOUTA_10[3]\, 
        ELINK_DOUTA_10(2) => \ELINK_DOUTA_10[2]\, 
        ELINK_DOUTA_10(1) => \ELINK_DOUTA_10[1]\, 
        ELINK_DOUTA_10(0) => \ELINK_DOUTA_10[0]\, ELKS_RWB => 
        ELKS_RWB, P_USB_MASTER_EN_c_0 => P_USB_MASTER_EN_c_0, 
        CLK_40M_GL => CLK_40M_GL, CLK60MHZ => CLK60MHZ, 
        ELKS_RAM_BLKB_EN => ELKS_RAM_BLKB_EN);
    
    \ELINK_ADDRA_1[1]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[1]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_20, E => un1_SM_BANK_SEL_19, Q => 
        \ELINK_ADDRA_1[1]_net_1\);
    
    \ELINK_ADDRA_12[7]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[7]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_3, E => un1_SM_BANK_SEL_7, Q => 
        \ELINK_ADDRA_12[7]_net_1\);
    
    \SI_CNT_RNO[1]\ : XA1B
      port map(A => \SI_CNT[1]_net_1\, B => \SI_CNT[0]_net_1\, C
         => N_678, Y => SI_CNT_n1);
    
    \USB_WR_BI\ : DFN1E1P0
      port map(D => un1_REG_STATE_26, CLK => CLK60MHZ, PRE => 
        P_USB_MASTER_EN_c_19, E => un1_REG_STATE_28, Q => 
        USB_WR_BI);
    
    \TFC_STOP_ADDR_T[1]\ : DFN1E1C0
      port map(D => \RD_USB_ADBUS[1]_net_1\, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_15, E => N_TFC_STOP_ADDR_T_0_sqmuxa, 
        Q => \TFC_STOP_ADDR_T[1]_net_1\);
    
    \SM_BANK_SEL_RNITHV62[12]\ : NOR3A
      port map(A => \SM_BANK_SEL[12]_net_1\, B => N_312_0, C => 
        N_1566_i_i_0, Y => un1_SM_BANK_SEL_37);
    
    \REG_STATE_0_RNIVAFF3[2]\ : OR2
      port map(A => N_454, B => N_1784, Y => un1_REG_STATE_18);
    
    USB_RD_BI_RNO_5 : NOR2B
      port map(A => \USB_RXF_B\, B => \REG_STATE[2]_net_1\, Y => 
        un1_REG_STATE_40_i_a2_0_0);
    
    \ELINK_DINA_19[7]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[7]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_1, E => un1_SM_BANK_SEL_11, Q => 
        \ELINK_DINA_19[7]_net_1\);
    
    \WR_USB_ADBUS_RNO_4[4]\ : AO1
      port map(A => \ELINK_DOUTA_8[4]\, B => un1_SM_BANK_SEL_38, 
        C => \ELINK_DOUTA_9_m[4]\, Y => 
        \N_WR_USB_ADBUS_0_iv_9[4]\);
    
    \REG_STATE_RNI5NQN_0[5]\ : NOR2B
      port map(A => \REG_STATE[5]_net_1\, B => 
        \REG_STATE[4]_net_1\, Y => N_1421_3);
    
    \WR_XFER_TYPE_RNIUT9V[5]\ : OAI1
      port map(A => \WR_XFER_TYPE[1]_net_1\, B => 
        \WR_XFER_TYPE[5]_net_1\, C => \ELK_N_ACTIVE\, Y => 
        \REG_STATE_ns_i_a2_0_0_0[5]\);
    
    \REG_STATE_RNIVPG2K2[2]\ : OR3A
      port map(A => N_513, B => \RD_USB_ADBUS_RNIP4GES[4]_net_1\, 
        C => \REG_STATE_ns_i_i_0[2]\, Y => 
        \REG_STATE_RNIVPG2K2[2]_net_1\);
    
    \WR_USB_ADBUS_RNO_31[1]\ : NOR2A
      port map(A => \TFC_STOP_ADDR[1]_net_1\, B => N_1501, Y => 
        \TFC_STOP_ADDR_m[1]\);
    
    \WR_USB_ADBUS_RNO_33[4]\ : NOR2A
      port map(A => \ELINKS_STRT_ADDR[4]_net_1\, B => N_1499, Y
         => \ELINKS_STRT_ADDR_m[4]\);
    
    \REG_ADDR[0]\ : DFN1E1C0
      port map(D => N_2624, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_10, E => REG_ADDRe, Q => 
        \REG_ADDR[0]_net_1\);
    
    \ELINK_DINA_8[1]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[1]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_18, E => un1_SM_BANK_SEL_21, Q => 
        \ELINK_DINA_8[1]_net_1\);
    
    \WR_USB_ADBUS_RNO_6[7]\ : OR3
      port map(A => \N_WR_USB_ADBUS_0_iv_3[7]\, B => 
        \N_WR_USB_ADBUS_0_iv_2[7]\, C => 
        \N_WR_USB_ADBUS_0_iv_4[7]\, Y => 
        \N_WR_USB_ADBUS_0_iv_6[7]\);
    
    U108_PATT_ELINK_BLK : DPRT_512X9_SRAM_8
      port map(ELINK_RWA_0 => \ELINK_RWA[8]_net_1\, 
        ELK_RX_SER_WORD_8(7) => ELK_RX_SER_WORD_8(7), 
        ELK_RX_SER_WORD_8(6) => ELK_RX_SER_WORD_8(6), 
        ELK_RX_SER_WORD_8(5) => ELK_RX_SER_WORD_8(5), 
        ELK_RX_SER_WORD_8(4) => ELK_RX_SER_WORD_8(4), 
        ELK_RX_SER_WORD_8(3) => ELK_RX_SER_WORD_8(3), 
        ELK_RX_SER_WORD_8(2) => ELK_RX_SER_WORD_8(2), 
        ELK_RX_SER_WORD_8(1) => ELK_RX_SER_WORD_8(1), 
        ELK_RX_SER_WORD_8(0) => ELK_RX_SER_WORD_8(0), 
        ELINK_DINA_8(7) => \ELINK_DINA_8[7]_net_1\, 
        ELINK_DINA_8(6) => \ELINK_DINA_8[6]_net_1\, 
        ELINK_DINA_8(5) => \ELINK_DINA_8[5]_net_1\, 
        ELINK_DINA_8(4) => \ELINK_DINA_8[4]_net_1\, 
        ELINK_DINA_8(3) => \ELINK_DINA_8[3]_net_1\, 
        ELINK_DINA_8(2) => \ELINK_DINA_8[2]_net_1\, 
        ELINK_DINA_8(1) => \ELINK_DINA_8[1]_net_1\, 
        ELINK_DINA_8(0) => \ELINK_DINA_8[0]_net_1\, ELINK_BLKA_0
         => \ELINK_BLKA[8]_net_1\, ELKS_ADDRB_0_d0 => 
        ELKS_ADDRB(0), ELKS_ADDRB_1 => ELKS_ADDRB(1), 
        ELKS_ADDRB_3 => ELKS_ADDRB(3), ELKS_ADDRB_5 => 
        ELKS_ADDRB(5), ELKS_ADDRB_7 => ELKS_ADDRB(7), 
        ELKS_ADDRB_0_0 => ELKS_ADDRB_0_0, ELKS_ADDRB_0_2 => 
        ELKS_ADDRB_0_2, ELKS_ADDRB_0_4 => ELKS_ADDRB_0_4, 
        ELINK_ADDRA_8(7) => \ELINK_ADDRA_8[7]_net_1\, 
        ELINK_ADDRA_8(6) => \ELINK_ADDRA_8[6]_net_1\, 
        ELINK_ADDRA_8(5) => \ELINK_ADDRA_8[5]_net_1\, 
        ELINK_ADDRA_8(4) => \ELINK_ADDRA_8[4]_net_1\, 
        ELINK_ADDRA_8(3) => \ELINK_ADDRA_8[3]_net_1\, 
        ELINK_ADDRA_8(2) => \ELINK_ADDRA_8[2]_net_1\, 
        ELINK_ADDRA_8(1) => \ELINK_ADDRA_8[1]_net_1\, 
        ELINK_ADDRA_8(0) => \ELINK_ADDRA_8[0]_net_1\, 
        PATT_ELK_DAT_8(7) => PATT_ELK_DAT_8(7), PATT_ELK_DAT_8(6)
         => PATT_ELK_DAT_8(6), PATT_ELK_DAT_8(5) => 
        PATT_ELK_DAT_8(5), PATT_ELK_DAT_8(4) => PATT_ELK_DAT_8(4), 
        PATT_ELK_DAT_8(3) => PATT_ELK_DAT_8(3), PATT_ELK_DAT_8(2)
         => PATT_ELK_DAT_8(2), PATT_ELK_DAT_8(1) => 
        PATT_ELK_DAT_8(1), PATT_ELK_DAT_8(0) => PATT_ELK_DAT_8(0), 
        ELINK_DOUTA_8(7) => \ELINK_DOUTA_8[7]\, ELINK_DOUTA_8(6)
         => \ELINK_DOUTA_8[6]\, ELINK_DOUTA_8(5) => 
        \ELINK_DOUTA_8[5]\, ELINK_DOUTA_8(4) => 
        \ELINK_DOUTA_8[4]\, ELINK_DOUTA_8(3) => 
        \ELINK_DOUTA_8[3]\, ELINK_DOUTA_8(2) => 
        \ELINK_DOUTA_8[2]\, ELINK_DOUTA_8(1) => 
        \ELINK_DOUTA_8[1]\, ELINK_DOUTA_8(0) => 
        \ELINK_DOUTA_8[0]\, ELKS_RWB => ELKS_RWB, 
        P_USB_MASTER_EN_c_0 => P_USB_MASTER_EN_c_0, CLK_40M_GL
         => CLK_40M_GL, CLK60MHZ => CLK60MHZ, ELKS_RAM_BLKB_EN
         => ELKS_RAM_BLKB_EN);
    
    \WR_USB_ADBUS_RNO_10[1]\ : AO1
      port map(A => \ELINK_DOUTA_6[1]\, B => un1_SM_BANK_SEL_30, 
        C => \ELINK_DOUTA_8_m[1]\, Y => 
        \N_WR_USB_ADBUS_0_iv_13[1]\);
    
    \ELINK_DINA_15[1]\ : DFN1E0C0
      port map(D => \N_TFC_DINA[1]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_16, E => N_199, Q => 
        \ELINK_DINA_15[1]_net_1\);
    
    \ELINKS_STOP_ADDR_T[6]\ : DFN1E1C0
      port map(D => \RD_USB_ADBUS[6]_net_1\, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_7, E => 
        N_ELINKS_STOP_ADDR_T_0_sqmuxa, Q => 
        \ELINKS_STOP_ADDR_T[6]_net_1\);
    
    \WR_USB_ADBUS_RNO_23[1]\ : NOR2B
      port map(A => \ELINK_DOUTA_9[1]\, B => un1_SM_BANK_SEL_42, 
        Y => \ELINK_DOUTA_9_m[1]\);
    
    \REG_STATE_RNI3LQN[5]\ : NOR2A
      port map(A => \REG_STATE[2]_net_1\, B => 
        \REG_STATE[5]_net_1\, Y => N_1778);
    
    USB_RXF_B_RNIN32A2_0 : NOR2B
      port map(A => N_2537_1, B => N_446, Y => un1_USB_RXF_B_m);
    
    USB_RXF_B_0_RNI7BA26 : AO1
      port map(A => \USB_RXF_B_0\, B => N_2467, C => 
        REG_STATE_ns_i_245_tz_0, Y => N_1282_tz);
    
    \SM_BANK_SEL[8]\ : DFN1E1C0
      port map(D => N_1836, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_8, E => un1_REG_STATE_30, Q => 
        \SM_BANK_SEL[8]_net_1\);
    
    \ELINK_ADDRA_17[2]\ : DFN1E0C0
      port map(D => \N_TFC_ADDRA[2]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_10, E => N_197, Q => 
        \ELINK_ADDRA_17[2]_net_1\);
    
    \SM_BANK_SEL_RNIAL9D[10]\ : OR3A
      port map(A => N_461, B => \SM_BANK_SEL[11]_net_1\, C => 
        \SM_BANK_SEL[10]_net_1\, Y => \N_ELINK_RWA_0[10]\);
    
    \ELINK_DINA_11[6]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[6]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_11, E => un1_SM_BANK_SEL_16, Q => 
        \ELINK_DINA_11[6]_net_1\);
    
    \ELINK_BLKA_RNO[9]\ : OA1B
      port map(A => N_392, B => \ELINK_BLKA[9]_net_1\, C => N_164, 
        Y => \N_ELINK_BLKA_0_iv[9]\);
    
    \WR_USB_ADBUS_RNO_27[3]\ : AO1
      port map(A => \ELINK_DOUTA_12[3]\, B => un1_SM_BANK_SEL_33, 
        C => \ELINK_DOUTA_13_m[3]\, Y => 
        \N_WR_USB_ADBUS_0_iv_16[3]\);
    
    \REG_ADDR_RNILTTH7[6]\ : OAI1
      port map(A => REG_STATE_tr73_9, B => REG_STATE_tr74_1, C
         => N_1404_8, Y => N_2576);
    
    \ELINK_DINA_10[7]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[7]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_9, E => un1_SM_BANK_SEL_20, Q => 
        \ELINK_DINA_10[7]_net_1\);
    
    \ELINK_ADDRA_1[4]\ : DFN1E1C0
      port map(D => \N_TFC_ADDRA[4]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_20, E => un1_SM_BANK_SEL_19, Q => 
        \ELINK_ADDRA_1[4]_net_1\);
    
    \ELINKS_STRT_ADDR[6]\ : DFN1E1C0
      port map(D => \ELINKS_STRT_ADDR_T[6]_net_1\, CLK => 
        CLK60MHZ, CLR => P_USB_MASTER_EN_c_17, E => 
        \REG_STATE_d[30]\, Q => \ELINKS_STRT_ADDR[6]_net_1\);
    
    U105_PATT_ELINK_BLK : DPRT_512X9_SRAM_5
      port map(ELINK_RWA_0 => \ELINK_RWA[5]_net_1\, 
        ELK_RX_SER_WORD_5(7) => ELK_RX_SER_WORD_5(7), 
        ELK_RX_SER_WORD_5(6) => ELK_RX_SER_WORD_5(6), 
        ELK_RX_SER_WORD_5(5) => ELK_RX_SER_WORD_5(5), 
        ELK_RX_SER_WORD_5(4) => ELK_RX_SER_WORD_5(4), 
        ELK_RX_SER_WORD_5(3) => ELK_RX_SER_WORD_5(3), 
        ELK_RX_SER_WORD_5(2) => ELK_RX_SER_WORD_5(2), 
        ELK_RX_SER_WORD_5(1) => ELK_RX_SER_WORD_5(1), 
        ELK_RX_SER_WORD_5(0) => ELK_RX_SER_WORD_5(0), 
        ELINK_DINA_5(7) => \ELINK_DINA_5[7]_net_1\, 
        ELINK_DINA_5(6) => \ELINK_DINA_5[6]_net_1\, 
        ELINK_DINA_5(5) => \ELINK_DINA_5[5]_net_1\, 
        ELINK_DINA_5(4) => \ELINK_DINA_5[4]_net_1\, 
        ELINK_DINA_5(3) => \ELINK_DINA_5[3]_net_1\, 
        ELINK_DINA_5(2) => \ELINK_DINA_5[2]_net_1\, 
        ELINK_DINA_5(1) => \ELINK_DINA_5[1]_net_1\, 
        ELINK_DINA_5(0) => \ELINK_DINA_5[0]_net_1\, ELINK_BLKA_0
         => \ELINK_BLKA[5]_net_1\, ELKS_ADDRB_0_d0 => 
        ELKS_ADDRB(0), ELKS_ADDRB_1 => ELKS_ADDRB(1), 
        ELKS_ADDRB_3 => ELKS_ADDRB(3), ELKS_ADDRB_5 => 
        ELKS_ADDRB(5), ELKS_ADDRB_7 => ELKS_ADDRB(7), 
        ELKS_ADDRB_0_0 => ELKS_ADDRB_0_0, ELKS_ADDRB_0_2 => 
        ELKS_ADDRB_0_2, ELKS_ADDRB_0_4 => ELKS_ADDRB_0_4, 
        ELINK_ADDRA_5(7) => \ELINK_ADDRA_5[7]_net_1\, 
        ELINK_ADDRA_5(6) => \ELINK_ADDRA_5[6]_net_1\, 
        ELINK_ADDRA_5(5) => \ELINK_ADDRA_5[5]_net_1\, 
        ELINK_ADDRA_5(4) => \ELINK_ADDRA_5[4]_net_1\, 
        ELINK_ADDRA_5(3) => \ELINK_ADDRA_5[3]_net_1\, 
        ELINK_ADDRA_5(2) => \ELINK_ADDRA_5[2]_net_1\, 
        ELINK_ADDRA_5(1) => \ELINK_ADDRA_5[1]_net_1\, 
        ELINK_ADDRA_5(0) => \ELINK_ADDRA_5[0]_net_1\, 
        PATT_ELK_DAT_5(7) => PATT_ELK_DAT_5(7), PATT_ELK_DAT_5(6)
         => PATT_ELK_DAT_5(6), PATT_ELK_DAT_5(5) => 
        PATT_ELK_DAT_5(5), PATT_ELK_DAT_5(4) => PATT_ELK_DAT_5(4), 
        PATT_ELK_DAT_5(3) => PATT_ELK_DAT_5(3), PATT_ELK_DAT_5(2)
         => PATT_ELK_DAT_5(2), PATT_ELK_DAT_5(1) => 
        PATT_ELK_DAT_5(1), PATT_ELK_DAT_5(0) => PATT_ELK_DAT_5(0), 
        ELINK_DOUTA_5(7) => \ELINK_DOUTA_5[7]\, ELINK_DOUTA_5(6)
         => \ELINK_DOUTA_5[6]\, ELINK_DOUTA_5(5) => 
        \ELINK_DOUTA_5[5]\, ELINK_DOUTA_5(4) => 
        \ELINK_DOUTA_5[4]\, ELINK_DOUTA_5(3) => 
        \ELINK_DOUTA_5[3]\, ELINK_DOUTA_5(2) => 
        \ELINK_DOUTA_5[2]\, ELINK_DOUTA_5(1) => 
        \ELINK_DOUTA_5[1]\, ELINK_DOUTA_5(0) => 
        \ELINK_DOUTA_5[0]\, ELKS_RWB => ELKS_RWB, 
        P_USB_MASTER_EN_c_0 => P_USB_MASTER_EN_c_0, CLK_40M_GL
         => CLK_40M_GL, CLK60MHZ => CLK60MHZ, ELKS_RAM_BLKB_EN
         => ELKS_RAM_BLKB_EN);
    
    \ELINK_DINA_17[2]\ : DFN1E0C0
      port map(D => \N_TFC_DINA[2]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_19, E => N_197, Q => 
        \ELINK_DINA_17[2]_net_1\);
    
    \CHKSUM[6]\ : DFN1E1C0
      port map(D => N_228, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_4, E => un1_REG_STATE_22, Q => 
        \CHKSUM[6]_net_1\);
    
    \WR_USB_ADBUS_RNO_28[0]\ : AO1
      port map(A => \WR_XFER_TYPE[0]_net_1\, B => N_398, C => 
        \ELINKS_STOP_ADDR_m[0]\, Y => \N_WR_USB_ADBUS_0_iv_3[0]\);
    
    \REG_ADDR_RNITLRI1[6]\ : NOR2B
      port map(A => REG_ADDR_c5, B => \REG_ADDR[6]_net_1\, Y => 
        REG_ADDR_c6);
    
    \WR_USB_ADBUS_RNO_3[4]\ : AO1
      port map(A => \ELINK_DOUTA_10[4]\, B => un1_SM_BANK_SEL_34, 
        C => \ELINK_DOUTA_11_m[4]\, Y => 
        \N_WR_USB_ADBUS_0_iv_10[4]\);
    
    \SI_CNT_RNO[3]\ : XA1C
      port map(A => \SI_CNT[3]_net_1\, B => N_1630, C => N_678, Y
         => SI_CNT_n3);
    
    \RD_USB_ADBUS_RNIOEOG3[3]\ : NOR2B
      port map(A => N_1882, B => \RD_USB_ADBUS[3]_net_1\, Y => 
        N_1892);
    
    \SM_BANK_SEL_RNISJLS1[0]\ : OR3B
      port map(A => N_394, B => N_464, C => 
        \SM_BANK_SEL[0]_net_1\, Y => N_131);
    
    \REG_ADDR[6]\ : DFN1E1C0
      port map(D => REG_ADDR_n6, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_10, E => REG_ADDRe, Q => 
        \REG_ADDR[6]_net_1\);
    
    \REG_STATE_RNILG2AC[5]\ : OR2A
      port map(A => N_2576, B => N_1374, Y => 
        \REG_STATE_ns_i_i_0[0]\);
    
    \RD_XFER_TYPE_RNINJMR[0]\ : XOR2
      port map(A => \RD_XFER_TYPE[1]_net_1\, B => 
        \RD_XFER_TYPE[0]_net_1\, Y => N_262_i);
    
    \RD_XFER_TYPE_RNO[0]\ : AO1
      port map(A => \RD_XFER_TYPE[0]_net_1\, B => N_1703, C => 
        N_1794, Y => \RD_XFER_TYPE_RNO[0]_net_1\);
    
    \REG_STATE_RNI0RN31[5]\ : NOR2B
      port map(A => N_1352_1, B => \REG_STATE[5]_net_1\, Y => 
        N_2616);
    
    \ELINK_ADDRA_15[6]\ : DFN1E0C0
      port map(D => \N_TFC_ADDRA[6]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_6, E => N_199, Q => 
        \ELINK_ADDRA_15[6]_net_1\);
    
    \WR_USB_ADBUS_RNO_14[4]\ : NOR2B
      port map(A => \ELINK_DOUTA_13[4]\, B => un1_SM_BANK_SEL_29, 
        Y => \ELINK_DOUTA_13_m[4]\);
    
    \TFC_STOP_ADDR_T[0]\ : DFN1E1C0
      port map(D => \RD_USB_ADBUS[0]_net_1\, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_15, E => N_TFC_STOP_ADDR_T_0_sqmuxa, 
        Q => \TFC_STOP_ADDR_T[0]_net_1\);
    
    \ELINK_DINA_18[1]\ : DFN1E0C0
      port map(D => \N_TFC_DINA[1]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_21, E => N_198, Q => 
        \ELINK_DINA_18[1]_net_1\);
    
    \WR_USB_ADBUS_RNO_13[7]\ : NOR2B
      port map(A => \ELINK_DOUTA_1[7]\, B => un1_SM_BANK_SEL_36, 
        Y => \ELINK_DOUTA_1_m[7]\);
    
    \ELINK_DINA_2[5]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[5]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_9, E => un1_SM_BANK_SEL_5, Q => 
        \ELINK_DINA_2[5]_net_1\);
    
    \ELINK_DINA_3[7]\ : DFN1E1C0
      port map(D => \N_TFC_DINA[7]\, CLK => CLK60MHZ, CLR => 
        P_USB_MASTER_EN_c_11, E => un1_SM_BANK_SEL_4, Q => 
        \ELINK_DINA_3[7]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SYNC_DAT_SEL is

    port( TFC_TX_DAT             : out   std_logic_vector(7 downto 0);
          PATT_TFC_DAT           : in    std_logic_vector(7 downto 0);
          OP_MODE_c_0_0          : in    std_logic;
          MASTER_DCB_POR_B_i_0_i : in    std_logic;
          CLK_40M_GL             : in    std_logic
        );

end SYNC_DAT_SEL;

architecture DEF_ARCH of SYNC_DAT_SEL is 

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \N_SERDAT[0]\, \N_SERDAT[1]\, \N_SERDAT[2]\, 
        \N_SERDAT[3]\, \N_SERDAT[4]\, \N_SERDAT[5]\, 
        \N_SERDAT[6]\, \N_SERDAT[7]\, \GND\, \VCC\ : std_logic;

begin 


    \SERDAT_RNO[4]\ : NOR2A
      port map(A => PATT_TFC_DAT(4), B => OP_MODE_c_0_0, Y => 
        \N_SERDAT[4]\);
    
    \SERDAT_RNO[0]\ : NOR2A
      port map(A => PATT_TFC_DAT(0), B => OP_MODE_c_0_0, Y => 
        \N_SERDAT[0]\);
    
    \SERDAT[6]\ : DFN1C0
      port map(D => \N_SERDAT[6]\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => TFC_TX_DAT(6));
    
    \SERDAT[4]\ : DFN1C0
      port map(D => \N_SERDAT[4]\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => TFC_TX_DAT(4));
    
    \SERDAT_RNO[7]\ : OR2
      port map(A => PATT_TFC_DAT(7), B => OP_MODE_c_0_0, Y => 
        \N_SERDAT[7]\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \SERDAT_RNO[3]\ : OR2
      port map(A => PATT_TFC_DAT(3), B => OP_MODE_c_0_0, Y => 
        \N_SERDAT[3]\);
    
    \SERDAT_RNO[2]\ : OR2
      port map(A => PATT_TFC_DAT(2), B => OP_MODE_c_0_0, Y => 
        \N_SERDAT[2]\);
    
    \SERDAT[5]\ : DFN1C0
      port map(D => \N_SERDAT[5]\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => TFC_TX_DAT(5));
    
    \SERDAT[7]\ : DFN1C0
      port map(D => \N_SERDAT[7]\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => TFC_TX_DAT(7));
    
    GND_i : GND
      port map(Y => \GND\);
    
    \SERDAT_RNO[5]\ : NOR2A
      port map(A => PATT_TFC_DAT(5), B => OP_MODE_c_0_0, Y => 
        \N_SERDAT[5]\);
    
    \SERDAT[0]\ : DFN1C0
      port map(D => \N_SERDAT[0]\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => TFC_TX_DAT(0));
    
    \SERDAT_RNO[6]\ : NOR2A
      port map(A => PATT_TFC_DAT(6), B => OP_MODE_c_0_0, Y => 
        \N_SERDAT[6]\);
    
    \SERDAT[1]\ : DFN1C0
      port map(D => \N_SERDAT[1]\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => TFC_TX_DAT(1));
    
    \SERDAT_RNO[1]\ : OR2
      port map(A => PATT_TFC_DAT(1), B => OP_MODE_c_0_0, Y => 
        \N_SERDAT[1]\);
    
    \SERDAT[3]\ : DFN1C0
      port map(D => \N_SERDAT[3]\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => TFC_TX_DAT(3));
    
    \SERDAT[2]\ : DFN1C0
      port map(D => \N_SERDAT[2]\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => TFC_TX_DAT(2));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity CLK_FXD_40_160_A60M is

    port( USBCLK60MHZ_c    : in    std_logic;
          CCC_MAIN_LOCK    : out   std_logic;
          CLK60MHZ_1       : out   std_logic;
          CCC_160M_FXD_1   : out   std_logic;
          CLK_40M_GL_1     : out   std_logic;
          CLK_40M_BUF_RECD : in    std_logic
        );

end CLK_FXD_40_160_A60M;

architecture DEF_ARCH of CLK_FXD_40_160_A60M is 

  component DYNCCC
    generic (VCOFREQUENCY:real := 0.0);

    port( CLKA      : in    std_logic := 'U';
          EXTFB     : in    std_logic := 'U';
          POWERDOWN : in    std_logic := 'U';
          GLA       : out   std_logic;
          LOCK      : out   std_logic;
          CLKB      : in    std_logic := 'U';
          GLB       : out   std_logic;
          YB        : out   std_logic;
          CLKC      : in    std_logic := 'U';
          GLC       : out   std_logic;
          YC        : out   std_logic;
          SDIN      : in    std_logic := 'U';
          SCLK      : in    std_logic := 'U';
          SSHIFT    : in    std_logic := 'U';
          SUPDATE   : in    std_logic := 'U';
          MODE      : in    std_logic := 'U';
          SDOUT     : out   std_logic;
          OADIV0    : in    std_logic := 'U';
          OADIV1    : in    std_logic := 'U';
          OADIV2    : in    std_logic := 'U';
          OADIV3    : in    std_logic := 'U';
          OADIV4    : in    std_logic := 'U';
          OAMUX0    : in    std_logic := 'U';
          OAMUX1    : in    std_logic := 'U';
          OAMUX2    : in    std_logic := 'U';
          DLYGLA0   : in    std_logic := 'U';
          DLYGLA1   : in    std_logic := 'U';
          DLYGLA2   : in    std_logic := 'U';
          DLYGLA3   : in    std_logic := 'U';
          DLYGLA4   : in    std_logic := 'U';
          OBDIV0    : in    std_logic := 'U';
          OBDIV1    : in    std_logic := 'U';
          OBDIV2    : in    std_logic := 'U';
          OBDIV3    : in    std_logic := 'U';
          OBDIV4    : in    std_logic := 'U';
          OBMUX0    : in    std_logic := 'U';
          OBMUX1    : in    std_logic := 'U';
          OBMUX2    : in    std_logic := 'U';
          DLYYB0    : in    std_logic := 'U';
          DLYYB1    : in    std_logic := 'U';
          DLYYB2    : in    std_logic := 'U';
          DLYYB3    : in    std_logic := 'U';
          DLYYB4    : in    std_logic := 'U';
          DLYGLB0   : in    std_logic := 'U';
          DLYGLB1   : in    std_logic := 'U';
          DLYGLB2   : in    std_logic := 'U';
          DLYGLB3   : in    std_logic := 'U';
          DLYGLB4   : in    std_logic := 'U';
          OCDIV0    : in    std_logic := 'U';
          OCDIV1    : in    std_logic := 'U';
          OCDIV2    : in    std_logic := 'U';
          OCDIV3    : in    std_logic := 'U';
          OCDIV4    : in    std_logic := 'U';
          OCMUX0    : in    std_logic := 'U';
          OCMUX1    : in    std_logic := 'U';
          OCMUX2    : in    std_logic := 'U';
          DLYYC0    : in    std_logic := 'U';
          DLYYC1    : in    std_logic := 'U';
          DLYYC2    : in    std_logic := 'U';
          DLYYC3    : in    std_logic := 'U';
          DLYYC4    : in    std_logic := 'U';
          DLYGLC0   : in    std_logic := 'U';
          DLYGLC1   : in    std_logic := 'U';
          DLYGLC2   : in    std_logic := 'U';
          DLYGLC3   : in    std_logic := 'U';
          DLYGLC4   : in    std_logic := 'U';
          FINDIV0   : in    std_logic := 'U';
          FINDIV1   : in    std_logic := 'U';
          FINDIV2   : in    std_logic := 'U';
          FINDIV3   : in    std_logic := 'U';
          FINDIV4   : in    std_logic := 'U';
          FINDIV5   : in    std_logic := 'U';
          FINDIV6   : in    std_logic := 'U';
          FBDIV0    : in    std_logic := 'U';
          FBDIV1    : in    std_logic := 'U';
          FBDIV2    : in    std_logic := 'U';
          FBDIV3    : in    std_logic := 'U';
          FBDIV4    : in    std_logic := 'U';
          FBDIV5    : in    std_logic := 'U';
          FBDIV6    : in    std_logic := 'U';
          FBDLY0    : in    std_logic := 'U';
          FBDLY1    : in    std_logic := 'U';
          FBDLY2    : in    std_logic := 'U';
          FBDLY3    : in    std_logic := 'U';
          FBDLY4    : in    std_logic := 'U';
          FBSEL0    : in    std_logic := 'U';
          FBSEL1    : in    std_logic := 'U';
          XDLYSEL   : in    std_logic := 'U';
          VCOSEL0   : in    std_logic := 'U';
          VCOSEL1   : in    std_logic := 'U';
          VCOSEL2   : in    std_logic := 'U'
        );
  end component;

  component PLLINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal CLKAP, SDOUT, Core_YB_0, Core_YC_0, 
        CLK_FXD_40_160_A60M_GND, CLKCP, CLK_FXD_40_160_A60M_VCC
         : std_logic;

begin 


    Core : DYNCCC
      generic map(VCOFREQUENCY => 160.0)

      port map(CLKA => CLKAP, EXTFB => CLK_FXD_40_160_A60M_GND, 
        POWERDOWN => CLK_FXD_40_160_A60M_VCC, GLA => CLK_40M_GL_1, 
        LOCK => CCC_MAIN_LOCK, CLKB => CLK_FXD_40_160_A60M_GND, 
        GLB => CCC_160M_FXD_1, YB => Core_YB_0, CLKC => CLKCP, 
        GLC => CLK60MHZ_1, YC => Core_YC_0, SDIN => 
        CLK_FXD_40_160_A60M_GND, SCLK => CLK_FXD_40_160_A60M_GND, 
        SSHIFT => CLK_FXD_40_160_A60M_GND, SUPDATE => 
        CLK_FXD_40_160_A60M_GND, MODE => CLK_FXD_40_160_A60M_GND, 
        SDOUT => SDOUT, OADIV0 => CLK_FXD_40_160_A60M_VCC, OADIV1
         => CLK_FXD_40_160_A60M_VCC, OADIV2 => 
        CLK_FXD_40_160_A60M_GND, OADIV3 => 
        CLK_FXD_40_160_A60M_GND, OADIV4 => 
        CLK_FXD_40_160_A60M_GND, OAMUX0 => 
        CLK_FXD_40_160_A60M_GND, OAMUX1 => 
        CLK_FXD_40_160_A60M_GND, OAMUX2 => 
        CLK_FXD_40_160_A60M_VCC, DLYGLA0 => 
        CLK_FXD_40_160_A60M_GND, DLYGLA1 => 
        CLK_FXD_40_160_A60M_GND, DLYGLA2 => 
        CLK_FXD_40_160_A60M_GND, DLYGLA3 => 
        CLK_FXD_40_160_A60M_GND, DLYGLA4 => 
        CLK_FXD_40_160_A60M_GND, OBDIV0 => 
        CLK_FXD_40_160_A60M_GND, OBDIV1 => 
        CLK_FXD_40_160_A60M_GND, OBDIV2 => 
        CLK_FXD_40_160_A60M_GND, OBDIV3 => 
        CLK_FXD_40_160_A60M_GND, OBDIV4 => 
        CLK_FXD_40_160_A60M_GND, OBMUX0 => 
        CLK_FXD_40_160_A60M_GND, OBMUX1 => 
        CLK_FXD_40_160_A60M_GND, OBMUX2 => 
        CLK_FXD_40_160_A60M_VCC, DLYYB0 => 
        CLK_FXD_40_160_A60M_GND, DLYYB1 => 
        CLK_FXD_40_160_A60M_GND, DLYYB2 => 
        CLK_FXD_40_160_A60M_GND, DLYYB3 => 
        CLK_FXD_40_160_A60M_GND, DLYYB4 => 
        CLK_FXD_40_160_A60M_GND, DLYGLB0 => 
        CLK_FXD_40_160_A60M_GND, DLYGLB1 => 
        CLK_FXD_40_160_A60M_GND, DLYGLB2 => 
        CLK_FXD_40_160_A60M_VCC, DLYGLB3 => 
        CLK_FXD_40_160_A60M_VCC, DLYGLB4 => 
        CLK_FXD_40_160_A60M_GND, OCDIV0 => 
        CLK_FXD_40_160_A60M_GND, OCDIV1 => 
        CLK_FXD_40_160_A60M_GND, OCDIV2 => 
        CLK_FXD_40_160_A60M_GND, OCDIV3 => 
        CLK_FXD_40_160_A60M_GND, OCDIV4 => 
        CLK_FXD_40_160_A60M_GND, OCMUX0 => 
        CLK_FXD_40_160_A60M_GND, OCMUX1 => 
        CLK_FXD_40_160_A60M_GND, OCMUX2 => 
        CLK_FXD_40_160_A60M_GND, DLYYC0 => 
        CLK_FXD_40_160_A60M_GND, DLYYC1 => 
        CLK_FXD_40_160_A60M_GND, DLYYC2 => 
        CLK_FXD_40_160_A60M_GND, DLYYC3 => 
        CLK_FXD_40_160_A60M_GND, DLYYC4 => 
        CLK_FXD_40_160_A60M_GND, DLYGLC0 => 
        CLK_FXD_40_160_A60M_VCC, DLYGLC1 => 
        CLK_FXD_40_160_A60M_GND, DLYGLC2 => 
        CLK_FXD_40_160_A60M_VCC, DLYGLC3 => 
        CLK_FXD_40_160_A60M_VCC, DLYGLC4 => 
        CLK_FXD_40_160_A60M_VCC, FINDIV0 => 
        CLK_FXD_40_160_A60M_VCC, FINDIV1 => 
        CLK_FXD_40_160_A60M_VCC, FINDIV2 => 
        CLK_FXD_40_160_A60M_VCC, FINDIV3 => 
        CLK_FXD_40_160_A60M_GND, FINDIV4 => 
        CLK_FXD_40_160_A60M_GND, FINDIV5 => 
        CLK_FXD_40_160_A60M_GND, FINDIV6 => 
        CLK_FXD_40_160_A60M_GND, FBDIV0 => 
        CLK_FXD_40_160_A60M_VCC, FBDIV1 => 
        CLK_FXD_40_160_A60M_VCC, FBDIV2 => 
        CLK_FXD_40_160_A60M_VCC, FBDIV3 => 
        CLK_FXD_40_160_A60M_VCC, FBDIV4 => 
        CLK_FXD_40_160_A60M_VCC, FBDIV5 => 
        CLK_FXD_40_160_A60M_GND, FBDIV6 => 
        CLK_FXD_40_160_A60M_GND, FBDLY0 => 
        CLK_FXD_40_160_A60M_GND, FBDLY1 => 
        CLK_FXD_40_160_A60M_GND, FBDLY2 => 
        CLK_FXD_40_160_A60M_VCC, FBDLY3 => 
        CLK_FXD_40_160_A60M_GND, FBDLY4 => 
        CLK_FXD_40_160_A60M_GND, FBSEL0 => 
        CLK_FXD_40_160_A60M_GND, FBSEL1 => 
        CLK_FXD_40_160_A60M_VCC, XDLYSEL => 
        CLK_FXD_40_160_A60M_GND, VCOSEL0 => 
        CLK_FXD_40_160_A60M_GND, VCOSEL1 => 
        CLK_FXD_40_160_A60M_GND, VCOSEL2 => 
        CLK_FXD_40_160_A60M_VCC);
    
    pllint1 : PLLINT
      port map(A => CLK_40M_BUF_RECD, Y => CLKAP);
    
    VCC_i : VCC
      port map(Y => CLK_FXD_40_160_A60M_VCC);
    
    pllint3 : PLLINT
      port map(A => USBCLK60MHZ_c, Y => CLKCP);
    
    GND_i : GND
      port map(Y => CLK_FXD_40_160_A60M_GND);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SLAVE_DES320S_1_17_16 is

    port( ELK_RX_SER_WORD_18     : out   std_logic_vector(7 downto 0);
          BIT_OS_SEL_2           : in    std_logic_vector(1 downto 0);
          BIT_OS_SEL_1           : in    std_logic_vector(2 downto 1);
          BIT_OS_SEL_0           : in    std_logic_vector(2 downto 1);
          CLK_40M_GL             : in    std_logic;
          CCC_160M_FXD           : in    std_logic;
          ELK_IN_R               : in    std_logic;
          ELK_IN_F               : in    std_logic;
          MASTER_DCB_POR_B_i_0_i : in    std_logic;
          CCC_160M_ADJ           : in    std_logic
        );

end SLAVE_DES320S_1_17_16;

architecture DEF_ARCH of SLAVE_DES320S_1_17_16 is 

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal N_17, \ARB_BYTE[0]_net_1\, \ARB_BYTE[4]_net_1\, N_18, 
        \ARB_BYTE[1]_net_1\, \ARB_BYTE[5]_net_1\, N_19, 
        \ARB_BYTE[2]_net_1\, \ARB_BYTE[6]_net_1\, N_20, 
        \ARB_BYTE[3]_net_1\, \ARB_BYTE[7]_net_1\, N_21, 
        \ARB_BYTE[8]_net_1\, N_22, \ARB_BYTE[9]_net_1\, N_23, 
        \ARB_BYTE[10]_net_1\, N_24, \ARB_BYTE[11]_net_1\, N_31, 
        \ARB_BYTE[12]_net_1\, N_32, \ARB_BYTE[13]_net_1\, N_33, 
        N_34, N_35, N_36, N_37, N_38, N_39, N_40, N_56, 
        \ARB_BYTE[14]_net_1\, N_64, \N_RECD_SER_WORD[0]\, 
        \N_RECD_SER_WORD[1]\, \N_RECD_SER_WORD[2]\, 
        \N_RECD_SER_WORD[3]\, \N_RECD_SER_WORD[4]\, 
        \N_RECD_SER_WORD[5]\, \N_RECD_SER_WORD[6]\, 
        \N_RECD_SER_WORD[7]\, \ADJ_SER_IN_F_0DEL\, 
        \ADJ_SER_IN_R_0DEL\, \ADJ_SER_IN_F_1DEL\, 
        \ADJ_SER_IN_R_1DEL\, \Q[0]_net_1\, \ADJ_Q[0]_net_1\, 
        \Q[1]_net_1\, \ADJ_Q[1]_net_1\, \Q[2]_net_1\, 
        \ADJ_Q[2]_net_1\, \Q[3]_net_1\, \ADJ_Q[3]_net_1\, 
        \Q[4]_net_1\, \ADJ_Q[4]_net_1\, \Q[5]_net_1\, 
        \ADJ_Q[5]_net_1\, \Q[6]_net_1\, \ADJ_Q[6]_net_1\, 
        \Q[7]_net_1\, \ADJ_Q[7]_net_1\, \Q[8]_net_1\, 
        \ADJ_Q[8]_net_1\, \Q[9]_net_1\, \ADJ_Q[9]_net_1\, 
        \Q[10]_net_1\, \ADJ_Q[10]_net_1\, \Q[11]_net_1\, 
        \ADJ_Q[11]_net_1\, \Q[12]_net_1\, \ADJ_Q[12]_net_1\, 
        \Q[13]_net_1\, \ADJ_Q[13]_net_1\, \Q[14]_net_1\, 
        \ADJ_Q[14]_net_1\, \ARB_WRD_40M_FIXED[0]_net_1\, 
        \ARB_WRD_40M_FIXED[1]_net_1\, 
        \ARB_WRD_40M_FIXED[2]_net_1\, 
        \ARB_WRD_40M_FIXED[3]_net_1\, 
        \ARB_WRD_40M_FIXED[4]_net_1\, 
        \ARB_WRD_40M_FIXED[5]_net_1\, 
        \ARB_WRD_40M_FIXED[6]_net_1\, 
        \ARB_WRD_40M_FIXED[7]_net_1\, 
        \ARB_WRD_40M_FIXED[8]_net_1\, 
        \ARB_WRD_40M_FIXED[9]_net_1\, 
        \ARB_WRD_40M_FIXED[10]_net_1\, 
        \ARB_WRD_40M_FIXED[11]_net_1\, 
        \ARB_WRD_40M_FIXED[12]_net_1\, 
        \ARB_WRD_40M_FIXED[13]_net_1\, 
        \ARB_WRD_40M_FIXED[14]_net_1\, \GND\, \VCC\ : std_logic;

begin 


    \RECD_SER_WORD_RNO[5]\ : MX2
      port map(A => N_38, B => N_39, S => BIT_OS_SEL_2(0), Y => 
        \N_RECD_SER_WORD[5]\);
    
    \ARB_WRD_40M_FIXED[9]\ : DFN1C0
      port map(D => \Q[9]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[9]_net_1\);
    
    \ADJ_Q[4]\ : DFN1C0
      port map(D => \ADJ_Q[2]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[4]_net_1\);
    
    \ARB_BYTE[6]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[6]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[6]_net_1\);
    
    ADJ_SER_IN_F_1DEL : DFN1C0
      port map(D => \ADJ_SER_IN_F_0DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_F_1DEL\);
    
    \ARB_BYTE[0]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[0]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[0]_net_1\);
    
    \Q[11]\ : DFN1C0
      port map(D => \ADJ_Q[11]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[11]_net_1\);
    
    \ADJ_Q[8]\ : DFN1C0
      port map(D => \ADJ_Q[6]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[8]_net_1\);
    
    \ARB_BYTE_RNICK681[4]\ : MX2
      port map(A => \ARB_BYTE[4]_net_1\, B => \ARB_BYTE[8]_net_1\, 
        S => BIT_OS_SEL_0(2), Y => N_21);
    
    \ARB_BYTE_RNIU6QV2[6]\ : MX2
      port map(A => N_23, B => N_31, S => BIT_OS_SEL_1(1), Y => 
        N_39);
    
    \ADJ_Q[6]\ : DFN1C0
      port map(D => \ADJ_Q[4]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[6]_net_1\);
    
    \ADJ_Q[12]\ : DFN1C0
      port map(D => \ADJ_Q[10]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[12]_net_1\);
    
    \RECD_SER_WORD_RNO_1[0]\ : MX2
      port map(A => \ARB_BYTE[0]_net_1\, B => \ARB_BYTE[4]_net_1\, 
        S => BIT_OS_SEL_0(2), Y => N_17);
    
    \Q[1]\ : DFN1C0
      port map(D => \ADJ_Q[1]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[1]_net_1\);
    
    \ARB_BYTE_RNI8G681[2]\ : MX2
      port map(A => \ARB_BYTE[2]_net_1\, B => \ARB_BYTE[6]_net_1\, 
        S => BIT_OS_SEL_0(2), Y => N_19);
    
    \ARB_BYTE[4]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[4]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[4]_net_1\);
    
    \ADJ_Q[2]\ : DFN1C0
      port map(D => \ADJ_Q[0]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[2]_net_1\);
    
    \RECD_SER_WORD_RNO_1[7]\ : MX2
      port map(A => \ARB_BYTE[10]_net_1\, B => 
        \ARB_BYTE[14]_net_1\, S => BIT_OS_SEL_1(2), Y => N_56);
    
    \RECD_SER_WORD[4]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[4]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_18(4));
    
    \Q[5]\ : DFN1C0
      port map(D => \ADJ_Q[5]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[5]_net_1\);
    
    \ADJ_Q[11]\ : DFN1C0
      port map(D => \ADJ_Q[9]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[11]_net_1\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \ADJ_Q[3]\ : DFN1C0
      port map(D => \ADJ_Q[1]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[3]_net_1\);
    
    \Q[10]\ : DFN1C0
      port map(D => \ADJ_Q[10]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[10]_net_1\);
    
    \ARB_WRD_40M_FIXED[6]\ : DFN1C0
      port map(D => \Q[6]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[6]_net_1\);
    
    \ARB_WRD_40M_FIXED[1]\ : DFN1C0
      port map(D => \Q[1]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[1]_net_1\);
    
    \RECD_SER_WORD[3]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[3]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_18(3));
    
    \ARB_BYTE_RNI3BJU2[3]\ : MX2
      port map(A => N_20, B => N_22, S => BIT_OS_SEL_0(1), Y => 
        N_36);
    
    \RECD_SER_WORD[0]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[0]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_18(0));
    
    \RECD_SER_WORD_RNO[3]\ : MX2
      port map(A => N_36, B => N_37, S => BIT_OS_SEL_2(0), Y => 
        \N_RECD_SER_WORD[3]\);
    
    \Q[0]\ : DFN1C0
      port map(D => \ADJ_Q[0]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[0]_net_1\);
    
    \RECD_SER_WORD_RNO_0[7]\ : MX2
      port map(A => N_31, B => N_56, S => BIT_OS_SEL_2(1), Y => 
        N_64);
    
    \Q[7]\ : DFN1C0
      port map(D => \ADJ_Q[7]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[7]_net_1\);
    
    \ARB_BYTE[14]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[14]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[14]_net_1\);
    
    \ARB_WRD_40M_FIXED[2]\ : DFN1C0
      port map(D => \Q[2]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[2]_net_1\);
    
    \ARB_WRD_40M_FIXED[14]\ : DFN1C0
      port map(D => \Q[14]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[14]_net_1\);
    
    \RECD_SER_WORD_RNO[2]\ : MX2
      port map(A => N_35, B => N_36, S => BIT_OS_SEL_2(0), Y => 
        \N_RECD_SER_WORD[2]\);
    
    \ARB_BYTE[2]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[2]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[2]_net_1\);
    
    \ADJ_Q[7]\ : DFN1C0
      port map(D => \ADJ_Q[5]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[7]_net_1\);
    
    \ARB_BYTE_RNIJCOV2[5]\ : MX2
      port map(A => N_22, B => N_24, S => BIT_OS_SEL_1(1), Y => 
        N_38);
    
    \ARB_BYTE[8]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[8]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[8]_net_1\);
    
    \RECD_SER_WORD[5]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[5]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_18(5));
    
    \ARB_BYTE[12]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[12]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[12]_net_1\);
    
    \RECD_SER_WORD[1]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[1]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_18(1));
    
    \ARB_BYTE_RNI2BQV2[13]\ : MX2
      port map(A => N_24, B => N_32, S => BIT_OS_SEL_1(1), Y => 
        N_40);
    
    \Q[3]\ : DFN1C0
      port map(D => \ADJ_Q[3]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[3]_net_1\);
    
    \ARB_BYTE_RNINE881[6]\ : MX2
      port map(A => \ARB_BYTE[6]_net_1\, B => 
        \ARB_BYTE[10]_net_1\, S => BIT_OS_SEL_0(2), Y => N_23);
    
    ADJ_SER_IN_F_0DEL : DFN1C0
      port map(D => ELK_IN_F, CLK => CCC_160M_ADJ, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_F_0DEL\);
    
    \RECD_SER_WORD_RNO[7]\ : MX2
      port map(A => N_40, B => N_64, S => BIT_OS_SEL_2(0), Y => 
        \N_RECD_SER_WORD[7]\);
    
    \RECD_SER_WORD_RNO[1]\ : MX2
      port map(A => N_34, B => N_35, S => BIT_OS_SEL_2(0), Y => 
        \N_RECD_SER_WORD[1]\);
    
    \ARB_WRD_40M_FIXED[4]\ : DFN1C0
      port map(D => \Q[4]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[4]_net_1\);
    
    \RECD_SER_WORD_RNO[0]\ : MX2
      port map(A => N_33, B => N_34, S => BIT_OS_SEL_2(0), Y => 
        \N_RECD_SER_WORD[0]\);
    
    \Q[6]\ : DFN1C0
      port map(D => \ADJ_Q[6]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[6]_net_1\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \ARB_WRD_40M_FIXED[8]\ : DFN1C0
      port map(D => \Q[8]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[8]_net_1\);
    
    \ARB_BYTE_RNITK881[13]\ : MX2
      port map(A => \ARB_BYTE[9]_net_1\, B => 
        \ARB_BYTE[13]_net_1\, S => BIT_OS_SEL_0(2), Y => N_32);
    
    \ARB_BYTE[11]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[11]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[11]_net_1\);
    
    \Q[9]\ : DFN1C0
      port map(D => \ADJ_Q[9]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[9]_net_1\);
    
    \ARB_BYTE_RNIV6JU2[2]\ : MX2
      port map(A => N_19, B => N_21, S => BIT_OS_SEL_0(1), Y => 
        N_35);
    
    \Q[14]\ : DFN1C0
      port map(D => \ADJ_Q[14]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[14]_net_1\);
    
    ADJ_SER_IN_R_0DEL : DFN1C0
      port map(D => ELK_IN_R, CLK => CCC_160M_ADJ, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_R_0DEL\);
    
    \Q[13]\ : DFN1C0
      port map(D => \ADJ_Q[13]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[13]_net_1\);
    
    \ARB_BYTE[9]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[9]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[9]_net_1\);
    
    ADJ_SER_IN_R_1DEL : DFN1C0
      port map(D => \ADJ_SER_IN_R_0DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_R_1DEL\);
    
    \ARB_BYTE[10]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[10]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[10]_net_1\);
    
    \ADJ_Q[9]\ : DFN1C0
      port map(D => \ADJ_Q[7]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[9]_net_1\);
    
    \RECD_SER_WORD[7]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[7]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_18(7));
    
    \ARB_WRD_40M_FIXED[5]\ : DFN1C0
      port map(D => \Q[5]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[5]_net_1\);
    
    \ARB_WRD_40M_FIXED[12]\ : DFN1C0
      port map(D => \Q[12]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[12]_net_1\);
    
    \ARB_WRD_40M_FIXED[11]\ : DFN1C0
      port map(D => \Q[11]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[11]_net_1\);
    
    \ARB_BYTE_RNIPG881[11]\ : MX2
      port map(A => \ARB_BYTE[7]_net_1\, B => 
        \ARB_BYTE[11]_net_1\, S => BIT_OS_SEL_0(2), Y => N_24);
    
    \ARB_WRD_40M_FIXED[0]\ : DFN1C0
      port map(D => \Q[0]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[0]_net_1\);
    
    \ARB_BYTE_RNIEM681[5]\ : MX2
      port map(A => \ARB_BYTE[5]_net_1\, B => \ARB_BYTE[9]_net_1\, 
        S => BIT_OS_SEL_0(2), Y => N_22);
    
    \ADJ_Q[10]\ : DFN1C0
      port map(D => \ADJ_Q[8]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[10]_net_1\);
    
    \Q[2]\ : DFN1C0
      port map(D => \ADJ_Q[2]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[2]_net_1\);
    
    \ARB_BYTE_RNIR2JU2[1]\ : MX2
      port map(A => N_18, B => N_20, S => BIT_OS_SEL_0(1), Y => 
        N_34);
    
    \ADJ_Q[1]\ : DFN1C0
      port map(D => \ADJ_SER_IN_F_1DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[1]_net_1\);
    
    \RECD_SER_WORD[6]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[6]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_18(6));
    
    \RECD_SER_WORD[2]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[2]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_18(2));
    
    \ADJ_Q[13]\ : DFN1C0
      port map(D => \ADJ_Q[11]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[13]_net_1\);
    
    \Q[8]\ : DFN1C0
      port map(D => \ADJ_Q[8]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[8]_net_1\);
    
    \ARB_BYTE[5]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[5]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[5]_net_1\);
    
    \ADJ_Q[14]\ : DFN1C0
      port map(D => \ADJ_Q[12]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[14]_net_1\);
    
    \RECD_SER_WORD_RNO[4]\ : MX2
      port map(A => N_37, B => N_38, S => BIT_OS_SEL_2(0), Y => 
        \N_RECD_SER_WORD[4]\);
    
    \Q[12]\ : DFN1C0
      port map(D => \ADJ_Q[12]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[12]_net_1\);
    
    \ARB_BYTE[13]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[13]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[13]_net_1\);
    
    \ARB_WRD_40M_FIXED[3]\ : DFN1C0
      port map(D => \Q[3]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[3]_net_1\);
    
    \ARB_BYTE[7]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[7]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[7]_net_1\);
    
    \RECD_SER_WORD_RNO_0[0]\ : MX2
      port map(A => N_17, B => N_19, S => BIT_OS_SEL_0(1), Y => 
        N_33);
    
    \ARB_BYTE_RNI6E681[1]\ : MX2
      port map(A => \ARB_BYTE[1]_net_1\, B => \ARB_BYTE[5]_net_1\, 
        S => BIT_OS_SEL_0(2), Y => N_18);
    
    \Q[4]\ : DFN1C0
      port map(D => \ADJ_Q[4]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[4]_net_1\);
    
    \ARB_WRD_40M_FIXED[7]\ : DFN1C0
      port map(D => \Q[7]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[7]_net_1\);
    
    \ARB_BYTE_RNIAI681[3]\ : MX2
      port map(A => \ARB_BYTE[3]_net_1\, B => \ARB_BYTE[7]_net_1\, 
        S => BIT_OS_SEL_0(2), Y => N_20);
    
    \RECD_SER_WORD_RNO[6]\ : MX2
      port map(A => N_39, B => N_40, S => BIT_OS_SEL_2(0), Y => 
        \N_RECD_SER_WORD[6]\);
    
    \ARB_BYTE_RNIRI881[12]\ : MX2
      port map(A => \ARB_BYTE[8]_net_1\, B => 
        \ARB_BYTE[12]_net_1\, S => BIT_OS_SEL_0(2), Y => N_31);
    
    \ARB_BYTE_RNIE5LU2[4]\ : MX2
      port map(A => N_21, B => N_23, S => BIT_OS_SEL_0(1), Y => 
        N_37);
    
    \ARB_BYTE[3]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[3]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[3]_net_1\);
    
    \ADJ_Q[5]\ : DFN1C0
      port map(D => \ADJ_Q[3]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[5]_net_1\);
    
    \ARB_BYTE[1]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[1]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[1]_net_1\);
    
    \ARB_WRD_40M_FIXED[13]\ : DFN1C0
      port map(D => \Q[13]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[13]_net_1\);
    
    \ADJ_Q[0]\ : DFN1C0
      port map(D => \ADJ_SER_IN_R_1DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[0]_net_1\);
    
    \ARB_WRD_40M_FIXED[10]\ : DFN1C0
      port map(D => \Q[10]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[10]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SER320M_3_34_18 is

    port( ELK_TX_DAT                 : in    std_logic_vector(7 downto 0);
          MASTER_SALT_POR_B_i_0_i_0  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_3  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_17 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_1  : in    std_logic;
          ELK_OUT_R                  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_4  : in    std_logic;
          ELK_OUT_F                  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_9  : in    std_logic;
          CCC_160M_FXD               : in    std_logic;
          CLK_40M_GL                 : in    std_logic
        );

end SER320M_3_34_18;

architecture DEF_ARCH of SER320M_3_34_18 is 

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \N_SER_CMD_WORD_R[0]\, \START_RISE\, 
        \N_SER_CMD_WORD_F[0]\, \N_SER_CMD_WORD_R[3]\, 
        \SER_CMD_WORD_R[2]_net_1\, \N_SER_CMD_WORD_R[2]\, 
        \SER_CMD_WORD_R[1]_net_1\, \N_SER_CMD_WORD_R[1]\, 
        \SER_CMD_WORD_R[0]_net_1\, \N_SER_CMD_WORD_F[3]\, 
        \SER_CMD_WORD_F[2]_net_1\, \N_SER_CMD_WORD_F[2]\, 
        \SER_CMD_WORD_F[1]_net_1\, \N_SER_CMD_WORD_F[1]\, 
        \SER_CMD_WORD_F[0]_net_1\, N_START_RISE, 
        \CLK40M_GEN_DEL0\, \SER_OUT_FI\, \SER_OUT_RI\, 
        \SER_CMD_WORD_F[3]_net_1\, \SER_CMD_WORD_R[3]_net_1\, 
        \GND\, \VCC\ : std_logic;

begin 


    SER_OUT_FI : DFN1C0
      port map(D => \SER_CMD_WORD_F[3]_net_1\, CLK => 
        CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_9, Q => 
        \SER_OUT_FI\);
    
    \SER_CMD_WORD_F[3]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[3]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_3, Q => 
        \SER_CMD_WORD_F[3]_net_1\);
    
    \SER_CMD_WORD_R[1]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[1]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_0, Q => 
        \SER_CMD_WORD_R[1]_net_1\);
    
    \SER_CMD_WORD_R[2]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[2]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_0, Q => 
        \SER_CMD_WORD_R[2]_net_1\);
    
    \SER_CMD_WORD_R_RNO[3]\ : MX2
      port map(A => \SER_CMD_WORD_R[2]_net_1\, B => ELK_TX_DAT(7), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_R[3]\);
    
    \SER_CMD_WORD_R_RNO[0]\ : NOR2B
      port map(A => \START_RISE\, B => ELK_TX_DAT(1), Y => 
        \N_SER_CMD_WORD_R[0]\);
    
    \SER_CMD_WORD_F[0]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[0]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_3, Q => 
        \SER_CMD_WORD_F[0]_net_1\);
    
    \SER_CMD_WORD_R_RNO[1]\ : MX2
      port map(A => \SER_CMD_WORD_R[0]_net_1\, B => ELK_TX_DAT(3), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_R[1]\);
    
    \SER_CMD_WORD_F_RNO[2]\ : MX2
      port map(A => \SER_CMD_WORD_F[1]_net_1\, B => ELK_TX_DAT(4), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_F[2]\);
    
    \SER_CMD_WORD_F_RNO[3]\ : MX2
      port map(A => \SER_CMD_WORD_F[2]_net_1\, B => ELK_TX_DAT(6), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_F[3]\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    CLK40M_GEN_DEL0 : DFN1C0
      port map(D => CLK_40M_GL, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_9, Q => \CLK40M_GEN_DEL0\);
    
    SER_OUT_RI : DFN1C0
      port map(D => \SER_CMD_WORD_R[3]_net_1\, CLK => 
        CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_9, Q => 
        \SER_OUT_RI\);
    
    \SER_CMD_WORD_F[2]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[2]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_3, Q => 
        \SER_CMD_WORD_F[2]_net_1\);
    
    \SER_CMD_WORD_F_RNO[1]\ : MX2
      port map(A => \SER_CMD_WORD_F[0]_net_1\, B => ELK_TX_DAT(2), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_F[1]\);
    
    \SER_CMD_WORD_R[0]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[0]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_0, Q => 
        \SER_CMD_WORD_R[0]_net_1\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    START_RISE : DFN1C0
      port map(D => N_START_RISE, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_17, Q => \START_RISE\);
    
    \SER_CMD_WORD_R[3]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[3]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_0, Q => 
        \SER_CMD_WORD_R[3]_net_1\);
    
    \SER_CMD_WORD_F_RNO[0]\ : NOR2B
      port map(A => \START_RISE\, B => ELK_TX_DAT(0), Y => 
        \N_SER_CMD_WORD_F[0]\);
    
    SER_OUT_RDEL : DFN1C0
      port map(D => \SER_OUT_RI\, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_1, Q => ELK_OUT_R);
    
    \SER_CMD_WORD_F[1]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[1]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_3, Q => 
        \SER_CMD_WORD_F[1]_net_1\);
    
    START_RISE_RNO : NOR2B
      port map(A => \CLK40M_GEN_DEL0\, B => CLK_40M_GL, Y => 
        N_START_RISE);
    
    \SER_CMD_WORD_R_RNO[2]\ : MX2
      port map(A => \SER_CMD_WORD_R[1]_net_1\, B => ELK_TX_DAT(5), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_R[2]\);
    
    SER_OUT_FDEL : DFN1C0
      port map(D => \SER_OUT_FI\, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_4, Q => ELK_OUT_F);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity DDR_BIDIR_LVDS_DUAL_CLK_18 is

    port( DCB_SALT_SEL_c_i : in    std_logic;
          ELK18_DAT_P      : inout std_logic := 'Z';
          ELK18_DAT_N      : inout std_logic := 'Z';
          ELK_OUT_R        : in    std_logic;
          ELK_OUT_F        : in    std_logic;
          CCC_160M_FXD     : in    std_logic;
          CCC_160M_ADJ     : in    std_logic;
          ELK_IN_DDR_R     : out   std_logic;
          ELK_IN_DDR_F     : out   std_logic
        );

end DDR_BIDIR_LVDS_DUAL_CLK_18;

architecture DEF_ARCH of DDR_BIDIR_LVDS_DUAL_CLK_18 is 

  component DDR_REG
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          QR  : out   std_logic;
          QF  : out   std_logic
        );
  end component;

  component DDR_OUT
    port( DR  : in    std_logic := 'U';
          DF  : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component BIBUF_LVDS
    port( PADP : inout   std_logic;
          PADN : inout   std_logic;
          D    : in    std_logic := 'U';
          E    : in    std_logic := 'U';
          Y    : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal DDR_BIDIR_LVDS_DUAL_CLK_18_GND, BIBUF_LVDS_0_Y, 
        DDR_OUT_0_Q, \VCC\ : std_logic;

begin 


    DDR_REG_0 : DDR_REG
      port map(D => BIBUF_LVDS_0_Y, CLK => CCC_160M_ADJ, CLR => 
        DDR_BIDIR_LVDS_DUAL_CLK_18_GND, QR => ELK_IN_DDR_R, QF
         => ELK_IN_DDR_F);
    
    DDR_OUT_0 : DDR_OUT
      port map(DR => ELK_OUT_R, DF => ELK_OUT_F, CLK => 
        CCC_160M_FXD, CLR => DDR_BIDIR_LVDS_DUAL_CLK_18_GND, Q
         => DDR_OUT_0_Q);
    
    BIBUF_LVDS_0 : BIBUF_LVDS
      port map(PADP => ELK18_DAT_P, PADN => ELK18_DAT_N, D => 
        DDR_OUT_0_Q, E => DCB_SALT_SEL_c_i, Y => BIBUF_LVDS_0_Y);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    GND_i : GND
      port map(Y => DDR_BIDIR_LVDS_DUAL_CLK_18_GND);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SYNC_DAT_SEL_18 is

    port( ELK_TX_DAT                 : out   std_logic_vector(7 downto 0);
          PATT_ELK_DAT_18            : in    std_logic_vector(7 downto 0);
          OP_MODE_c_2_0              : in    std_logic;
          OP_MODE_c_1_0              : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_13 : in    std_logic;
          CLK_40M_GL                 : in    std_logic
        );

end SYNC_DAT_SEL_18;

architecture DEF_ARCH of SYNC_DAT_SEL_18 is 

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \N_SERDAT[0]\, \N_SERDAT[1]\, \N_SERDAT[2]\, 
        \N_SERDAT[3]\, \N_SERDAT[4]\, \N_SERDAT[5]\, 
        \N_SERDAT[6]\, \N_SERDAT[7]\, \GND\, \VCC\ : std_logic;

begin 


    \SERDAT_RNO[4]\ : NOR2A
      port map(A => PATT_ELK_DAT_18(4), B => OP_MODE_c_2_0, Y => 
        \N_SERDAT[4]\);
    
    \SERDAT_RNO[0]\ : NOR2A
      port map(A => PATT_ELK_DAT_18(0), B => OP_MODE_c_1_0, Y => 
        \N_SERDAT[0]\);
    
    \SERDAT[6]\ : DFN1C0
      port map(D => \N_SERDAT[6]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_13, Q => ELK_TX_DAT(6));
    
    \SERDAT[4]\ : DFN1C0
      port map(D => \N_SERDAT[4]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_13, Q => ELK_TX_DAT(4));
    
    \SERDAT_RNO[7]\ : OR2
      port map(A => PATT_ELK_DAT_18(7), B => OP_MODE_c_2_0, Y => 
        \N_SERDAT[7]\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \SERDAT_RNO[3]\ : OR2
      port map(A => PATT_ELK_DAT_18(3), B => OP_MODE_c_1_0, Y => 
        \N_SERDAT[3]\);
    
    \SERDAT_RNO[2]\ : OR2
      port map(A => PATT_ELK_DAT_18(2), B => OP_MODE_c_1_0, Y => 
        \N_SERDAT[2]\);
    
    \SERDAT[5]\ : DFN1C0
      port map(D => \N_SERDAT[5]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_13, Q => ELK_TX_DAT(5));
    
    \SERDAT[7]\ : DFN1C0
      port map(D => \N_SERDAT[7]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_13, Q => ELK_TX_DAT(7));
    
    GND_i : GND
      port map(Y => \GND\);
    
    \SERDAT_RNO[5]\ : NOR2A
      port map(A => PATT_ELK_DAT_18(5), B => OP_MODE_c_2_0, Y => 
        \N_SERDAT[5]\);
    
    \SERDAT[0]\ : DFN1C0
      port map(D => \N_SERDAT[0]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_13, Q => ELK_TX_DAT(0));
    
    \SERDAT_RNO[6]\ : NOR2A
      port map(A => PATT_ELK_DAT_18(6), B => OP_MODE_c_2_0, Y => 
        \N_SERDAT[6]\);
    
    \SERDAT[1]\ : DFN1C0
      port map(D => \N_SERDAT[1]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_13, Q => ELK_TX_DAT(1));
    
    \SERDAT_RNO[1]\ : OR2
      port map(A => PATT_ELK_DAT_18(1), B => OP_MODE_c_1_0, Y => 
        \N_SERDAT[1]\);
    
    \SERDAT[3]\ : DFN1C0
      port map(D => \N_SERDAT[3]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_13, Q => ELK_TX_DAT(3));
    
    \SERDAT[2]\ : DFN1C0
      port map(D => \N_SERDAT[2]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_13, Q => ELK_TX_DAT(2));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity ELINK_SLAVE_15_13 is

    port( BIT_OS_SEL_0               : in    std_logic_vector(2 downto 1);
          BIT_OS_SEL_1               : in    std_logic_vector(2 downto 1);
          BIT_OS_SEL_2               : in    std_logic_vector(1 downto 0);
          ELK_RX_SER_WORD_18         : out   std_logic_vector(7 downto 0);
          OP_MODE_c_1_0              : in    std_logic;
          OP_MODE_c_2_0              : in    std_logic;
          PATT_ELK_DAT_18            : in    std_logic_vector(7 downto 0);
          MASTER_DCB_POR_B_i_0_i     : in    std_logic;
          ELK18_DAT_N                : inout std_logic := 'Z';
          ELK18_DAT_P                : inout std_logic := 'Z';
          DCB_SALT_SEL_c_i           : in    std_logic;
          CCC_160M_FXD               : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_9  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_4  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_1  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_17 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_3  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_0  : in    std_logic;
          CLK_40M_GL                 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_13 : in    std_logic;
          DEV_RST_B_c_0              : in    std_logic;
          CCC_160M_ADJ               : in    std_logic
        );

end ELINK_SLAVE_15_13;

architecture DEF_ARCH of ELINK_SLAVE_15_13 is 

  component SLAVE_DES320S_1_17_16
    port( ELK_RX_SER_WORD_18     : out   std_logic_vector(7 downto 0);
          BIT_OS_SEL_2           : in    std_logic_vector(1 downto 0) := (others => 'U');
          BIT_OS_SEL_1           : in    std_logic_vector(2 downto 1) := (others => 'U');
          BIT_OS_SEL_0           : in    std_logic_vector(2 downto 1) := (others => 'U');
          CLK_40M_GL             : in    std_logic := 'U';
          CCC_160M_FXD           : in    std_logic := 'U';
          ELK_IN_R               : in    std_logic := 'U';
          ELK_IN_F               : in    std_logic := 'U';
          MASTER_DCB_POR_B_i_0_i : in    std_logic := 'U';
          CCC_160M_ADJ           : in    std_logic := 'U'
        );
  end component;

  component SER320M_3_34_18
    port( ELK_TX_DAT                 : in    std_logic_vector(7 downto 0) := (others => 'U');
          MASTER_SALT_POR_B_i_0_i_0  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_3  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_17 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_1  : in    std_logic := 'U';
          ELK_OUT_R                  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_4  : in    std_logic := 'U';
          ELK_OUT_F                  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_9  : in    std_logic := 'U';
          CCC_160M_FXD               : in    std_logic := 'U';
          CLK_40M_GL                 : in    std_logic := 'U'
        );
  end component;

  component DDR_BIDIR_LVDS_DUAL_CLK_18
    port( DCB_SALT_SEL_c_i : in    std_logic := 'U';
          ELK18_DAT_P      : inout   std_logic;
          ELK18_DAT_N      : inout   std_logic;
          ELK_OUT_R        : in    std_logic := 'U';
          ELK_OUT_F        : in    std_logic := 'U';
          CCC_160M_FXD     : in    std_logic := 'U';
          CCC_160M_ADJ     : in    std_logic := 'U';
          ELK_IN_DDR_R     : out   std_logic;
          ELK_IN_DDR_F     : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component SYNC_DAT_SEL_18
    port( ELK_TX_DAT                 : out   std_logic_vector(7 downto 0);
          PATT_ELK_DAT_18            : in    std_logic_vector(7 downto 0) := (others => 'U');
          OP_MODE_c_2_0              : in    std_logic := 'U';
          OP_MODE_c_1_0              : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_13 : in    std_logic := 'U';
          CLK_40M_GL                 : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \ELK_IN_F\, ELK_IN_DDR_F, \ELK_IN_R\, ELK_IN_DDR_R, 
        \ELK_TX_DAT[0]\, \ELK_TX_DAT[1]\, \ELK_TX_DAT[2]\, 
        \ELK_TX_DAT[3]\, \ELK_TX_DAT[4]\, \ELK_TX_DAT[5]\, 
        \ELK_TX_DAT[6]\, \ELK_TX_DAT[7]\, ELK_OUT_R, ELK_OUT_F, 
        \GND\, \VCC\ : std_logic;

    for all : SLAVE_DES320S_1_17_16
	Use entity work.SLAVE_DES320S_1_17_16(DEF_ARCH);
    for all : SER320M_3_34_18
	Use entity work.SER320M_3_34_18(DEF_ARCH);
    for all : DDR_BIDIR_LVDS_DUAL_CLK_18
	Use entity work.DDR_BIDIR_LVDS_DUAL_CLK_18(DEF_ARCH);
    for all : SYNC_DAT_SEL_18
	Use entity work.SYNC_DAT_SEL_18(DEF_ARCH);
begin 


    U_SLAVE_1ELK : SLAVE_DES320S_1_17_16
      port map(ELK_RX_SER_WORD_18(7) => ELK_RX_SER_WORD_18(7), 
        ELK_RX_SER_WORD_18(6) => ELK_RX_SER_WORD_18(6), 
        ELK_RX_SER_WORD_18(5) => ELK_RX_SER_WORD_18(5), 
        ELK_RX_SER_WORD_18(4) => ELK_RX_SER_WORD_18(4), 
        ELK_RX_SER_WORD_18(3) => ELK_RX_SER_WORD_18(3), 
        ELK_RX_SER_WORD_18(2) => ELK_RX_SER_WORD_18(2), 
        ELK_RX_SER_WORD_18(1) => ELK_RX_SER_WORD_18(1), 
        ELK_RX_SER_WORD_18(0) => ELK_RX_SER_WORD_18(0), 
        BIT_OS_SEL_2(1) => BIT_OS_SEL_2(1), BIT_OS_SEL_2(0) => 
        BIT_OS_SEL_2(0), BIT_OS_SEL_1(2) => BIT_OS_SEL_1(2), 
        BIT_OS_SEL_1(1) => BIT_OS_SEL_1(1), BIT_OS_SEL_0(2) => 
        BIT_OS_SEL_0(2), BIT_OS_SEL_0(1) => BIT_OS_SEL_0(1), 
        CLK_40M_GL => CLK_40M_GL, CCC_160M_FXD => CCC_160M_FXD, 
        ELK_IN_R => \ELK_IN_R\, ELK_IN_F => \ELK_IN_F\, 
        MASTER_DCB_POR_B_i_0_i => MASTER_DCB_POR_B_i_0_i, 
        CCC_160M_ADJ => CCC_160M_ADJ);
    
    U_ELK1_CMD_TX : SER320M_3_34_18
      port map(ELK_TX_DAT(7) => \ELK_TX_DAT[7]\, ELK_TX_DAT(6)
         => \ELK_TX_DAT[6]\, ELK_TX_DAT(5) => \ELK_TX_DAT[5]\, 
        ELK_TX_DAT(4) => \ELK_TX_DAT[4]\, ELK_TX_DAT(3) => 
        \ELK_TX_DAT[3]\, ELK_TX_DAT(2) => \ELK_TX_DAT[2]\, 
        ELK_TX_DAT(1) => \ELK_TX_DAT[1]\, ELK_TX_DAT(0) => 
        \ELK_TX_DAT[0]\, MASTER_SALT_POR_B_i_0_i_0 => 
        MASTER_SALT_POR_B_i_0_i_0, MASTER_SALT_POR_B_i_0_i_3 => 
        MASTER_SALT_POR_B_i_0_i_3, MASTER_SALT_POR_B_i_0_i_17 => 
        MASTER_SALT_POR_B_i_0_i_17, MASTER_SALT_POR_B_i_0_i_1 => 
        MASTER_SALT_POR_B_i_0_i_1, ELK_OUT_R => ELK_OUT_R, 
        MASTER_SALT_POR_B_i_0_i_4 => MASTER_SALT_POR_B_i_0_i_4, 
        ELK_OUT_F => ELK_OUT_F, MASTER_SALT_POR_B_i_0_i_9 => 
        MASTER_SALT_POR_B_i_0_i_9, CCC_160M_FXD => CCC_160M_FXD, 
        CLK_40M_GL => CLK_40M_GL);
    
    U_DDR_ELK1 : DDR_BIDIR_LVDS_DUAL_CLK_18
      port map(DCB_SALT_SEL_c_i => DCB_SALT_SEL_c_i, ELK18_DAT_P
         => ELK18_DAT_P, ELK18_DAT_N => ELK18_DAT_N, ELK_OUT_R
         => ELK_OUT_R, ELK_OUT_F => ELK_OUT_F, CCC_160M_FXD => 
        CCC_160M_FXD, CCC_160M_ADJ => CCC_160M_ADJ, ELK_IN_DDR_R
         => ELK_IN_DDR_R, ELK_IN_DDR_F => ELK_IN_DDR_F);
    
    ELK_IN_F : DFN1C0
      port map(D => ELK_IN_DDR_F, CLK => CCC_160M_ADJ, CLR => 
        DEV_RST_B_c_0, Q => \ELK_IN_F\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    U_ELK1_SERDAT_SOURCE : SYNC_DAT_SEL_18
      port map(ELK_TX_DAT(7) => \ELK_TX_DAT[7]\, ELK_TX_DAT(6)
         => \ELK_TX_DAT[6]\, ELK_TX_DAT(5) => \ELK_TX_DAT[5]\, 
        ELK_TX_DAT(4) => \ELK_TX_DAT[4]\, ELK_TX_DAT(3) => 
        \ELK_TX_DAT[3]\, ELK_TX_DAT(2) => \ELK_TX_DAT[2]\, 
        ELK_TX_DAT(1) => \ELK_TX_DAT[1]\, ELK_TX_DAT(0) => 
        \ELK_TX_DAT[0]\, PATT_ELK_DAT_18(7) => PATT_ELK_DAT_18(7), 
        PATT_ELK_DAT_18(6) => PATT_ELK_DAT_18(6), 
        PATT_ELK_DAT_18(5) => PATT_ELK_DAT_18(5), 
        PATT_ELK_DAT_18(4) => PATT_ELK_DAT_18(4), 
        PATT_ELK_DAT_18(3) => PATT_ELK_DAT_18(3), 
        PATT_ELK_DAT_18(2) => PATT_ELK_DAT_18(2), 
        PATT_ELK_DAT_18(1) => PATT_ELK_DAT_18(1), 
        PATT_ELK_DAT_18(0) => PATT_ELK_DAT_18(0), OP_MODE_c_2_0
         => OP_MODE_c_2_0, OP_MODE_c_1_0 => OP_MODE_c_1_0, 
        MASTER_SALT_POR_B_i_0_i_13 => MASTER_SALT_POR_B_i_0_i_13, 
        CLK_40M_GL => CLK_40M_GL);
    
    ELK_IN_R : DFN1C0
      port map(D => ELK_IN_DDR_R, CLK => CCC_160M_ADJ, CLR => 
        DEV_RST_B_c_0, Q => \ELK_IN_R\);
    
    GND_i : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity tristate_buf_1 is

    port( P_USB_MASTER_EN_c : in    std_logic;
          USB_OE_BI         : in    std_logic;
          USB_OE_B          : out   std_logic
        );

end tristate_buf_1;

architecture DEF_ARCH of tristate_buf_1 is 

  component TRIBUFF_F_24U
    port( D   : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          PAD : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \GND\, \VCC\ : std_logic;

begin 


    \TRIBUFF_F_24U[0]\ : TRIBUFF_F_24U
      port map(D => USB_OE_BI, E => P_USB_MASTER_EN_c, PAD => 
        USB_OE_B);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    GND_i : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity BIDIR_LVDS_IO_0 is

    port( DCB_SALT_SEL_c : in    std_logic;
          CLK_40M_GL     : in    std_logic;
          EXTCLK_40MHZ_c : out   std_logic;
          REF_CLK_0P     : inout std_logic := 'Z';
          REF_CLK_0N     : inout std_logic := 'Z'
        );

end BIDIR_LVDS_IO_0;

architecture DEF_ARCH of BIDIR_LVDS_IO_0 is 

  component BIBUF_LVDS
    port( PADP : inout   std_logic;
          PADN : inout   std_logic;
          D    : in    std_logic := 'U';
          E    : in    std_logic := 'U';
          Y    : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \GND\, \VCC\ : std_logic;

begin 


    \BIBUF_LVDS[0]\ : BIBUF_LVDS
      port map(PADP => REF_CLK_0P, PADN => REF_CLK_0N, D => 
        CLK_40M_GL, E => DCB_SALT_SEL_c, Y => EXTCLK_40MHZ_c);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    GND_i : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SLAVE_DES320S_1_17_9 is

    port( ELK_RX_SER_WORD_11     : out   std_logic_vector(7 downto 0);
          BIT_OS_SEL_0           : in    std_logic;
          BIT_OS_SEL_6_0         : in    std_logic;
          BIT_OS_SEL_7_0         : in    std_logic;
          BIT_OS_SEL_5           : in    std_logic_vector(2 downto 1);
          BIT_OS_SEL_4           : in    std_logic_vector(2 downto 1);
          CLK_40M_GL             : in    std_logic;
          CCC_160M_FXD           : in    std_logic;
          ELK_IN_R               : in    std_logic;
          ELK_IN_F               : in    std_logic;
          MASTER_DCB_POR_B_i_0_i : in    std_logic;
          CCC_160M_ADJ           : in    std_logic
        );

end SLAVE_DES320S_1_17_9;

architecture DEF_ARCH of SLAVE_DES320S_1_17_9 is 

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal N_17, \ARB_BYTE[0]_net_1\, \ARB_BYTE[4]_net_1\, N_18, 
        \ARB_BYTE[1]_net_1\, \ARB_BYTE[5]_net_1\, N_19, 
        \ARB_BYTE[2]_net_1\, \ARB_BYTE[6]_net_1\, N_20, 
        \ARB_BYTE[3]_net_1\, \ARB_BYTE[7]_net_1\, N_21, 
        \ARB_BYTE[8]_net_1\, N_22, \ARB_BYTE[9]_net_1\, N_23, 
        \ARB_BYTE[10]_net_1\, N_24, \ARB_BYTE[11]_net_1\, N_31, 
        \ARB_BYTE[12]_net_1\, N_32, \ARB_BYTE[13]_net_1\, N_33, 
        N_34, N_35, N_36, N_37, N_38, N_39, N_40, N_56, 
        \ARB_BYTE[14]_net_1\, N_64, \N_RECD_SER_WORD[0]\, 
        \N_RECD_SER_WORD[1]\, \N_RECD_SER_WORD[2]\, 
        \N_RECD_SER_WORD[3]\, \N_RECD_SER_WORD[4]\, 
        \N_RECD_SER_WORD[5]\, \N_RECD_SER_WORD[6]\, 
        \N_RECD_SER_WORD[7]\, \ADJ_SER_IN_F_0DEL\, 
        \ADJ_SER_IN_R_0DEL\, \ADJ_SER_IN_F_1DEL\, 
        \ADJ_SER_IN_R_1DEL\, \Q[0]_net_1\, \ADJ_Q[0]_net_1\, 
        \Q[1]_net_1\, \ADJ_Q[1]_net_1\, \Q[2]_net_1\, 
        \ADJ_Q[2]_net_1\, \Q[3]_net_1\, \ADJ_Q[3]_net_1\, 
        \Q[4]_net_1\, \ADJ_Q[4]_net_1\, \Q[5]_net_1\, 
        \ADJ_Q[5]_net_1\, \Q[6]_net_1\, \ADJ_Q[6]_net_1\, 
        \Q[7]_net_1\, \ADJ_Q[7]_net_1\, \Q[8]_net_1\, 
        \ADJ_Q[8]_net_1\, \Q[9]_net_1\, \ADJ_Q[9]_net_1\, 
        \Q[10]_net_1\, \ADJ_Q[10]_net_1\, \Q[11]_net_1\, 
        \ADJ_Q[11]_net_1\, \Q[12]_net_1\, \ADJ_Q[12]_net_1\, 
        \Q[13]_net_1\, \ADJ_Q[13]_net_1\, \Q[14]_net_1\, 
        \ADJ_Q[14]_net_1\, \ARB_WRD_40M_FIXED[0]_net_1\, 
        \ARB_WRD_40M_FIXED[1]_net_1\, 
        \ARB_WRD_40M_FIXED[2]_net_1\, 
        \ARB_WRD_40M_FIXED[3]_net_1\, 
        \ARB_WRD_40M_FIXED[4]_net_1\, 
        \ARB_WRD_40M_FIXED[5]_net_1\, 
        \ARB_WRD_40M_FIXED[6]_net_1\, 
        \ARB_WRD_40M_FIXED[7]_net_1\, 
        \ARB_WRD_40M_FIXED[8]_net_1\, 
        \ARB_WRD_40M_FIXED[9]_net_1\, 
        \ARB_WRD_40M_FIXED[10]_net_1\, 
        \ARB_WRD_40M_FIXED[11]_net_1\, 
        \ARB_WRD_40M_FIXED[12]_net_1\, 
        \ARB_WRD_40M_FIXED[13]_net_1\, 
        \ARB_WRD_40M_FIXED[14]_net_1\, \GND\, \VCC\ : std_logic;

begin 


    \RECD_SER_WORD_RNO[5]\ : MX2
      port map(A => N_38, B => N_39, S => BIT_OS_SEL_0, Y => 
        \N_RECD_SER_WORD[5]\);
    
    \ARB_WRD_40M_FIXED[9]\ : DFN1C0
      port map(D => \Q[9]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[9]_net_1\);
    
    \ADJ_Q[4]\ : DFN1C0
      port map(D => \ADJ_Q[2]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[4]_net_1\);
    
    \ARB_BYTE[6]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[6]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[6]_net_1\);
    
    ADJ_SER_IN_F_1DEL : DFN1C0
      port map(D => \ADJ_SER_IN_F_0DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_F_1DEL\);
    
    \ARB_BYTE[0]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[0]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[0]_net_1\);
    
    \ARB_BYTE_RNIBM701[1]\ : MX2
      port map(A => N_18, B => N_20, S => BIT_OS_SEL_4(1), Y => 
        N_34);
    
    \Q[11]\ : DFN1C0
      port map(D => \ADJ_Q[11]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[11]_net_1\);
    
    \ADJ_Q[8]\ : DFN1C0
      port map(D => \ADJ_Q[6]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[8]_net_1\);
    
    \ADJ_Q[6]\ : DFN1C0
      port map(D => \ADJ_Q[4]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[6]_net_1\);
    
    \ADJ_Q[12]\ : DFN1C0
      port map(D => \ADJ_Q[10]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[12]_net_1\);
    
    \RECD_SER_WORD_RNO_1[0]\ : MX2
      port map(A => \ARB_BYTE[0]_net_1\, B => \ARB_BYTE[4]_net_1\, 
        S => BIT_OS_SEL_4(2), Y => N_17);
    
    \ARB_BYTE_RNIJU701[3]\ : MX2
      port map(A => N_20, B => N_22, S => BIT_OS_SEL_4(1), Y => 
        N_36);
    
    \Q[1]\ : DFN1C0
      port map(D => \ADJ_Q[1]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[1]_net_1\);
    
    \ARB_BYTE[4]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[4]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[4]_net_1\);
    
    \ADJ_Q[2]\ : DFN1C0
      port map(D => \ADJ_Q[0]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[2]_net_1\);
    
    \RECD_SER_WORD_RNO_1[7]\ : MX2
      port map(A => \ARB_BYTE[10]_net_1\, B => 
        \ARB_BYTE[14]_net_1\, S => BIT_OS_SEL_7_0, Y => N_56);
    
    \RECD_SER_WORD[4]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[4]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_11(4));
    
    \Q[5]\ : DFN1C0
      port map(D => \ADJ_Q[5]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[5]_net_1\);
    
    \ADJ_Q[11]\ : DFN1C0
      port map(D => \ADJ_Q[9]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[11]_net_1\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \ADJ_Q[3]\ : DFN1C0
      port map(D => \ADJ_Q[1]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[3]_net_1\);
    
    \Q[10]\ : DFN1C0
      port map(D => \ADJ_Q[10]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[10]_net_1\);
    
    \ARB_WRD_40M_FIXED[6]\ : DFN1C0
      port map(D => \Q[6]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[6]_net_1\);
    
    \ARB_WRD_40M_FIXED[1]\ : DFN1C0
      port map(D => \Q[1]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[1]_net_1\);
    
    \RECD_SER_WORD[3]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[3]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_11(3));
    
    \RECD_SER_WORD[0]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[0]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_11(0));
    
    \RECD_SER_WORD_RNO[3]\ : MX2
      port map(A => N_36, B => N_37, S => BIT_OS_SEL_0, Y => 
        \N_RECD_SER_WORD[3]\);
    
    \Q[0]\ : DFN1C0
      port map(D => \ADJ_Q[0]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[0]_net_1\);
    
    \ARB_BYTE_RNISHQE[1]\ : MX2
      port map(A => \ARB_BYTE[1]_net_1\, B => \ARB_BYTE[5]_net_1\, 
        S => BIT_OS_SEL_4(2), Y => N_18);
    
    \RECD_SER_WORD_RNO_0[7]\ : MX2
      port map(A => N_31, B => N_56, S => BIT_OS_SEL_6_0, Y => 
        N_64);
    
    \Q[7]\ : DFN1C0
      port map(D => \ADJ_Q[7]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[7]_net_1\);
    
    \ARB_BYTE[14]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[14]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[14]_net_1\);
    
    \ARB_WRD_40M_FIXED[2]\ : DFN1C0
      port map(D => \Q[2]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[2]_net_1\);
    
    \ARB_WRD_40M_FIXED[14]\ : DFN1C0
      port map(D => \Q[14]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[14]_net_1\);
    
    \RECD_SER_WORD_RNO[2]\ : MX2
      port map(A => N_35, B => N_36, S => BIT_OS_SEL_0, Y => 
        \N_RECD_SER_WORD[2]\);
    
    \ARB_BYTE[2]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[2]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[2]_net_1\);
    
    \ADJ_Q[7]\ : DFN1C0
      port map(D => \ADJ_Q[5]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[7]_net_1\);
    
    \ARB_BYTE[8]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[8]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[8]_net_1\);
    
    \ARB_BYTE_RNIUJQE[2]\ : MX2
      port map(A => \ARB_BYTE[2]_net_1\, B => \ARB_BYTE[6]_net_1\, 
        S => BIT_OS_SEL_4(2), Y => N_19);
    
    \RECD_SER_WORD[5]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[5]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_11(5));
    
    \ARB_BYTE[12]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[12]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[12]_net_1\);
    
    \RECD_SER_WORD[1]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[1]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_11(1));
    
    \Q[3]\ : DFN1C0
      port map(D => \ADJ_Q[3]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[3]_net_1\);
    
    \ARB_BYTE_RNIFQ701[2]\ : MX2
      port map(A => N_19, B => N_21, S => BIT_OS_SEL_4(1), Y => 
        N_35);
    
    ADJ_SER_IN_F_0DEL : DFN1C0
      port map(D => ELK_IN_F, CLK => CCC_160M_ADJ, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_F_0DEL\);
    
    \RECD_SER_WORD_RNO[7]\ : MX2
      port map(A => N_40, B => N_64, S => BIT_OS_SEL_0, Y => 
        \N_RECD_SER_WORD[7]\);
    
    \RECD_SER_WORD_RNO[1]\ : MX2
      port map(A => N_34, B => N_35, S => BIT_OS_SEL_0, Y => 
        \N_RECD_SER_WORD[1]\);
    
    \ARB_WRD_40M_FIXED[4]\ : DFN1C0
      port map(D => \Q[4]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[4]_net_1\);
    
    \RECD_SER_WORD_RNO[0]\ : MX2
      port map(A => N_33, B => N_34, S => BIT_OS_SEL_0, Y => 
        \N_RECD_SER_WORD[0]\);
    
    \Q[6]\ : DFN1C0
      port map(D => \ADJ_Q[6]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[6]_net_1\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \ARB_WRD_40M_FIXED[8]\ : DFN1C0
      port map(D => \Q[8]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[8]_net_1\);
    
    \ARB_BYTE[11]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[11]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[11]_net_1\);
    
    \Q[9]\ : DFN1C0
      port map(D => \ADJ_Q[9]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[9]_net_1\);
    
    \ARB_BYTE_RNIFDOI[11]\ : MX2
      port map(A => \ARB_BYTE[7]_net_1\, B => 
        \ARB_BYTE[11]_net_1\, S => BIT_OS_SEL_4(2), Y => N_24);
    
    \Q[14]\ : DFN1C0
      port map(D => \ADJ_Q[14]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[14]_net_1\);
    
    \ARB_BYTE_RNIUH541[4]\ : MX2
      port map(A => N_21, B => N_23, S => BIT_OS_SEL_4(1), Y => 
        N_37);
    
    \ARB_BYTE_RNIKKRJ[13]\ : MX2
      port map(A => \ARB_BYTE[9]_net_1\, B => 
        \ARB_BYTE[13]_net_1\, S => BIT_OS_SEL_5(2), Y => N_32);
    
    ADJ_SER_IN_R_0DEL : DFN1C0
      port map(D => ELK_IN_R, CLK => CCC_160M_ADJ, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_R_0DEL\);
    
    \Q[13]\ : DFN1C0
      port map(D => \ADJ_Q[13]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[13]_net_1\);
    
    \ARB_BYTE[9]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[9]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[9]_net_1\);
    
    ADJ_SER_IN_R_1DEL : DFN1C0
      port map(D => \ADJ_SER_IN_R_0DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_R_1DEL\);
    
    \ARB_BYTE_RNI2OQE[4]\ : MX2
      port map(A => \ARB_BYTE[4]_net_1\, B => \ARB_BYTE[8]_net_1\, 
        S => BIT_OS_SEL_4(2), Y => N_21);
    
    \ARB_BYTE[10]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[10]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[10]_net_1\);
    
    \ADJ_Q[9]\ : DFN1C0
      port map(D => \ADJ_Q[7]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[9]_net_1\);
    
    \RECD_SER_WORD[7]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[7]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_11(7));
    
    \ARB_WRD_40M_FIXED[5]\ : DFN1C0
      port map(D => \Q[5]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[5]_net_1\);
    
    \ARB_WRD_40M_FIXED[12]\ : DFN1C0
      port map(D => \Q[12]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[12]_net_1\);
    
    \ARB_BYTE_RNIJJ9A1[13]\ : MX2
      port map(A => N_24, B => N_32, S => BIT_OS_SEL_5(1), Y => 
        N_40);
    
    \ARB_WRD_40M_FIXED[11]\ : DFN1C0
      port map(D => \Q[11]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[11]_net_1\);
    
    \ARB_WRD_40M_FIXED[0]\ : DFN1C0
      port map(D => \Q[0]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[0]_net_1\);
    
    \ARB_BYTE_RNIDBOI[6]\ : MX2
      port map(A => \ARB_BYTE[6]_net_1\, B => 
        \ARB_BYTE[10]_net_1\, S => BIT_OS_SEL_4(2), Y => N_23);
    
    \ADJ_Q[10]\ : DFN1C0
      port map(D => \ADJ_Q[8]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[10]_net_1\);
    
    \Q[2]\ : DFN1C0
      port map(D => \ADJ_Q[2]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[2]_net_1\);
    
    \ARB_BYTE_RNIIIRJ[12]\ : MX2
      port map(A => \ARB_BYTE[8]_net_1\, B => 
        \ARB_BYTE[12]_net_1\, S => BIT_OS_SEL_5(2), Y => N_31);
    
    \ARB_BYTE_RNI4QQE[5]\ : MX2
      port map(A => \ARB_BYTE[5]_net_1\, B => \ARB_BYTE[9]_net_1\, 
        S => BIT_OS_SEL_4(2), Y => N_22);
    
    \ARB_BYTE_RNI2M541[5]\ : MX2
      port map(A => N_22, B => N_24, S => BIT_OS_SEL_4(1), Y => 
        N_38);
    
    \ADJ_Q[1]\ : DFN1C0
      port map(D => \ADJ_SER_IN_F_1DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[1]_net_1\);
    
    \RECD_SER_WORD[6]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[6]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_11(6));
    
    \RECD_SER_WORD[2]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[2]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_11(2));
    
    \ADJ_Q[13]\ : DFN1C0
      port map(D => \ADJ_Q[11]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[13]_net_1\);
    
    \Q[8]\ : DFN1C0
      port map(D => \ADJ_Q[8]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[8]_net_1\);
    
    \ARB_BYTE[5]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[5]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[5]_net_1\);
    
    \ADJ_Q[14]\ : DFN1C0
      port map(D => \ADJ_Q[12]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[14]_net_1\);
    
    \RECD_SER_WORD_RNO[4]\ : MX2
      port map(A => N_37, B => N_38, S => BIT_OS_SEL_0, Y => 
        \N_RECD_SER_WORD[4]\);
    
    \Q[12]\ : DFN1C0
      port map(D => \ADJ_Q[12]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[12]_net_1\);
    
    \ARB_BYTE[13]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[13]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[13]_net_1\);
    
    \ARB_BYTE_RNIFF9A1[6]\ : MX2
      port map(A => N_23, B => N_31, S => BIT_OS_SEL_5(1), Y => 
        N_39);
    
    \ARB_WRD_40M_FIXED[3]\ : DFN1C0
      port map(D => \Q[3]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[3]_net_1\);
    
    \ARB_BYTE[7]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[7]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[7]_net_1\);
    
    \RECD_SER_WORD_RNO_0[0]\ : MX2
      port map(A => N_17, B => N_19, S => BIT_OS_SEL_4(1), Y => 
        N_33);
    
    \Q[4]\ : DFN1C0
      port map(D => \ADJ_Q[4]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[4]_net_1\);
    
    \ARB_WRD_40M_FIXED[7]\ : DFN1C0
      port map(D => \Q[7]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[7]_net_1\);
    
    \RECD_SER_WORD_RNO[6]\ : MX2
      port map(A => N_39, B => N_40, S => BIT_OS_SEL_0, Y => 
        \N_RECD_SER_WORD[6]\);
    
    \ARB_BYTE_RNI0MQE[3]\ : MX2
      port map(A => \ARB_BYTE[3]_net_1\, B => \ARB_BYTE[7]_net_1\, 
        S => BIT_OS_SEL_4(2), Y => N_20);
    
    \ARB_BYTE[3]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[3]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[3]_net_1\);
    
    \ADJ_Q[5]\ : DFN1C0
      port map(D => \ADJ_Q[3]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[5]_net_1\);
    
    \ARB_BYTE[1]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[1]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[1]_net_1\);
    
    \ARB_WRD_40M_FIXED[13]\ : DFN1C0
      port map(D => \Q[13]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[13]_net_1\);
    
    \ADJ_Q[0]\ : DFN1C0
      port map(D => \ADJ_SER_IN_R_1DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[0]_net_1\);
    
    \ARB_WRD_40M_FIXED[10]\ : DFN1C0
      port map(D => \Q[10]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[10]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SER320M_3_34_11 is

    port( ELK_TX_DAT                 : in    std_logic_vector(7 downto 0);
          MASTER_SALT_POR_B_i_0_i_7  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_11 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_2  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_10 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_16 : in    std_logic;
          ELK_OUT_R                  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_0  : in    std_logic;
          ELK_OUT_F                  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_5  : in    std_logic;
          CCC_160M_FXD               : in    std_logic;
          CLK_40M_GL                 : in    std_logic
        );

end SER320M_3_34_11;

architecture DEF_ARCH of SER320M_3_34_11 is 

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \N_SER_CMD_WORD_R[0]\, \START_RISE\, 
        \N_SER_CMD_WORD_F[0]\, \N_SER_CMD_WORD_R[3]\, 
        \SER_CMD_WORD_R[2]_net_1\, \N_SER_CMD_WORD_R[2]\, 
        \SER_CMD_WORD_R[1]_net_1\, \N_SER_CMD_WORD_R[1]\, 
        \SER_CMD_WORD_R[0]_net_1\, \N_SER_CMD_WORD_F[3]\, 
        \SER_CMD_WORD_F[2]_net_1\, \N_SER_CMD_WORD_F[2]\, 
        \SER_CMD_WORD_F[1]_net_1\, \N_SER_CMD_WORD_F[1]\, 
        \SER_CMD_WORD_F[0]_net_1\, N_START_RISE, 
        \CLK40M_GEN_DEL0\, \SER_OUT_FI\, \SER_OUT_RI\, 
        \SER_CMD_WORD_F[3]_net_1\, \SER_CMD_WORD_R[3]_net_1\, 
        \GND\, \VCC\ : std_logic;

begin 


    SER_OUT_FI : DFN1C0
      port map(D => \SER_CMD_WORD_F[3]_net_1\, CLK => 
        CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_2, Q => 
        \SER_OUT_FI\);
    
    \SER_CMD_WORD_F[3]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[3]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_11, Q => 
        \SER_CMD_WORD_F[3]_net_1\);
    
    \SER_CMD_WORD_R[1]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[1]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_7, Q => 
        \SER_CMD_WORD_R[1]_net_1\);
    
    \SER_CMD_WORD_R[2]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[2]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_7, Q => 
        \SER_CMD_WORD_R[2]_net_1\);
    
    \SER_CMD_WORD_R_RNO[3]\ : MX2
      port map(A => \SER_CMD_WORD_R[2]_net_1\, B => ELK_TX_DAT(7), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_R[3]\);
    
    \SER_CMD_WORD_R_RNO[0]\ : NOR2B
      port map(A => \START_RISE\, B => ELK_TX_DAT(1), Y => 
        \N_SER_CMD_WORD_R[0]\);
    
    \SER_CMD_WORD_F[0]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[0]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_11, Q => 
        \SER_CMD_WORD_F[0]_net_1\);
    
    \SER_CMD_WORD_R_RNO[1]\ : MX2
      port map(A => \SER_CMD_WORD_R[0]_net_1\, B => ELK_TX_DAT(3), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_R[1]\);
    
    \SER_CMD_WORD_F_RNO[2]\ : MX2
      port map(A => \SER_CMD_WORD_F[1]_net_1\, B => ELK_TX_DAT(4), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_F[2]\);
    
    \SER_CMD_WORD_F_RNO[3]\ : MX2
      port map(A => \SER_CMD_WORD_F[2]_net_1\, B => ELK_TX_DAT(6), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_F[3]\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    CLK40M_GEN_DEL0 : DFN1C0
      port map(D => CLK_40M_GL, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_5, Q => \CLK40M_GEN_DEL0\);
    
    SER_OUT_RI : DFN1C0
      port map(D => \SER_CMD_WORD_R[3]_net_1\, CLK => 
        CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_2, Q => 
        \SER_OUT_RI\);
    
    \SER_CMD_WORD_F[2]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[2]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_11, Q => 
        \SER_CMD_WORD_F[2]_net_1\);
    
    \SER_CMD_WORD_F_RNO[1]\ : MX2
      port map(A => \SER_CMD_WORD_F[0]_net_1\, B => ELK_TX_DAT(2), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_F[1]\);
    
    \SER_CMD_WORD_R[0]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[0]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_7, Q => 
        \SER_CMD_WORD_R[0]_net_1\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    START_RISE : DFN1C0
      port map(D => N_START_RISE, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_10, Q => \START_RISE\);
    
    \SER_CMD_WORD_R[3]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[3]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_7, Q => 
        \SER_CMD_WORD_R[3]_net_1\);
    
    \SER_CMD_WORD_F_RNO[0]\ : NOR2B
      port map(A => \START_RISE\, B => ELK_TX_DAT(0), Y => 
        \N_SER_CMD_WORD_F[0]\);
    
    SER_OUT_RDEL : DFN1C0
      port map(D => \SER_OUT_RI\, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_16, Q => ELK_OUT_R);
    
    \SER_CMD_WORD_F[1]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[1]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_11, Q => 
        \SER_CMD_WORD_F[1]_net_1\);
    
    START_RISE_RNO : NOR2B
      port map(A => \CLK40M_GEN_DEL0\, B => CLK_40M_GL, Y => 
        N_START_RISE);
    
    \SER_CMD_WORD_R_RNO[2]\ : MX2
      port map(A => \SER_CMD_WORD_R[1]_net_1\, B => ELK_TX_DAT(5), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_R[2]\);
    
    SER_OUT_FDEL : DFN1C0
      port map(D => \SER_OUT_FI\, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_0, Q => ELK_OUT_F);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity DDR_BIDIR_LVDS_DUAL_CLK_11 is

    port( DCB_SALT_SEL_c_i : in    std_logic;
          ELK11_DAT_P      : inout std_logic := 'Z';
          ELK11_DAT_N      : inout std_logic := 'Z';
          ELK_OUT_R        : in    std_logic;
          ELK_OUT_F        : in    std_logic;
          CCC_160M_FXD     : in    std_logic;
          CCC_160M_ADJ     : in    std_logic;
          ELK_IN_DDR_R     : out   std_logic;
          ELK_IN_DDR_F     : out   std_logic
        );

end DDR_BIDIR_LVDS_DUAL_CLK_11;

architecture DEF_ARCH of DDR_BIDIR_LVDS_DUAL_CLK_11 is 

  component DDR_REG
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          QR  : out   std_logic;
          QF  : out   std_logic
        );
  end component;

  component DDR_OUT
    port( DR  : in    std_logic := 'U';
          DF  : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component BIBUF_LVDS
    port( PADP : inout   std_logic;
          PADN : inout   std_logic;
          D    : in    std_logic := 'U';
          E    : in    std_logic := 'U';
          Y    : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal DDR_BIDIR_LVDS_DUAL_CLK_11_GND, BIBUF_LVDS_0_Y, 
        DDR_OUT_0_Q, \VCC\ : std_logic;

begin 


    DDR_REG_0 : DDR_REG
      port map(D => BIBUF_LVDS_0_Y, CLK => CCC_160M_ADJ, CLR => 
        DDR_BIDIR_LVDS_DUAL_CLK_11_GND, QR => ELK_IN_DDR_R, QF
         => ELK_IN_DDR_F);
    
    DDR_OUT_0 : DDR_OUT
      port map(DR => ELK_OUT_R, DF => ELK_OUT_F, CLK => 
        CCC_160M_FXD, CLR => DDR_BIDIR_LVDS_DUAL_CLK_11_GND, Q
         => DDR_OUT_0_Q);
    
    BIBUF_LVDS_0 : BIBUF_LVDS
      port map(PADP => ELK11_DAT_P, PADN => ELK11_DAT_N, D => 
        DDR_OUT_0_Q, E => DCB_SALT_SEL_c_i, Y => BIBUF_LVDS_0_Y);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    GND_i : GND
      port map(Y => DDR_BIDIR_LVDS_DUAL_CLK_11_GND);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SYNC_DAT_SEL_11 is

    port( ELK_TX_DAT                : out   std_logic_vector(7 downto 0);
          PATT_ELK_DAT_11           : in    std_logic_vector(7 downto 0);
          OP_MODE_c_0               : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_0 : in    std_logic;
          CLK_40M_GL                : in    std_logic
        );

end SYNC_DAT_SEL_11;

architecture DEF_ARCH of SYNC_DAT_SEL_11 is 

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \N_SERDAT[0]\, \N_SERDAT[1]\, \N_SERDAT[2]\, 
        \N_SERDAT[3]\, \N_SERDAT[4]\, \N_SERDAT[5]\, 
        \N_SERDAT[7]\, \N_SERDAT[6]\, \GND\, \VCC\ : std_logic;

begin 


    \SERDAT_RNO[4]\ : NOR2A
      port map(A => PATT_ELK_DAT_11(4), B => OP_MODE_c_0, Y => 
        \N_SERDAT[4]\);
    
    \SERDAT_RNO[0]\ : NOR2A
      port map(A => PATT_ELK_DAT_11(0), B => OP_MODE_c_0, Y => 
        \N_SERDAT[0]\);
    
    \SERDAT[6]\ : DFN1C0
      port map(D => \N_SERDAT[6]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_0, Q => ELK_TX_DAT(6));
    
    \SERDAT[4]\ : DFN1C0
      port map(D => \N_SERDAT[4]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_0, Q => ELK_TX_DAT(4));
    
    \SERDAT_RNO[7]\ : OR2
      port map(A => PATT_ELK_DAT_11(7), B => OP_MODE_c_0, Y => 
        \N_SERDAT[7]\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \SERDAT_RNO[3]\ : OR2
      port map(A => PATT_ELK_DAT_11(3), B => OP_MODE_c_0, Y => 
        \N_SERDAT[3]\);
    
    \SERDAT_RNO[2]\ : OR2
      port map(A => PATT_ELK_DAT_11(2), B => OP_MODE_c_0, Y => 
        \N_SERDAT[2]\);
    
    \SERDAT[5]\ : DFN1C0
      port map(D => \N_SERDAT[5]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_0, Q => ELK_TX_DAT(5));
    
    \SERDAT[7]\ : DFN1C0
      port map(D => \N_SERDAT[7]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_0, Q => ELK_TX_DAT(7));
    
    GND_i : GND
      port map(Y => \GND\);
    
    \SERDAT_RNO[5]\ : NOR2A
      port map(A => PATT_ELK_DAT_11(5), B => OP_MODE_c_0, Y => 
        \N_SERDAT[5]\);
    
    \SERDAT[0]\ : DFN1C0
      port map(D => \N_SERDAT[0]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_0, Q => ELK_TX_DAT(0));
    
    \SERDAT_RNO[6]\ : NOR2A
      port map(A => PATT_ELK_DAT_11(6), B => OP_MODE_c_0, Y => 
        \N_SERDAT[6]\);
    
    \SERDAT[1]\ : DFN1C0
      port map(D => \N_SERDAT[1]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_0, Q => ELK_TX_DAT(1));
    
    \SERDAT_RNO[1]\ : OR2
      port map(A => PATT_ELK_DAT_11(1), B => OP_MODE_c_0, Y => 
        \N_SERDAT[1]\);
    
    \SERDAT[3]\ : DFN1C0
      port map(D => \N_SERDAT[3]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_0, Q => ELK_TX_DAT(3));
    
    \SERDAT[2]\ : DFN1C0
      port map(D => \N_SERDAT[2]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_0, Q => ELK_TX_DAT(2));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity ELINK_SLAVE_15_6 is

    port( BIT_OS_SEL_4               : in    std_logic_vector(2 downto 1);
          BIT_OS_SEL_5               : in    std_logic_vector(2 downto 1);
          BIT_OS_SEL_7_0             : in    std_logic;
          BIT_OS_SEL_6_0             : in    std_logic;
          BIT_OS_SEL_0               : in    std_logic;
          ELK_RX_SER_WORD_11         : out   std_logic_vector(7 downto 0);
          OP_MODE_c_0                : in    std_logic;
          PATT_ELK_DAT_11            : in    std_logic_vector(7 downto 0);
          MASTER_DCB_POR_B_i_0_i     : in    std_logic;
          ELK11_DAT_N                : inout std_logic := 'Z';
          ELK11_DAT_P                : inout std_logic := 'Z';
          DCB_SALT_SEL_c_i           : in    std_logic;
          CCC_160M_FXD               : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_5  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_16 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_10 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_2  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_11 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_7  : in    std_logic;
          CLK_40M_GL                 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_0  : in    std_logic;
          DEV_RST_B_c_0              : in    std_logic;
          CCC_160M_ADJ               : in    std_logic
        );

end ELINK_SLAVE_15_6;

architecture DEF_ARCH of ELINK_SLAVE_15_6 is 

  component SLAVE_DES320S_1_17_9
    port( ELK_RX_SER_WORD_11     : out   std_logic_vector(7 downto 0);
          BIT_OS_SEL_0           : in    std_logic := 'U';
          BIT_OS_SEL_6_0         : in    std_logic := 'U';
          BIT_OS_SEL_7_0         : in    std_logic := 'U';
          BIT_OS_SEL_5           : in    std_logic_vector(2 downto 1) := (others => 'U');
          BIT_OS_SEL_4           : in    std_logic_vector(2 downto 1) := (others => 'U');
          CLK_40M_GL             : in    std_logic := 'U';
          CCC_160M_FXD           : in    std_logic := 'U';
          ELK_IN_R               : in    std_logic := 'U';
          ELK_IN_F               : in    std_logic := 'U';
          MASTER_DCB_POR_B_i_0_i : in    std_logic := 'U';
          CCC_160M_ADJ           : in    std_logic := 'U'
        );
  end component;

  component SER320M_3_34_11
    port( ELK_TX_DAT                 : in    std_logic_vector(7 downto 0) := (others => 'U');
          MASTER_SALT_POR_B_i_0_i_7  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_11 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_2  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_10 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_16 : in    std_logic := 'U';
          ELK_OUT_R                  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_0  : in    std_logic := 'U';
          ELK_OUT_F                  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_5  : in    std_logic := 'U';
          CCC_160M_FXD               : in    std_logic := 'U';
          CLK_40M_GL                 : in    std_logic := 'U'
        );
  end component;

  component DDR_BIDIR_LVDS_DUAL_CLK_11
    port( DCB_SALT_SEL_c_i : in    std_logic := 'U';
          ELK11_DAT_P      : inout   std_logic;
          ELK11_DAT_N      : inout   std_logic;
          ELK_OUT_R        : in    std_logic := 'U';
          ELK_OUT_F        : in    std_logic := 'U';
          CCC_160M_FXD     : in    std_logic := 'U';
          CCC_160M_ADJ     : in    std_logic := 'U';
          ELK_IN_DDR_R     : out   std_logic;
          ELK_IN_DDR_F     : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component SYNC_DAT_SEL_11
    port( ELK_TX_DAT                : out   std_logic_vector(7 downto 0);
          PATT_ELK_DAT_11           : in    std_logic_vector(7 downto 0) := (others => 'U');
          OP_MODE_c_0               : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_0 : in    std_logic := 'U';
          CLK_40M_GL                : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \ELK_IN_F\, ELK_IN_DDR_F, \ELK_IN_R\, ELK_IN_DDR_R, 
        \ELK_TX_DAT[0]\, \ELK_TX_DAT[1]\, \ELK_TX_DAT[2]\, 
        \ELK_TX_DAT[3]\, \ELK_TX_DAT[4]\, \ELK_TX_DAT[5]\, 
        \ELK_TX_DAT[6]\, \ELK_TX_DAT[7]\, ELK_OUT_R, ELK_OUT_F, 
        \GND\, \VCC\ : std_logic;

    for all : SLAVE_DES320S_1_17_9
	Use entity work.SLAVE_DES320S_1_17_9(DEF_ARCH);
    for all : SER320M_3_34_11
	Use entity work.SER320M_3_34_11(DEF_ARCH);
    for all : DDR_BIDIR_LVDS_DUAL_CLK_11
	Use entity work.DDR_BIDIR_LVDS_DUAL_CLK_11(DEF_ARCH);
    for all : SYNC_DAT_SEL_11
	Use entity work.SYNC_DAT_SEL_11(DEF_ARCH);
begin 


    U_SLAVE_1ELK : SLAVE_DES320S_1_17_9
      port map(ELK_RX_SER_WORD_11(7) => ELK_RX_SER_WORD_11(7), 
        ELK_RX_SER_WORD_11(6) => ELK_RX_SER_WORD_11(6), 
        ELK_RX_SER_WORD_11(5) => ELK_RX_SER_WORD_11(5), 
        ELK_RX_SER_WORD_11(4) => ELK_RX_SER_WORD_11(4), 
        ELK_RX_SER_WORD_11(3) => ELK_RX_SER_WORD_11(3), 
        ELK_RX_SER_WORD_11(2) => ELK_RX_SER_WORD_11(2), 
        ELK_RX_SER_WORD_11(1) => ELK_RX_SER_WORD_11(1), 
        ELK_RX_SER_WORD_11(0) => ELK_RX_SER_WORD_11(0), 
        BIT_OS_SEL_0 => BIT_OS_SEL_0, BIT_OS_SEL_6_0 => 
        BIT_OS_SEL_6_0, BIT_OS_SEL_7_0 => BIT_OS_SEL_7_0, 
        BIT_OS_SEL_5(2) => BIT_OS_SEL_5(2), BIT_OS_SEL_5(1) => 
        BIT_OS_SEL_5(1), BIT_OS_SEL_4(2) => BIT_OS_SEL_4(2), 
        BIT_OS_SEL_4(1) => BIT_OS_SEL_4(1), CLK_40M_GL => 
        CLK_40M_GL, CCC_160M_FXD => CCC_160M_FXD, ELK_IN_R => 
        \ELK_IN_R\, ELK_IN_F => \ELK_IN_F\, 
        MASTER_DCB_POR_B_i_0_i => MASTER_DCB_POR_B_i_0_i, 
        CCC_160M_ADJ => CCC_160M_ADJ);
    
    U_ELK1_CMD_TX : SER320M_3_34_11
      port map(ELK_TX_DAT(7) => \ELK_TX_DAT[7]\, ELK_TX_DAT(6)
         => \ELK_TX_DAT[6]\, ELK_TX_DAT(5) => \ELK_TX_DAT[5]\, 
        ELK_TX_DAT(4) => \ELK_TX_DAT[4]\, ELK_TX_DAT(3) => 
        \ELK_TX_DAT[3]\, ELK_TX_DAT(2) => \ELK_TX_DAT[2]\, 
        ELK_TX_DAT(1) => \ELK_TX_DAT[1]\, ELK_TX_DAT(0) => 
        \ELK_TX_DAT[0]\, MASTER_SALT_POR_B_i_0_i_7 => 
        MASTER_SALT_POR_B_i_0_i_7, MASTER_SALT_POR_B_i_0_i_11 => 
        MASTER_SALT_POR_B_i_0_i_11, MASTER_SALT_POR_B_i_0_i_2 => 
        MASTER_SALT_POR_B_i_0_i_2, MASTER_SALT_POR_B_i_0_i_10 => 
        MASTER_SALT_POR_B_i_0_i_10, MASTER_SALT_POR_B_i_0_i_16
         => MASTER_SALT_POR_B_i_0_i_16, ELK_OUT_R => ELK_OUT_R, 
        MASTER_SALT_POR_B_i_0_i_0 => MASTER_SALT_POR_B_i_0_i_0, 
        ELK_OUT_F => ELK_OUT_F, MASTER_SALT_POR_B_i_0_i_5 => 
        MASTER_SALT_POR_B_i_0_i_5, CCC_160M_FXD => CCC_160M_FXD, 
        CLK_40M_GL => CLK_40M_GL);
    
    U_DDR_ELK1 : DDR_BIDIR_LVDS_DUAL_CLK_11
      port map(DCB_SALT_SEL_c_i => DCB_SALT_SEL_c_i, ELK11_DAT_P
         => ELK11_DAT_P, ELK11_DAT_N => ELK11_DAT_N, ELK_OUT_R
         => ELK_OUT_R, ELK_OUT_F => ELK_OUT_F, CCC_160M_FXD => 
        CCC_160M_FXD, CCC_160M_ADJ => CCC_160M_ADJ, ELK_IN_DDR_R
         => ELK_IN_DDR_R, ELK_IN_DDR_F => ELK_IN_DDR_F);
    
    ELK_IN_F : DFN1C0
      port map(D => ELK_IN_DDR_F, CLK => CCC_160M_ADJ, CLR => 
        DEV_RST_B_c_0, Q => \ELK_IN_F\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    U_ELK1_SERDAT_SOURCE : SYNC_DAT_SEL_11
      port map(ELK_TX_DAT(7) => \ELK_TX_DAT[7]\, ELK_TX_DAT(6)
         => \ELK_TX_DAT[6]\, ELK_TX_DAT(5) => \ELK_TX_DAT[5]\, 
        ELK_TX_DAT(4) => \ELK_TX_DAT[4]\, ELK_TX_DAT(3) => 
        \ELK_TX_DAT[3]\, ELK_TX_DAT(2) => \ELK_TX_DAT[2]\, 
        ELK_TX_DAT(1) => \ELK_TX_DAT[1]\, ELK_TX_DAT(0) => 
        \ELK_TX_DAT[0]\, PATT_ELK_DAT_11(7) => PATT_ELK_DAT_11(7), 
        PATT_ELK_DAT_11(6) => PATT_ELK_DAT_11(6), 
        PATT_ELK_DAT_11(5) => PATT_ELK_DAT_11(5), 
        PATT_ELK_DAT_11(4) => PATT_ELK_DAT_11(4), 
        PATT_ELK_DAT_11(3) => PATT_ELK_DAT_11(3), 
        PATT_ELK_DAT_11(2) => PATT_ELK_DAT_11(2), 
        PATT_ELK_DAT_11(1) => PATT_ELK_DAT_11(1), 
        PATT_ELK_DAT_11(0) => PATT_ELK_DAT_11(0), OP_MODE_c_0 => 
        OP_MODE_c_0, MASTER_SALT_POR_B_i_0_i_0 => 
        MASTER_SALT_POR_B_i_0_i_0, CLK_40M_GL => CLK_40M_GL);
    
    ELK_IN_R : DFN1C0
      port map(D => ELK_IN_DDR_R, CLK => CCC_160M_ADJ, CLR => 
        DEV_RST_B_c_0, Q => \ELK_IN_R\);
    
    GND_i : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity GP_PATT_GEN_1_0 is

    port( ELKS_ADDRB            : out   std_logic_vector(7 downto 0);
          ELK_RX_SER_WORD_0     : in    std_logic_vector(7 downto 0);
          ELKS_STOP_ADDR        : in    std_logic_vector(7 downto 0);
          ELKS_STRT_ADDR        : in    std_logic_vector(7 downto 0);
          OP_MODE_0             : in    std_logic;
          OP_MODE_c_0           : in    std_logic;
          ELKS_ADDRB_0_0        : out   std_logic;
          ELKS_ADDRB_0_2        : out   std_logic;
          ELKS_ADDRB_0_4        : out   std_logic;
          P_MASTER_POR_B_c_32   : in    std_logic;
          P_MASTER_POR_B_c_26   : in    std_logic;
          P_MASTER_POR_B_c_25   : in    std_logic;
          P_MASTER_POR_B_c_23   : in    std_logic;
          P_MASTER_POR_B_c_7    : in    std_logic;
          P_MASTER_POR_B_c_11   : in    std_logic;
          P_MASTER_POR_B_c_29   : in    std_logic;
          DCB_SALT_SEL_c_i      : in    std_logic;
          P_MASTER_POR_B_c_2    : in    std_logic;
          P_MASTER_POR_B_c_12   : in    std_logic;
          ELKS_RWB              : out   std_logic;
          P_MASTER_POR_B_c_13   : in    std_logic;
          ELKS_RAM_BLKB_EN      : out   std_logic;
          P_USB_MASTER_EN_c     : in    std_logic;
          ALIGN_ACTIVE          : in    std_logic;
          P_MASTER_POR_B_c_34_0 : in    std_logic;
          P_MASTER_POR_B_c_32_0 : in    std_logic;
          P_MASTER_POR_B_c_31_0 : in    std_logic;
          CLK_40M_GL            : in    std_logic
        );

end GP_PATT_GEN_1_0;

architecture DEF_ARCH of GP_PATT_GEN_1_0 is 

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component DFN1E1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E0P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component INV
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XNOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component AOI1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component AO1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

    signal N_34, N_30, N_26, \GP_PG_SM_0[10]_net_1\, 
        \GP_PG_SM_ns[0]\, \DWACT_ADD_CI_0_g_array_11[0]\, 
        \DWACT_ADD_CI_0_g_array_2[0]\, 
        \DWACT_ADD_CI_0_pog_array_1_1[0]\, 
        \DWACT_ADD_CI_0_g_array_1[0]\, 
        \DWACT_ADD_CI_0_pog_array_1[0]\, \DWACT_ADD_CI_0_TMP[0]\, 
        \ELKS_ADDRB[1]\, \DWACT_ADD_CI_0_g_array_12_1[0]\, 
        \ELKS_ADDRB[4]\, \DWACT_ADD_CI_0_g_array_12_2[0]\, 
        \ELKS_ADDRB[6]\, \DWACT_ADD_CI_0_g_array_12[0]\, 
        \ELKS_ADDRB[2]\, \RX_SER_WORD_2DEL_i[1]\, 
        \RX_SER_WORD_2DEL[1]_net_1\, \RX_SER_WORD_2DEL_i[2]\, 
        \RX_SER_WORD_2DEL[2]_net_1\, \RX_SER_WORD_2DEL_i[3]\, 
        \RX_SER_WORD_2DEL[3]_net_1\, \RX_SER_WORD_2DEL_i[7]\, 
        \RX_SER_WORD_2DEL[7]_net_1\, \N_ADDR_POINTER_i_o2_0[7]\, 
        N_39, N_214_li, \GP_PG_SM[10]_net_1\, 
        \GP_PG_SM_ns_0_a2_0[5]\, \GP_PG_SM[5]_net_1\, 
        \GP_PG_SM[4]_net_1\, \GP_PG_SM_ns_i_i_a4_0[7]\, 
        \GP_PG_SM[3]_net_1\, \GP_PG_SM[2]_net_1\, 
        \GP_PG_SM_ns_i_i_a4_1[1]\, \GP_PG_SM[9]_net_1\, N_45, 
        \GP_PG_SM_ns_i_i_a4_0_1[7]\, \GP_PG_SM[8]_net_1\, N_114, 
        \GP_PG_SM_ns_i_i_a4_0[2]\, N_213_li, 
        \GP_PG_SM_ns_0_a4_2[0]\, N_315, \GP_PG_SM_ns_0_a4_0[0]\, 
        N_50, \GP_PG_SM[1]_net_1\, \GP_PG_SM_ns_0_a2_0_1[5]\, 
        \GP_PG_SM_ns_0_a4_0[6]\, \GP_PG_SM[6]_net_1\, 
        un1_RX_SER_WORD_2DEL_NE_4, \RX_SER_WORD_2DEL[5]_net_1\, 
        \RX_SER_WORD_2DEL[4]_net_1\, un1_RX_SER_WORD_2DEL_NE_1, 
        un1_RX_SER_WORD_2DEL_NE_3, un1_RX_SER_WORD_2DEL_NE_2, 
        \RX_SER_WORD_2DEL[0]_net_1\, \RX_SER_WORD_2DEL[6]_net_1\, 
        un1_RX_SER_WORD_3DEL_NE_4, \RX_SER_WORD_3DEL[5]_net_1\, 
        \RX_SER_WORD_3DEL[4]_net_1\, un1_RX_SER_WORD_3DEL_NE_1, 
        un1_RX_SER_WORD_3DEL_NE_3, \RX_SER_WORD_3DEL_i_0[2]\, 
        \RX_SER_WORD_3DEL_i_0[3]\, un1_RX_SER_WORD_3DEL_NE_2, 
        \RX_SER_WORD_3DEL[0]_net_1\, \RX_SER_WORD_3DEL_i_0[1]\, 
        \RX_SER_WORD_3DEL[6]_net_1\, \RX_SER_WORD_3DEL_i_0[7]\, 
        un1_RX_SER_WORD_3DEL_1, un1_RX_SER_WORD_2DEL_1, N_64, 
        N_22, N_210_li, \GP_PG_SM[7]_net_1\, N_116, N_80, N_69, 
        N_160_3, N_76, N_47, N_61, N_107, N_40, 
        \GP_PG_SM_RNO_0[1]_net_1\, N_73, N_42, N_24, N_83, N_85, 
        N_84, N_86, N_88, N_87, N_28, N_89, N_374, N_373, N_376, 
        N_377, N_375, N_32, N_379, N_380, N_378, N_382, N_383, 
        N_381, N_36, N_102, N_103, N_101, N_38, N_105, N_106, 
        N_104, N_18, N_117, \GP_PG_SM_ns_0_a2_0_1[3]\, 
        \GP_PG_SM_ns[3]\, \GP_PG_SM_ns_0_a2_0[3]\, N_25, N_238, 
        N_74, N_65, \GP_PG_SM_ns[10]\, \GP_PG_SM[0]_net_1\, 
        \GP_PG_SM_RNO_0[2]_net_1\, N_72, N_110, 
        \GP_PG_SM_RNO_0[3]_net_1\, \GP_PG_SM_ns[5]\, 
        \GP_PG_SM_ns[6]\, N_79, \LOC_STRT_ADDR[0]_net_1\, 
        \DWACT_ADD_CI_0_partial_sum[0]\, \LOC_STRT_ADDR[1]_net_1\, 
        I_30_0, \LOC_STRT_ADDR[2]_net_1\, I_29_0, 
        \LOC_STRT_ADDR[3]_net_1\, I_27_0, 
        \LOC_STRT_ADDR[4]_net_1\, I_33_0, 
        \LOC_STRT_ADDR[5]_net_1\, I_28_0, 
        \LOC_STRT_ADDR[6]_net_1\, I_31_0, 
        \LOC_STRT_ADDR[7]_net_1\, I_34_0, 
        \GP_PG_SM_RNIFMVG1[10]_net_1\, \LOC_STOP_ADDR[0]_net_1\, 
        \LOC_STOP_ADDR[1]_net_1\, \LOC_STOP_ADDR[2]_net_1\, 
        \LOC_STOP_ADDR[3]_net_1\, \LOC_STOP_ADDR[4]_net_1\, 
        \LOC_STOP_ADDR[5]_net_1\, \LOC_STOP_ADDR[6]_net_1\, 
        \LOC_STOP_ADDR[7]_net_1\, \RX_SER_WORD_1DEL[0]_net_1\, 
        \RX_SER_WORD_1DEL[1]_net_1\, \RX_SER_WORD_1DEL[2]_net_1\, 
        \RX_SER_WORD_1DEL[3]_net_1\, \RX_SER_WORD_1DEL[4]_net_1\, 
        \RX_SER_WORD_1DEL[5]_net_1\, \RX_SER_WORD_1DEL[6]_net_1\, 
        \RX_SER_WORD_1DEL[7]_net_1\, \ELKS_ADDRB[0]\, 
        \ELKS_ADDRB[3]\, \ELKS_ADDRB[5]\, \ELKS_ADDRB[7]\, 
        \DWACT_COMP0_E[1]\, \DWACT_COMP0_E[2]\, 
        \DWACT_COMP0_E[0]\, N_11, N_10, N_9, N_6, N_8, N_7, N_5, 
        N_2, N_3, N_4, \ACT_LT3_E[3]\, \ACT_LT3_E[4]\, 
        \ACT_LT3_E[5]\, \ACT_LT3_E[0]\, \ACT_LT3_E[1]\, 
        \ACT_LT3_E[2]\, \DWACT_BL_EQUAL_0_E[2]\, 
        \DWACT_BL_EQUAL_0_E[1]\, \DWACT_BL_EQUAL_0_E[0]\, \GND\, 
        \VCC\ : std_logic;

begin 

    ELKS_ADDRB(7) <= \ELKS_ADDRB[7]\;
    ELKS_ADDRB(6) <= \ELKS_ADDRB[6]\;
    ELKS_ADDRB(5) <= \ELKS_ADDRB[5]\;
    ELKS_ADDRB(4) <= \ELKS_ADDRB[4]\;
    ELKS_ADDRB(3) <= \ELKS_ADDRB[3]\;
    ELKS_ADDRB(2) <= \ELKS_ADDRB[2]\;
    ELKS_ADDRB(1) <= \ELKS_ADDRB[1]\;
    ELKS_ADDRB(0) <= \ELKS_ADDRB[0]\;

    \GP_PG_SM_RNIDKBH[6]\ : NOR2
      port map(A => \GP_PG_SM[6]_net_1\, B => \GP_PG_SM[7]_net_1\, 
        Y => N_114);
    
    \ADDR_POINTER_RNO_2[1]\ : OA1B
      port map(A => N_107, B => \N_ADDR_POINTER_i_o2_0[7]\, C => 
        ELKS_STRT_ADDR(1), Y => N_101);
    
    un1_ADDR_POINTER_2_I_46 : AND2
      port map(A => \ELKS_ADDRB[2]\, B => \ELKS_ADDRB[3]\, Y => 
        \DWACT_ADD_CI_0_pog_array_1[0]\);
    
    \GP_PG.un1_ADDR_POINTER_0_I_25\ : AO1
      port map(A => \DWACT_COMP0_E[1]\, B => \DWACT_COMP0_E[2]\, 
        C => \DWACT_COMP0_E[0]\, Y => N_214_li);
    
    \GP_PG_SM_RNO_0[8]\ : NOR2B
      port map(A => \GP_PG_SM[9]_net_1\, B => N_213_li, Y => 
        \GP_PG_SM_ns_i_i_a4_0[2]\);
    
    un1_ADDR_POINTER_2_I_45 : NOR2B
      port map(A => \DWACT_ADD_CI_0_g_array_1[0]\, B => 
        \ELKS_ADDRB[2]\, Y => \DWACT_ADD_CI_0_g_array_12[0]\);
    
    \GP_PG_SM_RNO_1[4]\ : NOR3C
      port map(A => N_214_li, B => N_117, C => 
        \GP_PG_SM[4]_net_1\, Y => N_79);
    
    \GP_PG_SM_RNIF42K1[1]\ : NOR2A
      port map(A => N_110, B => N_61, Y => N_116);
    
    \ADDR_POINTER_0[6]\ : DFN1C0
      port map(D => N_26, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_32_0, Q => ELKS_ADDRB_0_4);
    
    \ADDR_POINTER[2]\ : DFN1C0
      port map(D => N_34, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_31_0, Q => \ELKS_ADDRB[2]\);
    
    \RX_SER_WORD_1DEL[7]\ : DFN1C0
      port map(D => ELK_RX_SER_WORD_0(7), CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_23, Q => \RX_SER_WORD_1DEL[7]_net_1\);
    
    \GP_PG.un1_ADDR_POINTER_0_I_21\ : OR2A
      port map(A => \ELKS_ADDRB[4]\, B => 
        \LOC_STOP_ADDR[4]_net_1\, Y => N_9);
    
    \GP_PG_SM_RNO_2[2]\ : OR2B
      port map(A => N_47, B => \GP_PG_SM[2]_net_1\, Y => N_65);
    
    \RX_SER_WORD_3DEL[7]\ : DFN1P0
      port map(D => \RX_SER_WORD_2DEL_i[7]\, CLK => CLK_40M_GL, 
        PRE => P_MASTER_POR_B_c_31_0, Q => 
        \RX_SER_WORD_3DEL_i_0[7]\);
    
    \LOC_STOP_ADDR[2]\ : DFN1E1C0
      port map(D => ELKS_STOP_ADDR(2), CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_7, E => \GP_PG_SM_0[10]_net_1\, Q => 
        \LOC_STOP_ADDR[2]_net_1\);
    
    un1_ADDR_POINTER_2_I_28 : XOR2
      port map(A => \ELKS_ADDRB[5]\, B => 
        \DWACT_ADD_CI_0_g_array_12_1[0]\, Y => I_28_0);
    
    \ADDR_POINTER_RNO[5]\ : NOR3
      port map(A => N_89, B => N_374, C => N_373, Y => N_28);
    
    \LOC_STOP_ADDR[1]\ : DFN1E1C0
      port map(D => ELKS_STOP_ADDR(1), CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_7, E => \GP_PG_SM_0[10]_net_1\, Q => 
        \LOC_STOP_ADDR[1]_net_1\);
    
    \GP_PG_SM_RNO[8]\ : NOR3C
      port map(A => N_315, B => \GP_PG_SM_ns_i_i_a4_0[2]\, C => 
        N_116, Y => N_80);
    
    \GP_PG_SM_RNIL4A1K[10]\ : OA1B
      port map(A => N_107, B => \N_ADDR_POINTER_i_o2_0[7]\, C => 
        ELKS_STRT_ADDR(2), Y => N_381);
    
    \RX_SER_WORD_1DEL[0]\ : DFN1C0
      port map(D => ELK_RX_SER_WORD_0(0), CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_23, Q => \RX_SER_WORD_1DEL[0]_net_1\);
    
    \ADDR_POINTER_RNO_0[5]\ : OA1B
      port map(A => N_107, B => \N_ADDR_POINTER_i_o2_0[7]\, C => 
        ELKS_STRT_ADDR(5), Y => N_89);
    
    \RX_SER_WORD_3DEL[0]\ : DFN1C0
      port map(D => \RX_SER_WORD_2DEL[0]_net_1\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_31_0, Q => 
        \RX_SER_WORD_3DEL[0]_net_1\);
    
    \LOC_STRT_ADDR_RNIM80EA1[2]\ : NOR3
      port map(A => N_382, B => N_383, C => N_381, Y => N_34);
    
    un1_ADDR_POINTER_2_I_31 : XOR2
      port map(A => \ELKS_ADDRB[6]\, B => 
        \DWACT_ADD_CI_0_g_array_11[0]\, Y => I_31_0);
    
    \RX_SER_WORD_2DEL_RNISQ9J1[0]\ : OR3
      port map(A => un1_RX_SER_WORD_2DEL_NE_3, B => 
        un1_RX_SER_WORD_2DEL_NE_2, C => un1_RX_SER_WORD_2DEL_NE_4, 
        Y => un1_RX_SER_WORD_2DEL_1);
    
    \ADDR_POINTER_RNO[3]\ : NOR3
      port map(A => N_379, B => N_380, C => N_378, Y => N_32);
    
    \ADDR_POINTER[1]\ : DFN1C0
      port map(D => N_36, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_31_0, Q => \ELKS_ADDRB[1]\);
    
    \GP_PG_SM[0]\ : DFN1C0
      port map(D => \GP_PG_SM_ns[10]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_29, Q => \GP_PG_SM[0]_net_1\);
    
    \LOC_STRT_ADDR[5]\ : DFN1E1C0
      port map(D => ELKS_STRT_ADDR(5), CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_11, E => \GP_PG_SM_0[10]_net_1\, Q => 
        \LOC_STRT_ADDR[5]_net_1\);
    
    \LOC_STRT_ADDR_RNIVDV4B1[4]\ : NOR3
      port map(A => N_376, B => N_377, C => N_375, Y => N_30);
    
    \GP_PG_SM_RNIUFCB1[5]\ : NOR2A
      port map(A => N_117, B => N_40, Y => N_25);
    
    \ADDR_POINTER_RNO_2[7]\ : NOR3A
      port map(A => N_42, B => \GP_PG_SM[10]_net_1\, C => I_34_0, 
        Y => N_84);
    
    \GP_PG_SM_RNI3PVC[0]\ : NOR2A
      port map(A => \GP_PG_SM[0]_net_1\, B => OP_MODE_c_0, Y => 
        N_72);
    
    \ADDR_POINTER_RNO_1[0]\ : NOR3A
      port map(A => N_39, B => N_214_li, C => 
        \LOC_STRT_ADDR[0]_net_1\, Y => N_106);
    
    \GP_PG_SM_RNO_0[3]\ : NOR3C
      port map(A => OP_MODE_0, B => \GP_PG_SM[8]_net_1\, C => 
        N_114, Y => \GP_PG_SM_ns_i_i_a4_0_1[7]\);
    
    \GP_PG.un1_ADDR_POINTER_0_I_17\ : OR2A
      port map(A => \LOC_STOP_ADDR[4]_net_1\, B => 
        \ELKS_ADDRB[4]\, Y => N_5);
    
    \RX_SER_WORD_3DEL_RNINOOL[2]\ : OR2
      port map(A => \RX_SER_WORD_3DEL_i_0[2]\, B => 
        \RX_SER_WORD_3DEL_i_0[3]\, Y => un1_RX_SER_WORD_3DEL_NE_3);
    
    \ADDR_POINTER_RNO_2[0]\ : OA1B
      port map(A => N_107, B => \N_ADDR_POINTER_i_o2_0[7]\, C => 
        ELKS_STRT_ADDR(0), Y => N_104);
    
    R_BLKB : DFN1E0P0
      port map(D => N_160_3, CLK => CLK_40M_GL, PRE => 
        P_MASTER_POR_B_c_13, E => N_238, Q => ELKS_RAM_BLKB_EN);
    
    \LOC_STRT_ADDR[0]\ : DFN1E1C0
      port map(D => ELKS_STRT_ADDR(0), CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_11, E => \GP_PG_SM_0[10]_net_1\, Q => 
        \LOC_STRT_ADDR[0]_net_1\);
    
    \RX_SER_WORD_3DEL_RNIJKOL[0]\ : OR2
      port map(A => \RX_SER_WORD_3DEL[0]_net_1\, B => 
        \RX_SER_WORD_3DEL_i_0[1]\, Y => un1_RX_SER_WORD_3DEL_NE_2);
    
    \ADDR_POINTER_0[4]\ : DFN1C0
      port map(D => N_30, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_32_0, Q => ELKS_ADDRB_0_2);
    
    \GP_PG_SM_RNO[7]\ : OA1
      port map(A => \GP_PG_SM_ns_0_a2_0[3]\, B => 
        \GP_PG_SM_ns_0_a2_0_1[3]\, C => N_25, Y => 
        \GP_PG_SM_ns[3]\);
    
    \RX_SER_WORD_3DEL_RNO[2]\ : INV
      port map(A => \RX_SER_WORD_2DEL[2]_net_1\, Y => 
        \RX_SER_WORD_2DEL_i[2]\);
    
    \RX_SER_WORD_2DEL_RNIH8QC[0]\ : OR2A
      port map(A => \RX_SER_WORD_2DEL[1]_net_1\, B => 
        \RX_SER_WORD_2DEL[0]_net_1\, Y => 
        un1_RX_SER_WORD_2DEL_NE_2);
    
    \GP_PG_SM_RNO_1[5]\ : NOR3C
      port map(A => N_214_li, B => N_117, C => 
        \GP_PG_SM_ns_0_a2_0[5]\, Y => N_18);
    
    \RX_SER_WORD_1DEL[4]\ : DFN1C0
      port map(D => ELK_RX_SER_WORD_0(4), CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_23, Q => \RX_SER_WORD_1DEL[4]_net_1\);
    
    \ADDR_POINTER[6]\ : DFN1C0
      port map(D => N_26, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_32, Q => \ELKS_ADDRB[6]\);
    
    \GP_PG.un1_ADDR_POINTER_0_I_7\ : NOR2A
      port map(A => \LOC_STOP_ADDR[5]_net_1\, B => 
        \ELKS_ADDRB[5]\, Y => \ACT_LT3_E[0]\);
    
    \RX_SER_WORD_1DEL[2]\ : DFN1C0
      port map(D => ELK_RX_SER_WORD_0(2), CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_23, Q => \RX_SER_WORD_1DEL[2]_net_1\);
    
    \RX_SER_WORD_3DEL[4]\ : DFN1C0
      port map(D => \RX_SER_WORD_2DEL[4]_net_1\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_31_0, Q => 
        \RX_SER_WORD_3DEL[4]_net_1\);
    
    R_BLKB_RNO : OR3A
      port map(A => OP_MODE_c_0, B => \GP_PG_SM[1]_net_1\, C => 
        N_45, Y => N_160_3);
    
    \RX_SER_WORD_3DEL[2]\ : DFN1P0
      port map(D => \RX_SER_WORD_2DEL_i[2]\, CLK => CLK_40M_GL, 
        PRE => P_MASTER_POR_B_c_31_0, Q => 
        \RX_SER_WORD_3DEL_i_0[2]\);
    
    \GP_PG.un1_ADDR_POINTER_0_I_13\ : AOI1A
      port map(A => \ACT_LT3_E[3]\, B => \ACT_LT3_E[4]\, C => 
        \ACT_LT3_E[5]\, Y => \DWACT_COMP0_E[0]\);
    
    \GP_PG_SM_RNO[9]\ : NOR3C
      port map(A => \GP_PG_SM_ns_i_i_a4_1[1]\, B => N_315, C => 
        N_116, Y => N_69);
    
    \GP_PG.un1_ADDR_POINTER_0_I_1\ : XNOR2
      port map(A => \ELKS_ADDRB[7]\, B => 
        \LOC_STOP_ADDR[7]_net_1\, Y => \DWACT_BL_EQUAL_0_E[2]\);
    
    \ADDR_POINTER_RNO_0[7]\ : OA1B
      port map(A => N_107, B => \N_ADDR_POINTER_i_o2_0[7]\, C => 
        ELKS_STRT_ADDR(7), Y => N_83);
    
    \GP_PG_SM_RNIP8A1K[10]\ : OA1B
      port map(A => N_107, B => \N_ADDR_POINTER_i_o2_0[7]\, C => 
        ELKS_STRT_ADDR(6), Y => N_86);
    
    \GP_PG_SM_RNIO67Q9[5]\ : NOR3A
      port map(A => N_40, B => N_39, C => N_214_li, Y => N_107);
    
    \GP_PG.un1_ADDR_POINTER_0_I_4\ : AND3
      port map(A => \DWACT_BL_EQUAL_0_E[2]\, B => 
        \DWACT_BL_EQUAL_0_E[1]\, C => \DWACT_BL_EQUAL_0_E[0]\, Y
         => \DWACT_COMP0_E[1]\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    un1_ADDR_POINTER_2_I_34 : XOR2
      port map(A => \ELKS_ADDRB[7]\, B => 
        \DWACT_ADD_CI_0_g_array_12_2[0]\, Y => I_34_0);
    
    \GP_PG_SM_RNI18BH[1]\ : OR2
      port map(A => \GP_PG_SM[0]_net_1\, B => \GP_PG_SM[1]_net_1\, 
        Y => N_61);
    
    \GP_PG.un1_ADDR_POINTER_0_I_24\ : OA1
      port map(A => N_11, B => N_10, C => N_9, Y => 
        \DWACT_COMP0_E[2]\);
    
    un1_ADDR_POINTER_2_I_33 : XOR2
      port map(A => \ELKS_ADDRB[4]\, B => 
        \DWACT_ADD_CI_0_g_array_2[0]\, Y => I_33_0);
    
    \GP_PG_SM[6]\ : DFN1C0
      port map(D => N_22, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_29, Q => \GP_PG_SM[6]_net_1\);
    
    \GP_PG_SM_RNO_1[2]\ : AOI1B
      port map(A => \GP_PG_SM[6]_net_1\, B => OP_MODE_0, C => 
        N_65, Y => N_74);
    
    \LOC_STOP_ADDR[4]\ : DFN1E1C0
      port map(D => ELKS_STOP_ADDR(4), CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_7, E => \GP_PG_SM_0[10]_net_1\, Q => 
        \LOC_STOP_ADDR[4]_net_1\);
    
    \LOC_STOP_ADDR[5]\ : DFN1E1C0
      port map(D => ELKS_STOP_ADDR(5), CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_7, E => \GP_PG_SM_0[10]_net_1\, Q => 
        \LOC_STOP_ADDR[5]_net_1\);
    
    \ADDR_POINTER_RNO_0[0]\ : NOR3A
      port map(A => N_42, B => \GP_PG_SM[10]_net_1\, C => 
        \DWACT_ADD_CI_0_partial_sum[0]\, Y => N_105);
    
    un1_ADDR_POINTER_2_I_36 : NOR2B
      port map(A => \DWACT_ADD_CI_0_TMP[0]\, B => \ELKS_ADDRB[1]\, 
        Y => \DWACT_ADD_CI_0_g_array_1[0]\);
    
    \GP_PG.un1_ADDR_POINTER_0_I_12\ : AND2A
      port map(A => \LOC_STOP_ADDR[7]_net_1\, B => 
        \ELKS_ADDRB[7]\, Y => \ACT_LT3_E[5]\);
    
    un1_ADDR_POINTER_2_I_29 : XOR2
      port map(A => \ELKS_ADDRB[2]\, B => 
        \DWACT_ADD_CI_0_g_array_1[0]\, Y => I_29_0);
    
    \GP_PG_SM[5]\ : DFN1C0
      port map(D => \GP_PG_SM_ns[5]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_29, Q => \GP_PG_SM[5]_net_1\);
    
    un1_ADDR_POINTER_2_I_35 : NOR2B
      port map(A => \DWACT_ADD_CI_0_g_array_1[0]\, B => 
        \DWACT_ADD_CI_0_pog_array_1[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_2[0]\);
    
    \ADDR_POINTER[0]\ : DFN1C0
      port map(D => N_38, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_31_0, Q => \ELKS_ADDRB[0]\);
    
    \ADDR_POINTER_0[2]\ : DFN1C0
      port map(D => N_34, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_31_0, Q => ELKS_ADDRB_0_0);
    
    \GP_PG_SM_RNO_0[9]\ : NOR3A
      port map(A => OP_MODE_c_0, B => \GP_PG_SM[9]_net_1\, C => 
        N_45, Y => \GP_PG_SM_ns_i_i_a4_1[1]\);
    
    \RX_SER_WORD_2DEL_RNILCQC[2]\ : OR2B
      port map(A => \RX_SER_WORD_2DEL[2]_net_1\, B => 
        \RX_SER_WORD_2DEL[3]_net_1\, Y => 
        un1_RX_SER_WORD_2DEL_NE_3);
    
    \GP_PG_SM_RNO[2]\ : AOI1
      port map(A => N_64, B => \GP_PG_SM[0]_net_1\, C => N_74, Y
         => \GP_PG_SM_RNO_0[2]_net_1\);
    
    \LOC_STRT_ADDR_RNIT6OG9[6]\ : NOR3A
      port map(A => N_39, B => N_214_li, C => 
        \LOC_STRT_ADDR[6]_net_1\, Y => N_88);
    
    \ADDR_POINTER_RNO[0]\ : NOR3
      port map(A => N_105, B => N_106, C => N_104, Y => N_38);
    
    \RX_SER_WORD_3DEL_RNIV0PL[6]\ : OR2
      port map(A => \RX_SER_WORD_3DEL[6]_net_1\, B => 
        \RX_SER_WORD_3DEL_i_0[7]\, Y => un1_RX_SER_WORD_3DEL_NE_1);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \LOC_STRT_ADDR_RNIR4OG9[4]\ : NOR3A
      port map(A => N_39, B => N_214_li, C => 
        \LOC_STRT_ADDR[4]_net_1\, Y => N_377);
    
    \GP_PG_SM[7]\ : DFN1C0
      port map(D => \GP_PG_SM_ns[3]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_29, Q => \GP_PG_SM[7]_net_1\);
    
    \GP_PG_SM_RNIETPL[0]\ : AO1C
      port map(A => \GP_PG_SM[0]_net_1\, B => N_45, C => 
        OP_MODE_c_0, Y => N_50);
    
    \GP_PG_SM_RNO_2[5]\ : NOR2A
      port map(A => \GP_PG_SM[5]_net_1\, B => \GP_PG_SM[4]_net_1\, 
        Y => \GP_PG_SM_ns_0_a2_0[5]\);
    
    \GP_PG_SM[1]\ : DFN1C0
      port map(D => \GP_PG_SM_RNO_0[1]_net_1\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_29, Q => \GP_PG_SM[1]_net_1\);
    
    \GP_PG_SM_RNIM7S9E[10]\ : NOR3A
      port map(A => N_42, B => \GP_PG_SM[10]_net_1\, C => I_31_0, 
        Y => N_87);
    
    \GP_PG.un1_ADDR_POINTER_0_I_19\ : OA1A
      port map(A => \ELKS_ADDRB[3]\, B => 
        \LOC_STOP_ADDR[3]_net_1\, C => N_3, Y => N_7);
    
    un1_ADDR_POINTER_2_I_1 : AND2
      port map(A => \ELKS_ADDRB[0]\, B => 
        \GP_PG_SM_RNIFMVG1[10]_net_1\, Y => 
        \DWACT_ADD_CI_0_TMP[0]\);
    
    \GP_PG_SM_RNO_1[3]\ : NOR3B
      port map(A => \GP_PG_SM_ns_i_i_a4_0[7]\, B => N_47, C => 
        N_61, Y => N_76);
    
    \GP_PG_SM_RNO_2[3]\ : NOR2A
      port map(A => \GP_PG_SM[3]_net_1\, B => \GP_PG_SM[2]_net_1\, 
        Y => \GP_PG_SM_ns_i_i_a4_0[7]\);
    
    \GP_PG_SM_RNO[4]\ : AO1
      port map(A => \GP_PG_SM_ns_0_a4_0[6]\, B => N_117, C => 
        N_79, Y => \GP_PG_SM_ns[6]\);
    
    LOC_DIR_MODE : DFN1E1C0
      port map(D => DCB_SALT_SEL_c_i, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_2, E => \GP_PG_SM_0[10]_net_1\, Q => 
        N_213_li);
    
    \ADDR_POINTER_RNO_2[3]\ : OA1B
      port map(A => N_107, B => \N_ADDR_POINTER_i_o2_0[7]\, C => 
        ELKS_STRT_ADDR(3), Y => N_378);
    
    un1_ADDR_POINTER_2_I_27 : XOR2
      port map(A => \ELKS_ADDRB[3]\, B => 
        \DWACT_ADD_CI_0_g_array_12[0]\, Y => I_27_0);
    
    \ADDR_POINTER_RNO_1[7]\ : NOR3A
      port map(A => N_39, B => N_214_li, C => 
        \LOC_STRT_ADDR[7]_net_1\, Y => N_85);
    
    \RX_SER_WORD_3DEL_RNO[1]\ : INV
      port map(A => \RX_SER_WORD_2DEL[1]_net_1\, Y => 
        \RX_SER_WORD_2DEL_i[1]\);
    
    \GP_PG_SM[10]\ : DFN1P0
      port map(D => \GP_PG_SM_ns[0]\, CLK => CLK_40M_GL, PRE => 
        P_MASTER_POR_B_c_34_0, Q => \GP_PG_SM[10]_net_1\);
    
    un1_ADDR_POINTER_2_I_49 : AND2
      port map(A => \ELKS_ADDRB[4]\, B => \ELKS_ADDRB[5]\, Y => 
        \DWACT_ADD_CI_0_pog_array_1_1[0]\);
    
    \GP_PG_SM_RNIFMVG1[10]\ : OR2A
      port map(A => N_110, B => \GP_PG_SM[10]_net_1\, Y => 
        \GP_PG_SM_RNIFMVG1[10]_net_1\);
    
    \ADDR_POINTER[4]\ : DFN1C0
      port map(D => N_30, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_32, Q => \ELKS_ADDRB[4]\);
    
    \GP_PG.un1_ADDR_POINTER_0_I_20\ : AO1C
      port map(A => \ELKS_ADDRB[2]\, B => 
        \LOC_STOP_ADDR[2]_net_1\, C => N_2, Y => N_8);
    
    \GP_PG_SM_ns_i_i_o2[7]\ : OR2
      port map(A => N_214_li, B => OP_MODE_c_0, Y => N_47);
    
    \GP_PG.un1_ADDR_POINTER_0_I_15\ : OR2A
      port map(A => \ELKS_ADDRB[2]\, B => 
        \LOC_STOP_ADDR[2]_net_1\, Y => N_3);
    
    \GP_PG_SM[4]\ : DFN1C0
      port map(D => \GP_PG_SM_ns[6]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_29, Q => \GP_PG_SM[4]_net_1\);
    
    \GP_PG_SM_RNI5CBH[3]\ : OR2
      port map(A => \GP_PG_SM[3]_net_1\, B => \GP_PG_SM[2]_net_1\, 
        Y => N_39);
    
    \GP_PG_SM_RNO_0[2]\ : OR3C
      port map(A => OP_MODE_c_0, B => \GP_PG_SM[2]_net_1\, C => 
        N_214_li, Y => N_64);
    
    \GP_PG_SM_RNIAHBH[9]\ : NOR2
      port map(A => \GP_PG_SM[9]_net_1\, B => \GP_PG_SM[1]_net_1\, 
        Y => \GP_PG_SM_ns_0_a4_0[0]\);
    
    \RX_SER_WORD_2DEL[6]\ : DFN1C0
      port map(D => \RX_SER_WORD_1DEL[6]_net_1\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_26, Q => 
        \RX_SER_WORD_2DEL[6]_net_1\);
    
    \GP_PG.un1_ADDR_POINTER_0_I_11\ : OR2A
      port map(A => \LOC_STOP_ADDR[7]_net_1\, B => 
        \ELKS_ADDRB[7]\, Y => \ACT_LT3_E[4]\);
    
    \RX_SER_WORD_3DEL_RNIQTHB1[4]\ : OR3
      port map(A => \RX_SER_WORD_3DEL[5]_net_1\, B => 
        \RX_SER_WORD_3DEL[4]_net_1\, C => 
        un1_RX_SER_WORD_3DEL_NE_1, Y => un1_RX_SER_WORD_3DEL_NE_4);
    
    \RX_SER_WORD_3DEL_RNI4B3N2[0]\ : OR3
      port map(A => un1_RX_SER_WORD_3DEL_NE_3, B => 
        un1_RX_SER_WORD_3DEL_NE_2, C => un1_RX_SER_WORD_3DEL_NE_4, 
        Y => un1_RX_SER_WORD_3DEL_1);
    
    \GP_PG_SM_RNO_0[4]\ : NOR2A
      port map(A => \GP_PG_SM[6]_net_1\, B => OP_MODE_0, Y => 
        \GP_PG_SM_ns_0_a4_0[6]\);
    
    \LOC_STOP_ADDR[7]\ : DFN1E1C0
      port map(D => ELKS_STOP_ADDR(7), CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_7, E => \GP_PG_SM_0[10]_net_1\, Q => 
        \LOC_STOP_ADDR[7]_net_1\);
    
    \ADDR_POINTER_RNO[1]\ : NOR3
      port map(A => N_102, B => N_103, C => N_101, Y => N_36);
    
    \GP_PG_SM_0[10]\ : DFN1P0
      port map(D => \GP_PG_SM_ns[0]\, CLK => CLK_40M_GL, PRE => 
        P_MASTER_POR_B_c_34_0, Q => \GP_PG_SM_0[10]_net_1\);
    
    LOC_DIR_MODE_RNIB4Q8 : AO1C
      port map(A => N_213_li, B => ALIGN_ACTIVE, C => 
        P_USB_MASTER_EN_c, Y => N_45);
    
    \LOC_STRT_ADDR[2]\ : DFN1E1C0
      port map(D => ELKS_STRT_ADDR(2), CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_11, E => \GP_PG_SM_0[10]_net_1\, Q => 
        \LOC_STRT_ADDR[2]_net_1\);
    
    \RX_SER_WORD_2DEL[5]\ : DFN1C0
      port map(D => \RX_SER_WORD_1DEL[5]_net_1\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_26, Q => 
        \RX_SER_WORD_2DEL[5]_net_1\);
    
    \ADDR_POINTER_RNO_0[1]\ : NOR3A
      port map(A => N_42, B => \GP_PG_SM[10]_net_1\, C => I_30_0, 
        Y => N_102);
    
    \RX_SER_WORD_2DEL[3]\ : DFN1C0
      port map(D => \RX_SER_WORD_1DEL[3]_net_1\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_25, Q => 
        \RX_SER_WORD_2DEL[3]_net_1\);
    
    \GP_PG_SM_RNIN6A1K[10]\ : OA1B
      port map(A => N_107, B => \N_ADDR_POINTER_i_o2_0[7]\, C => 
        ELKS_STRT_ADDR(4), Y => N_375);
    
    \GP_PG_SM_RNO[6]\ : NOR3C
      port map(A => N_210_li, B => \GP_PG_SM[7]_net_1\, C => 
        N_116, Y => N_22);
    
    \GP_PG_SM_RNIGG4N9[10]\ : OA1A
      port map(A => N_39, B => N_214_li, C => 
        \GP_PG_SM[10]_net_1\, Y => \N_ADDR_POINTER_i_o2_0[7]\);
    
    \ADDR_POINTER_RNO_1[5]\ : NOR3A
      port map(A => N_39, B => N_214_li, C => 
        \LOC_STRT_ADDR[5]_net_1\, Y => N_374);
    
    \LOC_STRT_ADDR[3]\ : DFN1E1C0
      port map(D => ELKS_STRT_ADDR(3), CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_11, E => \GP_PG_SM_0[10]_net_1\, Q => 
        \LOC_STRT_ADDR[3]_net_1\);
    
    \LOC_STRT_ADDR[1]\ : DFN1E1C0
      port map(D => ELKS_STRT_ADDR(1), CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_11, E => \GP_PG_SM_0[10]_net_1\, Q => 
        \LOC_STRT_ADDR[1]_net_1\);
    
    \LOC_STRT_ADDR[7]\ : DFN1E1C0
      port map(D => ELKS_STRT_ADDR(7), CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_12, E => \GP_PG_SM[10]_net_1\, Q => 
        \LOC_STRT_ADDR[7]_net_1\);
    
    \RX_SER_WORD_2DEL_RNITKQC[6]\ : OR2A
      port map(A => \RX_SER_WORD_2DEL[7]_net_1\, B => 
        \RX_SER_WORD_2DEL[6]_net_1\, Y => 
        un1_RX_SER_WORD_2DEL_NE_1);
    
    \LOC_STRT_ADDR_RNIP2OG9[2]\ : NOR3A
      port map(A => N_39, B => N_214_li, C => 
        \LOC_STRT_ADDR[2]_net_1\, Y => N_383);
    
    \GP_PG_SM[8]\ : DFN1C0
      port map(D => N_80, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_29, Q => \GP_PG_SM[8]_net_1\);
    
    \GP_PG.un1_ADDR_POINTER_0_I_9\ : AND2A
      port map(A => \LOC_STOP_ADDR[6]_net_1\, B => 
        \ELKS_ADDRB[6]\, Y => \ACT_LT3_E[2]\);
    
    \GP_PG.un1_ADDR_POINTER_0_I_3\ : XNOR2
      port map(A => \ELKS_ADDRB[5]\, B => 
        \LOC_STOP_ADDR[5]_net_1\, Y => \DWACT_BL_EQUAL_0_E[0]\);
    
    \ADDR_POINTER_RNO_1[1]\ : NOR3A
      port map(A => N_39, B => N_214_li, C => 
        \LOC_STRT_ADDR[1]_net_1\, Y => N_103);
    
    \RX_SER_WORD_2DEL_RNIM5LP[4]\ : OR3
      port map(A => \RX_SER_WORD_2DEL[5]_net_1\, B => 
        \RX_SER_WORD_2DEL[4]_net_1\, C => 
        un1_RX_SER_WORD_2DEL_NE_1, Y => un1_RX_SER_WORD_2DEL_NE_4);
    
    \GP_PG_SM[3]\ : DFN1C0
      port map(D => \GP_PG_SM_RNO_0[3]_net_1\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_29, Q => \GP_PG_SM[3]_net_1\);
    
    \RX_SER_WORD_3DEL_RNO[7]\ : INV
      port map(A => \RX_SER_WORD_2DEL[7]_net_1\, Y => 
        \RX_SER_WORD_2DEL_i[7]\);
    
    \ADDR_POINTER[3]\ : DFN1C0
      port map(D => N_32, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_32, Q => \ELKS_ADDRB[3]\);
    
    \RX_SER_WORD_2DEL[1]\ : DFN1C0
      port map(D => \RX_SER_WORD_1DEL[1]_net_1\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_25, Q => 
        \RX_SER_WORD_2DEL[1]_net_1\);
    
    \GP_PG_SM_RNO_0[5]\ : NOR3B
      port map(A => \GP_PG_SM[8]_net_1\, B => N_114, C => 
        OP_MODE_0, Y => \GP_PG_SM_ns_0_a2_0_1[5]\);
    
    \GP_PG_SM_RNI81URC[10]\ : NOR3A
      port map(A => N_42, B => \GP_PG_SM[10]_net_1\, C => I_29_0, 
        Y => N_382);
    
    \GP_PG.un1_ADDR_POINTER_0_I_23\ : OA1A
      port map(A => N_6, B => N_8, C => N_7, Y => N_11);
    
    \GP_PG.un1_ADDR_POINTER_0_I_2\ : XNOR2
      port map(A => \ELKS_ADDRB[6]\, B => 
        \LOC_STOP_ADDR[6]_net_1\, Y => \DWACT_BL_EQUAL_0_E[1]\);
    
    \LOC_STRT_ADDR_RNICNURB1[6]\ : NOR3
      port map(A => N_86, B => N_88, C => N_87, Y => N_26);
    
    \GP_PG.un1_ADDR_POINTER_0_I_14\ : OR2A
      port map(A => \LOC_STOP_ADDR[1]_net_1\, B => 
        \ELKS_ADDRB[1]\, Y => N_2);
    
    \RX_SER_WORD_3DEL_RNO[3]\ : INV
      port map(A => \RX_SER_WORD_2DEL[3]_net_1\, Y => 
        \RX_SER_WORD_2DEL_i[3]\);
    
    \ADDR_POINTER_RNO[7]\ : NOR3
      port map(A => N_83, B => N_85, C => N_84, Y => N_24);
    
    \GP_PG.un1_ADDR_POINTER_0_I_8\ : OR2A
      port map(A => \LOC_STOP_ADDR[6]_net_1\, B => 
        \ELKS_ADDRB[6]\, Y => \ACT_LT3_E[1]\);
    
    \ADDR_POINTER[7]\ : DFN1C0
      port map(D => N_24, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_32, Q => \ELKS_ADDRB[7]\);
    
    \LOC_STOP_ADDR[3]\ : DFN1E1C0
      port map(D => ELKS_STOP_ADDR(3), CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_7, E => \GP_PG_SM_0[10]_net_1\, Q => 
        \LOC_STOP_ADDR[3]_net_1\);
    
    \RX_SER_WORD_1DEL[6]\ : DFN1C0
      port map(D => ELK_RX_SER_WORD_0(6), CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_23, Q => \RX_SER_WORD_1DEL[6]_net_1\);
    
    \RX_SER_WORD_2DEL[7]\ : DFN1C0
      port map(D => \RX_SER_WORD_1DEL[7]_net_1\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_26, Q => 
        \RX_SER_WORD_2DEL[7]_net_1\);
    
    \GP_PG_SM_RNO_1[7]\ : NOR3B
      port map(A => \GP_PG_SM[9]_net_1\, B => N_315, C => 
        N_213_li, Y => \GP_PG_SM_ns_0_a2_0_1[3]\);
    
    \GP_PG_SM_RNI5G1Q[8]\ : NOR2A
      port map(A => N_114, B => \GP_PG_SM[8]_net_1\, Y => N_315);
    
    un1_ADDR_POINTER_2_I_24 : XOR2
      port map(A => \ELKS_ADDRB[0]\, B => 
        \GP_PG_SM_RNIFMVG1[10]_net_1\, Y => 
        \DWACT_ADD_CI_0_partial_sum[0]\);
    
    \RX_SER_WORD_3DEL[6]\ : DFN1C0
      port map(D => \RX_SER_WORD_2DEL[6]_net_1\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_31_0, Q => 
        \RX_SER_WORD_3DEL[6]_net_1\);
    
    \GP_PG_SM_RNO[0]\ : AO1
      port map(A => \GP_PG_SM[0]_net_1\, B => OP_MODE_c_0, C => 
        \GP_PG_SM[1]_net_1\, Y => \GP_PG_SM_ns[10]\);
    
    \GP_PG_SM[9]\ : DFN1C0
      port map(D => N_69, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_29, Q => \GP_PG_SM[9]_net_1\);
    
    \ADDR_POINTER_RNO_2[5]\ : NOR3A
      port map(A => N_42, B => \GP_PG_SM[10]_net_1\, C => I_28_0, 
        Y => N_373);
    
    un1_ADDR_POINTER_2_I_41 : NOR2B
      port map(A => \DWACT_ADD_CI_0_g_array_2[0]\, B => 
        \DWACT_ADD_CI_0_pog_array_1_1[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_11[0]\);
    
    \GP_PG_SM_RNITU612[0]\ : NOR3C
      port map(A => N_315, B => \GP_PG_SM_ns_0_a4_0[0]\, C => 
        N_50, Y => \GP_PG_SM_ns_0_a4_2[0]\);
    
    \GP_PG.un1_ADDR_POINTER_0_I_22\ : AO1C
      port map(A => \ELKS_ADDRB[3]\, B => 
        \LOC_STOP_ADDR[3]_net_1\, C => N_5, Y => N_10);
    
    \RX_SER_WORD_2DEL[0]\ : DFN1C0
      port map(D => \RX_SER_WORD_1DEL[0]_net_1\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_25, Q => 
        \RX_SER_WORD_2DEL[0]_net_1\);
    
    \GP_PG_SM_RNILV0Q[0]\ : NOR2
      port map(A => \GP_PG_SM[0]_net_1\, B => N_39, Y => N_117);
    
    \GP_PG_SM_RNI9GBH[5]\ : OR2
      port map(A => \GP_PG_SM[5]_net_1\, B => \GP_PG_SM[4]_net_1\, 
        Y => N_40);
    
    \LOC_STOP_ADDR[0]\ : DFN1E1C0
      port map(D => ELKS_STOP_ADDR(0), CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_7, E => \GP_PG_SM_0[10]_net_1\, Q => 
        \LOC_STOP_ADDR[0]_net_1\);
    
    \RX_SER_WORD_1DEL[5]\ : DFN1C0
      port map(D => ELK_RX_SER_WORD_0(5), CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_23, Q => \RX_SER_WORD_1DEL[5]_net_1\);
    
    \GP_PG.un1_ADDR_POINTER_0_I_18\ : AO1C
      port map(A => \LOC_STOP_ADDR[1]_net_1\, B => 
        \ELKS_ADDRB[1]\, C => N_4, Y => N_6);
    
    \RX_SER_WORD_1DEL[3]\ : DFN1C0
      port map(D => ELK_RX_SER_WORD_0(3), CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_23, Q => \RX_SER_WORD_1DEL[3]_net_1\);
    
    \GP_PG_SM[2]\ : DFN1C0
      port map(D => \GP_PG_SM_RNO_0[2]_net_1\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_29, Q => \GP_PG_SM[2]_net_1\);
    
    un1_ADDR_POINTER_2_I_30 : XOR2
      port map(A => \ELKS_ADDRB[1]\, B => \DWACT_ADD_CI_0_TMP[0]\, 
        Y => I_30_0);
    
    \RX_SER_WORD_3DEL[5]\ : DFN1C0
      port map(D => \RX_SER_WORD_2DEL[5]_net_1\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_31_0, Q => 
        \RX_SER_WORD_3DEL[5]_net_1\);
    
    \GP_PG_SM_RNO[5]\ : AO1
      port map(A => \GP_PG_SM_ns_0_a2_0_1[5]\, B => N_25, C => 
        N_18, Y => \GP_PG_SM_ns[5]\);
    
    \GP_PG_SM_RNIO67Q9_0[5]\ : OR2
      port map(A => N_110, B => N_214_li, Y => N_42);
    
    \RX_SER_WORD_3DEL[3]\ : DFN1P0
      port map(D => \RX_SER_WORD_2DEL_i[3]\, CLK => CLK_40M_GL, 
        PRE => P_MASTER_POR_B_c_31_0, Q => 
        \RX_SER_WORD_3DEL_i_0[3]\);
    
    \GP_PG_SM_RNO[3]\ : AO1
      port map(A => \GP_PG_SM_ns_i_i_a4_0_1[7]\, B => N_116, C
         => N_76, Y => \GP_PG_SM_RNO_0[3]_net_1\);
    
    \GP_PG_SM_RNO_0[7]\ : NOR2A
      port map(A => \GP_PG_SM[7]_net_1\, B => N_210_li, Y => 
        \GP_PG_SM_ns_0_a2_0[3]\);
    
    \LOC_STRT_ADDR[4]\ : DFN1E1C0
      port map(D => ELKS_STRT_ADDR(4), CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_11, E => \GP_PG_SM_0[10]_net_1\, Q => 
        \LOC_STRT_ADDR[4]_net_1\);
    
    \GP_PG_SM_RNIESM21[5]\ : NOR2
      port map(A => N_40, B => N_39, Y => N_110);
    
    \GP_PG_SM_RNO[1]\ : NOR3
      port map(A => N_73, B => N_61, C => N_42, Y => 
        \GP_PG_SM_RNO_0[1]_net_1\);
    
    \ADDR_POINTER[5]\ : DFN1C0
      port map(D => N_28, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_32, Q => \ELKS_ADDRB[5]\);
    
    R_RWB : DFN1E1P0
      port map(D => N_213_li, CLK => CLK_40M_GL, PRE => 
        P_MASTER_POR_B_c_12, E => \GP_PG_SM[10]_net_1\, Q => 
        ELKS_RWB);
    
    R_BLKB_RNO_0 : NOR2
      port map(A => \GP_PG_SM[1]_net_1\, B => 
        \GP_PG_SM[10]_net_1\, Y => N_238);
    
    \ADDR_POINTER_RNO_1[3]\ : NOR3A
      port map(A => N_39, B => N_214_li, C => 
        \LOC_STRT_ADDR[3]_net_1\, Y => N_380);
    
    \GP_PG_SM_RNIEKTG3[0]\ : AO1
      port map(A => \GP_PG_SM_ns_0_a4_2[0]\, B => N_110, C => 
        N_72, Y => \GP_PG_SM_ns[0]\);
    
    \RX_SER_WORD_2DEL_RNI06DA4[0]\ : NOR2B
      port map(A => un1_RX_SER_WORD_2DEL_1, B => 
        un1_RX_SER_WORD_3DEL_1, Y => N_210_li);
    
    \RX_SER_WORD_2DEL[4]\ : DFN1C0
      port map(D => \RX_SER_WORD_1DEL[4]_net_1\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_25, Q => 
        \RX_SER_WORD_2DEL[4]_net_1\);
    
    \LOC_STRT_ADDR[6]\ : DFN1E1C0
      port map(D => ELKS_STRT_ADDR(6), CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_12, E => \GP_PG_SM[10]_net_1\, Q => 
        \LOC_STRT_ADDR[6]_net_1\);
    
    un1_ADDR_POINTER_2_I_44 : NOR2B
      port map(A => \DWACT_ADD_CI_0_g_array_11[0]\, B => 
        \ELKS_ADDRB[6]\, Y => \DWACT_ADD_CI_0_g_array_12_2[0]\);
    
    \RX_SER_WORD_2DEL[2]\ : DFN1C0
      port map(D => \RX_SER_WORD_1DEL[2]_net_1\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_25, Q => 
        \RX_SER_WORD_2DEL[2]_net_1\);
    
    \GP_PG_SM_RNO_0[1]\ : NOR2B
      port map(A => N_39, B => OP_MODE_c_0, Y => N_73);
    
    \LOC_STOP_ADDR[6]\ : DFN1E1C0
      port map(D => ELKS_STOP_ADDR(6), CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_7, E => \GP_PG_SM_0[10]_net_1\, Q => 
        \LOC_STOP_ADDR[6]_net_1\);
    
    \GP_PG.un1_ADDR_POINTER_0_I_10\ : AOI1A
      port map(A => \ACT_LT3_E[0]\, B => \ACT_LT3_E[1]\, C => 
        \ACT_LT3_E[2]\, Y => \ACT_LT3_E[3]\);
    
    \GP_PG_SM_RNID2TID[10]\ : NOR3A
      port map(A => N_42, B => \GP_PG_SM[10]_net_1\, C => I_33_0, 
        Y => N_376);
    
    \RX_SER_WORD_1DEL[1]\ : DFN1C0
      port map(D => ELK_RX_SER_WORD_0(1), CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_23, Q => \RX_SER_WORD_1DEL[1]_net_1\);
    
    un1_ADDR_POINTER_2_I_43 : NOR2B
      port map(A => \DWACT_ADD_CI_0_g_array_2[0]\, B => 
        \ELKS_ADDRB[4]\, Y => \DWACT_ADD_CI_0_g_array_12_1[0]\);
    
    \GP_PG.un1_ADDR_POINTER_0_I_16\ : NOR2A
      port map(A => \LOC_STOP_ADDR[0]_net_1\, B => 
        \ELKS_ADDRB[0]\, Y => N_4);
    
    \RX_SER_WORD_3DEL[1]\ : DFN1P0
      port map(D => \RX_SER_WORD_2DEL_i[1]\, CLK => CLK_40M_GL, 
        PRE => P_MASTER_POR_B_c_31_0, Q => 
        \RX_SER_WORD_3DEL_i_0[1]\);
    
    \ADDR_POINTER_RNO_0[3]\ : NOR3A
      port map(A => N_42, B => \GP_PG_SM[10]_net_1\, C => I_27_0, 
        Y => N_379);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SER320M_3_34 is

    port( TFC_TX_DAT             : in    std_logic_vector(7 downto 0);
          TFC_OUT_R              : out   std_logic;
          TFC_OUT_F              : out   std_logic;
          MASTER_DCB_POR_B_i_0_i : in    std_logic;
          CCC_160M_FXD           : in    std_logic;
          CLK_40M_GL             : in    std_logic
        );

end SER320M_3_34;

architecture DEF_ARCH of SER320M_3_34 is 

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \N_SER_CMD_WORD_R[0]\, \START_RISE\, 
        \N_SER_CMD_WORD_F[0]\, \N_SER_CMD_WORD_R[3]\, 
        \SER_CMD_WORD_R[2]_net_1\, \N_SER_CMD_WORD_R[2]\, 
        \SER_CMD_WORD_R[1]_net_1\, \N_SER_CMD_WORD_R[1]\, 
        \SER_CMD_WORD_R[0]_net_1\, \N_SER_CMD_WORD_F[3]\, 
        \SER_CMD_WORD_F[2]_net_1\, \N_SER_CMD_WORD_F[2]\, 
        \SER_CMD_WORD_F[1]_net_1\, \N_SER_CMD_WORD_F[1]\, 
        \SER_CMD_WORD_F[0]_net_1\, N_START_RISE, 
        \CLK40M_GEN_DEL0\, \SER_OUT_FI\, \SER_OUT_RI\, 
        \SER_CMD_WORD_F[3]_net_1\, \SER_CMD_WORD_R[3]_net_1\, 
        \GND\, \VCC\ : std_logic;

begin 


    SER_OUT_FI : DFN1C0
      port map(D => \SER_CMD_WORD_F[3]_net_1\, CLK => 
        CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \SER_OUT_FI\);
    
    \SER_CMD_WORD_F[3]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[3]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \SER_CMD_WORD_F[3]_net_1\);
    
    \SER_CMD_WORD_R[1]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[1]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \SER_CMD_WORD_R[1]_net_1\);
    
    \SER_CMD_WORD_R[2]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[2]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \SER_CMD_WORD_R[2]_net_1\);
    
    \SER_CMD_WORD_R_RNO[3]\ : MX2
      port map(A => \SER_CMD_WORD_R[2]_net_1\, B => TFC_TX_DAT(7), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_R[3]\);
    
    \SER_CMD_WORD_R_RNO[0]\ : NOR2B
      port map(A => \START_RISE\, B => TFC_TX_DAT(1), Y => 
        \N_SER_CMD_WORD_R[0]\);
    
    \SER_CMD_WORD_F[0]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[0]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \SER_CMD_WORD_F[0]_net_1\);
    
    \SER_CMD_WORD_R_RNO[1]\ : MX2
      port map(A => \SER_CMD_WORD_R[0]_net_1\, B => TFC_TX_DAT(3), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_R[1]\);
    
    \SER_CMD_WORD_F_RNO[2]\ : MX2
      port map(A => \SER_CMD_WORD_F[1]_net_1\, B => TFC_TX_DAT(4), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_F[2]\);
    
    \SER_CMD_WORD_F_RNO[3]\ : MX2
      port map(A => \SER_CMD_WORD_F[2]_net_1\, B => TFC_TX_DAT(6), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_F[3]\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    CLK40M_GEN_DEL0 : DFN1C0
      port map(D => CLK_40M_GL, CLK => CCC_160M_FXD, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \CLK40M_GEN_DEL0\);
    
    SER_OUT_RI : DFN1C0
      port map(D => \SER_CMD_WORD_R[3]_net_1\, CLK => 
        CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \SER_OUT_RI\);
    
    \SER_CMD_WORD_F[2]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[2]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \SER_CMD_WORD_F[2]_net_1\);
    
    \SER_CMD_WORD_F_RNO[1]\ : MX2
      port map(A => \SER_CMD_WORD_F[0]_net_1\, B => TFC_TX_DAT(2), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_F[1]\);
    
    \SER_CMD_WORD_R[0]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[0]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \SER_CMD_WORD_R[0]_net_1\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    START_RISE : DFN1C0
      port map(D => N_START_RISE, CLK => CCC_160M_FXD, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \START_RISE\);
    
    \SER_CMD_WORD_R[3]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[3]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \SER_CMD_WORD_R[3]_net_1\);
    
    \SER_CMD_WORD_F_RNO[0]\ : NOR2B
      port map(A => \START_RISE\, B => TFC_TX_DAT(0), Y => 
        \N_SER_CMD_WORD_F[0]\);
    
    SER_OUT_RDEL : DFN1C0
      port map(D => \SER_OUT_RI\, CLK => CCC_160M_FXD, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => TFC_OUT_R);
    
    \SER_CMD_WORD_F[1]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[1]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \SER_CMD_WORD_F[1]_net_1\);
    
    START_RISE_RNO : NOR2B
      port map(A => \CLK40M_GEN_DEL0\, B => CLK_40M_GL, Y => 
        N_START_RISE);
    
    \SER_CMD_WORD_R_RNO[2]\ : MX2
      port map(A => \SER_CMD_WORD_R[1]_net_1\, B => TFC_TX_DAT(5), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_R[2]\);
    
    SER_OUT_FDEL : DFN1C0
      port map(D => \SER_OUT_FI\, CLK => CCC_160M_FXD, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => TFC_OUT_F);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SER320M_3_34_0 is

    port( ELK0_TX_DAT                : in    std_logic_vector(7 downto 0);
          MASTER_SALT_POR_B_i_0_i_17 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_3  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_7  : in    std_logic;
          ELK0_OUT_R_i_0             : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_10 : in    std_logic;
          ELK0_OUT_F_i_0             : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_5  : in    std_logic;
          CLK_40M_GL                 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_13 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_14 : in    std_logic;
          CCC_160M_FXD               : in    std_logic
        );

end SER320M_3_34_0;

architecture DEF_ARCH of SER320M_3_34_0 is 

  component DFI1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          QN  : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component DFN1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

    signal SER_OUT_RI_i, \SER_CMD_WORD_R[3]_net_1\, SER_OUT_FI_i, 
        \SER_CMD_WORD_F[3]_net_1\, \N_SER_CMD_WORD_R[0]\, 
        \START_RISE\, \N_SER_CMD_WORD_F[0]\, 
        \N_SER_CMD_WORD_R[3]\, \SER_CMD_WORD_R[2]_net_1\, 
        \N_SER_CMD_WORD_R[2]\, \SER_CMD_WORD_R[1]_net_1\, 
        \N_SER_CMD_WORD_R[1]\, \SER_CMD_WORD_R[0]_net_1\, 
        \N_SER_CMD_WORD_F[3]\, \SER_CMD_WORD_F[2]_net_1\, 
        \N_SER_CMD_WORD_F[2]\, \SER_CMD_WORD_F[1]_net_1\, 
        \N_SER_CMD_WORD_F[1]\, \SER_CMD_WORD_F[0]_net_1\, 
        N_START_RISE, \CLK40M_GEN_DEL0\, \GND\, \VCC\
         : std_logic;

begin 


    SER_OUT_FI : DFI1C0
      port map(D => \SER_CMD_WORD_F[3]_net_1\, CLK => 
        CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_13, QN => 
        SER_OUT_FI_i);
    
    \SER_CMD_WORD_F[3]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[3]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_17, Q => 
        \SER_CMD_WORD_F[3]_net_1\);
    
    \SER_CMD_WORD_R[1]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[1]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_14, Q => 
        \SER_CMD_WORD_R[1]_net_1\);
    
    \SER_CMD_WORD_R[2]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[2]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_14, Q => 
        \SER_CMD_WORD_R[2]_net_1\);
    
    \SER_CMD_WORD_R_RNO[3]\ : MX2
      port map(A => \SER_CMD_WORD_R[2]_net_1\, B => 
        ELK0_TX_DAT(7), S => \START_RISE\, Y => 
        \N_SER_CMD_WORD_R[3]\);
    
    \SER_CMD_WORD_R_RNO[0]\ : NOR2B
      port map(A => \START_RISE\, B => ELK0_TX_DAT(1), Y => 
        \N_SER_CMD_WORD_R[0]\);
    
    \SER_CMD_WORD_F[0]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[0]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_17, Q => 
        \SER_CMD_WORD_F[0]_net_1\);
    
    \SER_CMD_WORD_R_RNO[1]\ : MX2
      port map(A => \SER_CMD_WORD_R[0]_net_1\, B => 
        ELK0_TX_DAT(3), S => \START_RISE\, Y => 
        \N_SER_CMD_WORD_R[1]\);
    
    \SER_CMD_WORD_F_RNO[2]\ : MX2
      port map(A => \SER_CMD_WORD_F[1]_net_1\, B => 
        ELK0_TX_DAT(4), S => \START_RISE\, Y => 
        \N_SER_CMD_WORD_F[2]\);
    
    \SER_CMD_WORD_F_RNO[3]\ : MX2
      port map(A => \SER_CMD_WORD_F[2]_net_1\, B => 
        ELK0_TX_DAT(6), S => \START_RISE\, Y => 
        \N_SER_CMD_WORD_F[3]\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    CLK40M_GEN_DEL0 : DFN1C0
      port map(D => CLK_40M_GL, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_5, Q => \CLK40M_GEN_DEL0\);
    
    SER_OUT_RI : DFI1C0
      port map(D => \SER_CMD_WORD_R[3]_net_1\, CLK => 
        CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_14, QN => 
        SER_OUT_RI_i);
    
    \SER_CMD_WORD_F[2]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[2]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_17, Q => 
        \SER_CMD_WORD_F[2]_net_1\);
    
    \SER_CMD_WORD_F_RNO[1]\ : MX2
      port map(A => \SER_CMD_WORD_F[0]_net_1\, B => 
        ELK0_TX_DAT(2), S => \START_RISE\, Y => 
        \N_SER_CMD_WORD_F[1]\);
    
    \SER_CMD_WORD_R[0]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[0]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_14, Q => 
        \SER_CMD_WORD_R[0]_net_1\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    START_RISE : DFN1C0
      port map(D => N_START_RISE, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_3, Q => \START_RISE\);
    
    \SER_CMD_WORD_R[3]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[3]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_14, Q => 
        \SER_CMD_WORD_R[3]_net_1\);
    
    \SER_CMD_WORD_F_RNO[0]\ : NOR2B
      port map(A => \START_RISE\, B => ELK0_TX_DAT(0), Y => 
        \N_SER_CMD_WORD_F[0]\);
    
    SER_OUT_RDEL : DFN1P0
      port map(D => SER_OUT_RI_i, CLK => CCC_160M_FXD, PRE => 
        MASTER_SALT_POR_B_i_0_i_7, Q => ELK0_OUT_R_i_0);
    
    \SER_CMD_WORD_F[1]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[1]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_17, Q => 
        \SER_CMD_WORD_F[1]_net_1\);
    
    START_RISE_RNO : NOR2B
      port map(A => \CLK40M_GEN_DEL0\, B => CLK_40M_GL, Y => 
        N_START_RISE);
    
    \SER_CMD_WORD_R_RNO[2]\ : MX2
      port map(A => \SER_CMD_WORD_R[1]_net_1\, B => 
        ELK0_TX_DAT(5), S => \START_RISE\, Y => 
        \N_SER_CMD_WORD_R[2]\);
    
    SER_OUT_FDEL : DFN1P0
      port map(D => SER_OUT_FI_i, CLK => CCC_160M_FXD, PRE => 
        MASTER_SALT_POR_B_i_0_i_10, Q => ELK0_OUT_F_i_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SLAVE_DES320S_1_17_10 is

    port( ELK_RX_SER_WORD_12     : out   std_logic_vector(7 downto 0);
          BIT_OS_SEL_5_0         : in    std_logic;
          BIT_OS_SEL_6           : in    std_logic_vector(2 downto 1);
          BIT_OS_SEL_4           : in    std_logic_vector(2 downto 1);
          BIT_OS_SEL_3_0         : in    std_logic;
          CLK_40M_GL             : in    std_logic;
          CCC_160M_FXD           : in    std_logic;
          ELK_IN_R               : in    std_logic;
          ELK_IN_F               : in    std_logic;
          MASTER_DCB_POR_B_i_0_i : in    std_logic;
          CCC_160M_ADJ           : in    std_logic
        );

end SLAVE_DES320S_1_17_10;

architecture DEF_ARCH of SLAVE_DES320S_1_17_10 is 

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal N_17, \ARB_BYTE[0]_net_1\, \ARB_BYTE[4]_net_1\, N_18, 
        \ARB_BYTE[1]_net_1\, \ARB_BYTE[5]_net_1\, N_19, 
        \ARB_BYTE[2]_net_1\, \ARB_BYTE[6]_net_1\, N_20, 
        \ARB_BYTE[3]_net_1\, \ARB_BYTE[7]_net_1\, N_21, 
        \ARB_BYTE[8]_net_1\, N_22, \ARB_BYTE[9]_net_1\, N_23, 
        \ARB_BYTE[10]_net_1\, N_24, \ARB_BYTE[11]_net_1\, N_31, 
        \ARB_BYTE[12]_net_1\, N_32, \ARB_BYTE[13]_net_1\, N_33, 
        N_34, N_35, N_36, N_37, N_38, N_39, N_40, N_56, 
        \ARB_BYTE[14]_net_1\, N_64, \N_RECD_SER_WORD[0]\, 
        \N_RECD_SER_WORD[1]\, \N_RECD_SER_WORD[2]\, 
        \N_RECD_SER_WORD[3]\, \N_RECD_SER_WORD[4]\, 
        \N_RECD_SER_WORD[5]\, \N_RECD_SER_WORD[6]\, 
        \N_RECD_SER_WORD[7]\, \ADJ_SER_IN_F_0DEL\, 
        \ADJ_SER_IN_R_0DEL\, \ADJ_SER_IN_F_1DEL\, 
        \ADJ_SER_IN_R_1DEL\, \Q[0]_net_1\, \ADJ_Q[0]_net_1\, 
        \Q[1]_net_1\, \ADJ_Q[1]_net_1\, \Q[2]_net_1\, 
        \ADJ_Q[2]_net_1\, \Q[3]_net_1\, \ADJ_Q[3]_net_1\, 
        \Q[4]_net_1\, \ADJ_Q[4]_net_1\, \Q[5]_net_1\, 
        \ADJ_Q[5]_net_1\, \Q[6]_net_1\, \ADJ_Q[6]_net_1\, 
        \Q[7]_net_1\, \ADJ_Q[7]_net_1\, \Q[8]_net_1\, 
        \ADJ_Q[8]_net_1\, \Q[9]_net_1\, \ADJ_Q[9]_net_1\, 
        \Q[10]_net_1\, \ADJ_Q[10]_net_1\, \Q[11]_net_1\, 
        \ADJ_Q[11]_net_1\, \Q[12]_net_1\, \ADJ_Q[12]_net_1\, 
        \Q[13]_net_1\, \ADJ_Q[13]_net_1\, \Q[14]_net_1\, 
        \ADJ_Q[14]_net_1\, \ARB_WRD_40M_FIXED[0]_net_1\, 
        \ARB_WRD_40M_FIXED[1]_net_1\, 
        \ARB_WRD_40M_FIXED[2]_net_1\, 
        \ARB_WRD_40M_FIXED[3]_net_1\, 
        \ARB_WRD_40M_FIXED[4]_net_1\, 
        \ARB_WRD_40M_FIXED[5]_net_1\, 
        \ARB_WRD_40M_FIXED[6]_net_1\, 
        \ARB_WRD_40M_FIXED[7]_net_1\, 
        \ARB_WRD_40M_FIXED[8]_net_1\, 
        \ARB_WRD_40M_FIXED[9]_net_1\, 
        \ARB_WRD_40M_FIXED[10]_net_1\, 
        \ARB_WRD_40M_FIXED[11]_net_1\, 
        \ARB_WRD_40M_FIXED[12]_net_1\, 
        \ARB_WRD_40M_FIXED[13]_net_1\, 
        \ARB_WRD_40M_FIXED[14]_net_1\, \GND\, \VCC\ : std_logic;

begin 


    \RECD_SER_WORD_RNO[5]\ : MX2
      port map(A => N_38, B => N_39, S => BIT_OS_SEL_5_0, Y => 
        \N_RECD_SER_WORD[5]\);
    
    \ARB_WRD_40M_FIXED[9]\ : DFN1C0
      port map(D => \Q[9]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[9]_net_1\);
    
    \ADJ_Q[4]\ : DFN1C0
      port map(D => \ADJ_Q[2]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[4]_net_1\);
    
    \ARB_BYTE[6]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[6]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[6]_net_1\);
    
    ADJ_SER_IN_F_1DEL : DFN1C0
      port map(D => \ADJ_SER_IN_F_0DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_F_1DEL\);
    
    \ARB_BYTE[0]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[0]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[0]_net_1\);
    
    \Q[11]\ : DFN1C0
      port map(D => \ADJ_Q[11]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[11]_net_1\);
    
    \ADJ_Q[8]\ : DFN1C0
      port map(D => \ADJ_Q[6]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[8]_net_1\);
    
    \ARB_BYTE_RNILV6T1[13]\ : MX2
      port map(A => N_24, B => N_32, S => BIT_OS_SEL_4(1), Y => 
        N_40);
    
    \ADJ_Q[6]\ : DFN1C0
      port map(D => \ADJ_Q[4]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[6]_net_1\);
    
    \ADJ_Q[12]\ : DFN1C0
      port map(D => \ADJ_Q[10]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[12]_net_1\);
    
    \RECD_SER_WORD_RNO_1[0]\ : MX2
      port map(A => \ARB_BYTE[0]_net_1\, B => \ARB_BYTE[4]_net_1\, 
        S => BIT_OS_SEL_3_0, Y => N_17);
    
    \Q[1]\ : DFN1C0
      port map(D => \ADJ_Q[1]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[1]_net_1\);
    
    \ARB_BYTE[4]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[4]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[4]_net_1\);
    
    \ADJ_Q[2]\ : DFN1C0
      port map(D => \ADJ_Q[0]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[2]_net_1\);
    
    \RECD_SER_WORD_RNO_1[7]\ : MX2
      port map(A => \ARB_BYTE[10]_net_1\, B => 
        \ARB_BYTE[14]_net_1\, S => BIT_OS_SEL_6(2), Y => N_56);
    
    \RECD_SER_WORD[4]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[4]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_12(4));
    
    \Q[5]\ : DFN1C0
      port map(D => \ADJ_Q[5]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[5]_net_1\);
    
    \ADJ_Q[11]\ : DFN1C0
      port map(D => \ADJ_Q[9]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[11]_net_1\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \ADJ_Q[3]\ : DFN1C0
      port map(D => \ADJ_Q[1]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[3]_net_1\);
    
    \Q[10]\ : DFN1C0
      port map(D => \ADJ_Q[10]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[10]_net_1\);
    
    \ARB_BYTE_RNI1BDT[3]\ : MX2
      port map(A => \ARB_BYTE[3]_net_1\, B => \ARB_BYTE[7]_net_1\, 
        S => BIT_OS_SEL_3_0, Y => N_20);
    
    \ARB_WRD_40M_FIXED[6]\ : DFN1C0
      port map(D => \Q[6]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[6]_net_1\);
    
    \ARB_WRD_40M_FIXED[1]\ : DFN1C0
      port map(D => \Q[1]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[1]_net_1\);
    
    \RECD_SER_WORD[3]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[3]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_12(3));
    
    \RECD_SER_WORD[0]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[0]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_12(0));
    
    \RECD_SER_WORD_RNO[3]\ : MX2
      port map(A => N_36, B => N_37, S => BIT_OS_SEL_5_0, Y => 
        \N_RECD_SER_WORD[3]\);
    
    \Q[0]\ : DFN1C0
      port map(D => \ADJ_Q[0]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[0]_net_1\);
    
    \ARB_BYTE_RNIL8DT1[3]\ : MX2
      port map(A => N_20, B => N_22, S => BIT_OS_SEL_4(1), Y => 
        N_36);
    
    \ARB_BYTE_RNIHR6T1[10]\ : MX2
      port map(A => N_23, B => N_31, S => BIT_OS_SEL_4(1), Y => 
        N_39);
    
    \RECD_SER_WORD_RNO_0[7]\ : MX2
      port map(A => N_31, B => N_56, S => BIT_OS_SEL_6(1), Y => 
        N_64);
    
    \Q[7]\ : DFN1C0
      port map(D => \ADJ_Q[7]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[7]_net_1\);
    
    \ARB_BYTE_RNIT6DT[1]\ : MX2
      port map(A => \ARB_BYTE[1]_net_1\, B => \ARB_BYTE[5]_net_1\, 
        S => BIT_OS_SEL_3_0, Y => N_18);
    
    \ARB_BYTE[14]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[14]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[14]_net_1\);
    
    \ARB_WRD_40M_FIXED[2]\ : DFN1C0
      port map(D => \Q[2]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[2]_net_1\);
    
    \ARB_WRD_40M_FIXED[14]\ : DFN1C0
      port map(D => \Q[14]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[14]_net_1\);
    
    \RECD_SER_WORD_RNO[2]\ : MX2
      port map(A => N_35, B => N_36, S => BIT_OS_SEL_5_0, Y => 
        \N_RECD_SER_WORD[2]\);
    
    \ARB_BYTE[2]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[2]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[2]_net_1\);
    
    \ARB_BYTE_RNI10AT1[10]\ : MX2
      port map(A => N_21, B => N_23, S => BIT_OS_SEL_4(1), Y => 
        N_37);
    
    \ADJ_Q[7]\ : DFN1C0
      port map(D => \ADJ_Q[5]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[7]_net_1\);
    
    \ARB_BYTE_RNID0DT1[1]\ : MX2
      port map(A => N_18, B => N_20, S => BIT_OS_SEL_4(1), Y => 
        N_34);
    
    \ARB_BYTE[8]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[8]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[8]_net_1\);
    
    \RECD_SER_WORD[5]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[5]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_12(5));
    
    \ARB_BYTE[12]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[12]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[12]_net_1\);
    
    \RECD_SER_WORD[1]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[1]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_12(1));
    
    \Q[3]\ : DFN1C0
      port map(D => \ADJ_Q[3]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[3]_net_1\);
    
    \ARB_BYTE_RNIF4AT[10]\ : MX2
      port map(A => \ARB_BYTE[6]_net_1\, B => 
        \ARB_BYTE[10]_net_1\, S => BIT_OS_SEL_4(2), Y => N_23);
    
    ADJ_SER_IN_F_0DEL : DFN1C0
      port map(D => ELK_IN_F, CLK => CCC_160M_ADJ, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_F_0DEL\);
    
    \RECD_SER_WORD_RNO[7]\ : MX2
      port map(A => N_40, B => N_64, S => BIT_OS_SEL_5_0, Y => 
        \N_RECD_SER_WORD[7]\);
    
    \RECD_SER_WORD_RNO[1]\ : MX2
      port map(A => N_34, B => N_35, S => BIT_OS_SEL_5_0, Y => 
        \N_RECD_SER_WORD[1]\);
    
    \ARB_WRD_40M_FIXED[4]\ : DFN1C0
      port map(D => \Q[4]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[4]_net_1\);
    
    \RECD_SER_WORD_RNO[0]\ : MX2
      port map(A => N_33, B => N_34, S => BIT_OS_SEL_5_0, Y => 
        \N_RECD_SER_WORD[0]\);
    
    \Q[6]\ : DFN1C0
      port map(D => \ADJ_Q[6]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[6]_net_1\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \ARB_WRD_40M_FIXED[8]\ : DFN1C0
      port map(D => \Q[8]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[8]_net_1\);
    
    \ARB_BYTE[11]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[11]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[11]_net_1\);
    
    \Q[9]\ : DFN1C0
      port map(D => \ADJ_Q[9]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[9]_net_1\);
    
    \Q[14]\ : DFN1C0
      port map(D => \ADJ_Q[14]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[14]_net_1\);
    
    ADJ_SER_IN_R_0DEL : DFN1C0
      port map(D => ELK_IN_R, CLK => CCC_160M_ADJ, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_R_0DEL\);
    
    \Q[13]\ : DFN1C0
      port map(D => \ADJ_Q[13]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[13]_net_1\);
    
    \ARB_BYTE_RNIJ8AT[12]\ : MX2
      port map(A => \ARB_BYTE[8]_net_1\, B => 
        \ARB_BYTE[12]_net_1\, S => BIT_OS_SEL_4(2), Y => N_31);
    
    \ARB_BYTE[9]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[9]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[9]_net_1\);
    
    ADJ_SER_IN_R_1DEL : DFN1C0
      port map(D => \ADJ_SER_IN_R_0DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_R_1DEL\);
    
    \ARB_BYTE[10]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[10]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[10]_net_1\);
    
    \ADJ_Q[9]\ : DFN1C0
      port map(D => \ADJ_Q[7]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[9]_net_1\);
    
    \RECD_SER_WORD[7]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[7]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_12(7));
    
    \ARB_WRD_40M_FIXED[5]\ : DFN1C0
      port map(D => \Q[5]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[5]_net_1\);
    
    \ARB_WRD_40M_FIXED[12]\ : DFN1C0
      port map(D => \Q[12]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[12]_net_1\);
    
    \ARB_BYTE_RNILAAT[13]\ : MX2
      port map(A => \ARB_BYTE[9]_net_1\, B => 
        \ARB_BYTE[13]_net_1\, S => BIT_OS_SEL_4(2), Y => N_32);
    
    \ARB_WRD_40M_FIXED[11]\ : DFN1C0
      port map(D => \Q[11]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[11]_net_1\);
    
    \ARB_WRD_40M_FIXED[0]\ : DFN1C0
      port map(D => \Q[0]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[0]_net_1\);
    
    \ADJ_Q[10]\ : DFN1C0
      port map(D => \ADJ_Q[8]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[10]_net_1\);
    
    \Q[2]\ : DFN1C0
      port map(D => \ADJ_Q[2]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[2]_net_1\);
    
    \ARB_BYTE_RNIH4DT1[2]\ : MX2
      port map(A => N_19, B => N_21, S => BIT_OS_SEL_4(1), Y => 
        N_35);
    
    \ARB_BYTE_RNI54AT1[11]\ : MX2
      port map(A => N_22, B => N_24, S => BIT_OS_SEL_4(1), Y => 
        N_38);
    
    \ADJ_Q[1]\ : DFN1C0
      port map(D => \ADJ_SER_IN_F_1DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[1]_net_1\);
    
    \RECD_SER_WORD[6]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[6]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_12(6));
    
    \RECD_SER_WORD[2]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[2]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_12(2));
    
    \ADJ_Q[13]\ : DFN1C0
      port map(D => \ADJ_Q[11]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[13]_net_1\);
    
    \ARB_BYTE_RNIV8DT[2]\ : MX2
      port map(A => \ARB_BYTE[2]_net_1\, B => \ARB_BYTE[6]_net_1\, 
        S => BIT_OS_SEL_3_0, Y => N_19);
    
    \Q[8]\ : DFN1C0
      port map(D => \ADJ_Q[8]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[8]_net_1\);
    
    \ARB_BYTE[5]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[5]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[5]_net_1\);
    
    \ADJ_Q[14]\ : DFN1C0
      port map(D => \ADJ_Q[12]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[14]_net_1\);
    
    \RECD_SER_WORD_RNO[4]\ : MX2
      port map(A => N_37, B => N_38, S => BIT_OS_SEL_5_0, Y => 
        \N_RECD_SER_WORD[4]\);
    
    \Q[12]\ : DFN1C0
      port map(D => \ADJ_Q[12]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[12]_net_1\);
    
    \ARB_BYTE[13]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[13]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[13]_net_1\);
    
    \ARB_BYTE_RNI3DDT[4]\ : MX2
      port map(A => \ARB_BYTE[4]_net_1\, B => \ARB_BYTE[8]_net_1\, 
        S => BIT_OS_SEL_3_0, Y => N_21);
    
    \ARB_WRD_40M_FIXED[3]\ : DFN1C0
      port map(D => \Q[3]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[3]_net_1\);
    
    \ARB_BYTE[7]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[7]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[7]_net_1\);
    
    \RECD_SER_WORD_RNO_0[0]\ : MX2
      port map(A => N_17, B => N_19, S => BIT_OS_SEL_4(1), Y => 
        N_33);
    
    \Q[4]\ : DFN1C0
      port map(D => \ADJ_Q[4]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[4]_net_1\);
    
    \ARB_WRD_40M_FIXED[7]\ : DFN1C0
      port map(D => \Q[7]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[7]_net_1\);
    
    \ARB_BYTE_RNI5FDT[5]\ : MX2
      port map(A => \ARB_BYTE[5]_net_1\, B => \ARB_BYTE[9]_net_1\, 
        S => BIT_OS_SEL_3_0, Y => N_22);
    
    \RECD_SER_WORD_RNO[6]\ : MX2
      port map(A => N_39, B => N_40, S => BIT_OS_SEL_5_0, Y => 
        \N_RECD_SER_WORD[6]\);
    
    \ARB_BYTE[3]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[3]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[3]_net_1\);
    
    \ARB_BYTE_RNIH6AT[11]\ : MX2
      port map(A => \ARB_BYTE[7]_net_1\, B => 
        \ARB_BYTE[11]_net_1\, S => BIT_OS_SEL_4(2), Y => N_24);
    
    \ADJ_Q[5]\ : DFN1C0
      port map(D => \ADJ_Q[3]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[5]_net_1\);
    
    \ARB_BYTE[1]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[1]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[1]_net_1\);
    
    \ARB_WRD_40M_FIXED[13]\ : DFN1C0
      port map(D => \Q[13]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[13]_net_1\);
    
    \ADJ_Q[0]\ : DFN1C0
      port map(D => \ADJ_SER_IN_R_1DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[0]_net_1\);
    
    \ARB_WRD_40M_FIXED[10]\ : DFN1C0
      port map(D => \Q[10]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[10]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SER320M_3_34_12 is

    port( ELK_TX_DAT                 : in    std_logic_vector(7 downto 0);
          MASTER_SALT_POR_B_i_0_i_15 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_10 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_0  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_8  : in    std_logic;
          ELK_OUT_R                  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_12 : in    std_logic;
          ELK_OUT_F                  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_6  : in    std_logic;
          CCC_160M_FXD               : in    std_logic;
          CLK_40M_GL                 : in    std_logic
        );

end SER320M_3_34_12;

architecture DEF_ARCH of SER320M_3_34_12 is 

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \N_SER_CMD_WORD_R[0]\, \START_RISE\, 
        \N_SER_CMD_WORD_F[0]\, \N_SER_CMD_WORD_R[3]\, 
        \SER_CMD_WORD_R[2]_net_1\, \N_SER_CMD_WORD_R[2]\, 
        \SER_CMD_WORD_R[1]_net_1\, \N_SER_CMD_WORD_R[1]\, 
        \SER_CMD_WORD_R[0]_net_1\, \N_SER_CMD_WORD_F[3]\, 
        \SER_CMD_WORD_F[2]_net_1\, \N_SER_CMD_WORD_F[2]\, 
        \SER_CMD_WORD_F[1]_net_1\, \N_SER_CMD_WORD_F[1]\, 
        \SER_CMD_WORD_F[0]_net_1\, N_START_RISE, 
        \CLK40M_GEN_DEL0\, \SER_OUT_FI\, \SER_OUT_RI\, 
        \SER_CMD_WORD_F[3]_net_1\, \SER_CMD_WORD_R[3]_net_1\, 
        \GND\, \VCC\ : std_logic;

begin 


    SER_OUT_FI : DFN1C0
      port map(D => \SER_CMD_WORD_F[3]_net_1\, CLK => 
        CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_10, Q => 
        \SER_OUT_FI\);
    
    \SER_CMD_WORD_F[3]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[3]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_15, Q => 
        \SER_CMD_WORD_F[3]_net_1\);
    
    \SER_CMD_WORD_R[1]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[1]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_12, Q => 
        \SER_CMD_WORD_R[1]_net_1\);
    
    \SER_CMD_WORD_R[2]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[2]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_12, Q => 
        \SER_CMD_WORD_R[2]_net_1\);
    
    \SER_CMD_WORD_R_RNO[3]\ : MX2
      port map(A => \SER_CMD_WORD_R[2]_net_1\, B => ELK_TX_DAT(7), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_R[3]\);
    
    \SER_CMD_WORD_R_RNO[0]\ : NOR2B
      port map(A => \START_RISE\, B => ELK_TX_DAT(1), Y => 
        \N_SER_CMD_WORD_R[0]\);
    
    \SER_CMD_WORD_F[0]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[0]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_15, Q => 
        \SER_CMD_WORD_F[0]_net_1\);
    
    \SER_CMD_WORD_R_RNO[1]\ : MX2
      port map(A => \SER_CMD_WORD_R[0]_net_1\, B => ELK_TX_DAT(3), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_R[1]\);
    
    \SER_CMD_WORD_F_RNO[2]\ : MX2
      port map(A => \SER_CMD_WORD_F[1]_net_1\, B => ELK_TX_DAT(4), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_F[2]\);
    
    \SER_CMD_WORD_F_RNO[3]\ : MX2
      port map(A => \SER_CMD_WORD_F[2]_net_1\, B => ELK_TX_DAT(6), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_F[3]\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    CLK40M_GEN_DEL0 : DFN1C0
      port map(D => CLK_40M_GL, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_6, Q => \CLK40M_GEN_DEL0\);
    
    SER_OUT_RI : DFN1C0
      port map(D => \SER_CMD_WORD_R[3]_net_1\, CLK => 
        CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_10, Q => 
        \SER_OUT_RI\);
    
    \SER_CMD_WORD_F[2]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[2]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_15, Q => 
        \SER_CMD_WORD_F[2]_net_1\);
    
    \SER_CMD_WORD_F_RNO[1]\ : MX2
      port map(A => \SER_CMD_WORD_F[0]_net_1\, B => ELK_TX_DAT(2), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_F[1]\);
    
    \SER_CMD_WORD_R[0]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[0]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_12, Q => 
        \SER_CMD_WORD_R[0]_net_1\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    START_RISE : DFN1C0
      port map(D => N_START_RISE, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_0, Q => \START_RISE\);
    
    \SER_CMD_WORD_R[3]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[3]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_12, Q => 
        \SER_CMD_WORD_R[3]_net_1\);
    
    \SER_CMD_WORD_F_RNO[0]\ : NOR2B
      port map(A => \START_RISE\, B => ELK_TX_DAT(0), Y => 
        \N_SER_CMD_WORD_F[0]\);
    
    SER_OUT_RDEL : DFN1C0
      port map(D => \SER_OUT_RI\, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_8, Q => ELK_OUT_R);
    
    \SER_CMD_WORD_F[1]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[1]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_15, Q => 
        \SER_CMD_WORD_F[1]_net_1\);
    
    START_RISE_RNO : NOR2B
      port map(A => \CLK40M_GEN_DEL0\, B => CLK_40M_GL, Y => 
        N_START_RISE);
    
    \SER_CMD_WORD_R_RNO[2]\ : MX2
      port map(A => \SER_CMD_WORD_R[1]_net_1\, B => ELK_TX_DAT(5), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_R[2]\);
    
    SER_OUT_FDEL : DFN1C0
      port map(D => \SER_OUT_FI\, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_12, Q => ELK_OUT_F);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity DDR_BIDIR_LVDS_DUAL_CLK_12 is

    port( DCB_SALT_SEL_c_i : in    std_logic;
          ELK12_DAT_P      : inout std_logic := 'Z';
          ELK12_DAT_N      : inout std_logic := 'Z';
          ELK_OUT_R        : in    std_logic;
          ELK_OUT_F        : in    std_logic;
          CCC_160M_FXD     : in    std_logic;
          CCC_160M_ADJ     : in    std_logic;
          ELK_IN_DDR_R     : out   std_logic;
          ELK_IN_DDR_F     : out   std_logic
        );

end DDR_BIDIR_LVDS_DUAL_CLK_12;

architecture DEF_ARCH of DDR_BIDIR_LVDS_DUAL_CLK_12 is 

  component DDR_REG
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          QR  : out   std_logic;
          QF  : out   std_logic
        );
  end component;

  component DDR_OUT
    port( DR  : in    std_logic := 'U';
          DF  : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component BIBUF_LVDS
    port( PADP : inout   std_logic;
          PADN : inout   std_logic;
          D    : in    std_logic := 'U';
          E    : in    std_logic := 'U';
          Y    : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal DDR_BIDIR_LVDS_DUAL_CLK_12_GND, BIBUF_LVDS_0_Y, 
        DDR_OUT_0_Q, \VCC\ : std_logic;

begin 


    DDR_REG_0 : DDR_REG
      port map(D => BIBUF_LVDS_0_Y, CLK => CCC_160M_ADJ, CLR => 
        DDR_BIDIR_LVDS_DUAL_CLK_12_GND, QR => ELK_IN_DDR_R, QF
         => ELK_IN_DDR_F);
    
    DDR_OUT_0 : DDR_OUT
      port map(DR => ELK_OUT_R, DF => ELK_OUT_F, CLK => 
        CCC_160M_FXD, CLR => DDR_BIDIR_LVDS_DUAL_CLK_12_GND, Q
         => DDR_OUT_0_Q);
    
    BIBUF_LVDS_0 : BIBUF_LVDS
      port map(PADP => ELK12_DAT_P, PADN => ELK12_DAT_N, D => 
        DDR_OUT_0_Q, E => DCB_SALT_SEL_c_i, Y => BIBUF_LVDS_0_Y);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    GND_i : GND
      port map(Y => DDR_BIDIR_LVDS_DUAL_CLK_12_GND);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SYNC_DAT_SEL_12 is

    port( ELK_TX_DAT                : out   std_logic_vector(7 downto 0);
          PATT_ELK_DAT_12           : in    std_logic_vector(7 downto 0);
          OP_MODE_c_3_0             : in    std_logic;
          OP_MODE_c_2_0             : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_2 : in    std_logic;
          CLK_40M_GL                : in    std_logic
        );

end SYNC_DAT_SEL_12;

architecture DEF_ARCH of SYNC_DAT_SEL_12 is 

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \N_SERDAT[0]\, \N_SERDAT[1]\, \N_SERDAT[2]\, 
        \N_SERDAT[3]\, \N_SERDAT[4]\, \N_SERDAT[5]\, 
        \N_SERDAT[6]\, \N_SERDAT[7]\, \GND\, \VCC\ : std_logic;

begin 


    \SERDAT_RNO[4]\ : NOR2A
      port map(A => PATT_ELK_DAT_12(4), B => OP_MODE_c_3_0, Y => 
        \N_SERDAT[4]\);
    
    \SERDAT_RNO[0]\ : NOR2A
      port map(A => PATT_ELK_DAT_12(0), B => OP_MODE_c_2_0, Y => 
        \N_SERDAT[0]\);
    
    \SERDAT[6]\ : DFN1C0
      port map(D => \N_SERDAT[6]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_2, Q => ELK_TX_DAT(6));
    
    \SERDAT[4]\ : DFN1C0
      port map(D => \N_SERDAT[4]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_2, Q => ELK_TX_DAT(4));
    
    \SERDAT_RNO[7]\ : OR2
      port map(A => PATT_ELK_DAT_12(7), B => OP_MODE_c_3_0, Y => 
        \N_SERDAT[7]\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \SERDAT_RNO[3]\ : OR2
      port map(A => PATT_ELK_DAT_12(3), B => OP_MODE_c_3_0, Y => 
        \N_SERDAT[3]\);
    
    \SERDAT_RNO[2]\ : OR2
      port map(A => PATT_ELK_DAT_12(2), B => OP_MODE_c_3_0, Y => 
        \N_SERDAT[2]\);
    
    \SERDAT[5]\ : DFN1C0
      port map(D => \N_SERDAT[5]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_2, Q => ELK_TX_DAT(5));
    
    \SERDAT[7]\ : DFN1C0
      port map(D => \N_SERDAT[7]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_2, Q => ELK_TX_DAT(7));
    
    GND_i : GND
      port map(Y => \GND\);
    
    \SERDAT_RNO[5]\ : NOR2A
      port map(A => PATT_ELK_DAT_12(5), B => OP_MODE_c_3_0, Y => 
        \N_SERDAT[5]\);
    
    \SERDAT[0]\ : DFN1C0
      port map(D => \N_SERDAT[0]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_2, Q => ELK_TX_DAT(0));
    
    \SERDAT_RNO[6]\ : NOR2A
      port map(A => PATT_ELK_DAT_12(6), B => OP_MODE_c_3_0, Y => 
        \N_SERDAT[6]\);
    
    \SERDAT[1]\ : DFN1C0
      port map(D => \N_SERDAT[1]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_2, Q => ELK_TX_DAT(1));
    
    \SERDAT_RNO[1]\ : OR2
      port map(A => PATT_ELK_DAT_12(1), B => OP_MODE_c_2_0, Y => 
        \N_SERDAT[1]\);
    
    \SERDAT[3]\ : DFN1C0
      port map(D => \N_SERDAT[3]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_2, Q => ELK_TX_DAT(3));
    
    \SERDAT[2]\ : DFN1C0
      port map(D => \N_SERDAT[2]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_2, Q => ELK_TX_DAT(2));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity ELINK_SLAVE_15_7 is

    port( BIT_OS_SEL_3_0             : in    std_logic;
          BIT_OS_SEL_4               : in    std_logic_vector(2 downto 1);
          BIT_OS_SEL_6               : in    std_logic_vector(2 downto 1);
          BIT_OS_SEL_5_0             : in    std_logic;
          ELK_RX_SER_WORD_12         : out   std_logic_vector(7 downto 0);
          OP_MODE_c_2_0              : in    std_logic;
          OP_MODE_c_3_0              : in    std_logic;
          PATT_ELK_DAT_12            : in    std_logic_vector(7 downto 0);
          MASTER_DCB_POR_B_i_0_i     : in    std_logic;
          ELK12_DAT_N                : inout std_logic := 'Z';
          ELK12_DAT_P                : inout std_logic := 'Z';
          DCB_SALT_SEL_c_i           : in    std_logic;
          CCC_160M_FXD               : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_6  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_12 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_8  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_0  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_10 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_15 : in    std_logic;
          CLK_40M_GL                 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_2  : in    std_logic;
          DEV_RST_B_c                : in    std_logic;
          CCC_160M_ADJ               : in    std_logic
        );

end ELINK_SLAVE_15_7;

architecture DEF_ARCH of ELINK_SLAVE_15_7 is 

  component SLAVE_DES320S_1_17_10
    port( ELK_RX_SER_WORD_12     : out   std_logic_vector(7 downto 0);
          BIT_OS_SEL_5_0         : in    std_logic := 'U';
          BIT_OS_SEL_6           : in    std_logic_vector(2 downto 1) := (others => 'U');
          BIT_OS_SEL_4           : in    std_logic_vector(2 downto 1) := (others => 'U');
          BIT_OS_SEL_3_0         : in    std_logic := 'U';
          CLK_40M_GL             : in    std_logic := 'U';
          CCC_160M_FXD           : in    std_logic := 'U';
          ELK_IN_R               : in    std_logic := 'U';
          ELK_IN_F               : in    std_logic := 'U';
          MASTER_DCB_POR_B_i_0_i : in    std_logic := 'U';
          CCC_160M_ADJ           : in    std_logic := 'U'
        );
  end component;

  component SER320M_3_34_12
    port( ELK_TX_DAT                 : in    std_logic_vector(7 downto 0) := (others => 'U');
          MASTER_SALT_POR_B_i_0_i_15 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_10 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_0  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_8  : in    std_logic := 'U';
          ELK_OUT_R                  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_12 : in    std_logic := 'U';
          ELK_OUT_F                  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_6  : in    std_logic := 'U';
          CCC_160M_FXD               : in    std_logic := 'U';
          CLK_40M_GL                 : in    std_logic := 'U'
        );
  end component;

  component DDR_BIDIR_LVDS_DUAL_CLK_12
    port( DCB_SALT_SEL_c_i : in    std_logic := 'U';
          ELK12_DAT_P      : inout   std_logic;
          ELK12_DAT_N      : inout   std_logic;
          ELK_OUT_R        : in    std_logic := 'U';
          ELK_OUT_F        : in    std_logic := 'U';
          CCC_160M_FXD     : in    std_logic := 'U';
          CCC_160M_ADJ     : in    std_logic := 'U';
          ELK_IN_DDR_R     : out   std_logic;
          ELK_IN_DDR_F     : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component SYNC_DAT_SEL_12
    port( ELK_TX_DAT                : out   std_logic_vector(7 downto 0);
          PATT_ELK_DAT_12           : in    std_logic_vector(7 downto 0) := (others => 'U');
          OP_MODE_c_3_0             : in    std_logic := 'U';
          OP_MODE_c_2_0             : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_2 : in    std_logic := 'U';
          CLK_40M_GL                : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \ELK_IN_F\, ELK_IN_DDR_F, \ELK_IN_R\, ELK_IN_DDR_R, 
        \ELK_TX_DAT[0]\, \ELK_TX_DAT[1]\, \ELK_TX_DAT[2]\, 
        \ELK_TX_DAT[3]\, \ELK_TX_DAT[4]\, \ELK_TX_DAT[5]\, 
        \ELK_TX_DAT[6]\, \ELK_TX_DAT[7]\, ELK_OUT_R, ELK_OUT_F, 
        \GND\, \VCC\ : std_logic;

    for all : SLAVE_DES320S_1_17_10
	Use entity work.SLAVE_DES320S_1_17_10(DEF_ARCH);
    for all : SER320M_3_34_12
	Use entity work.SER320M_3_34_12(DEF_ARCH);
    for all : DDR_BIDIR_LVDS_DUAL_CLK_12
	Use entity work.DDR_BIDIR_LVDS_DUAL_CLK_12(DEF_ARCH);
    for all : SYNC_DAT_SEL_12
	Use entity work.SYNC_DAT_SEL_12(DEF_ARCH);
begin 


    U_SLAVE_1ELK : SLAVE_DES320S_1_17_10
      port map(ELK_RX_SER_WORD_12(7) => ELK_RX_SER_WORD_12(7), 
        ELK_RX_SER_WORD_12(6) => ELK_RX_SER_WORD_12(6), 
        ELK_RX_SER_WORD_12(5) => ELK_RX_SER_WORD_12(5), 
        ELK_RX_SER_WORD_12(4) => ELK_RX_SER_WORD_12(4), 
        ELK_RX_SER_WORD_12(3) => ELK_RX_SER_WORD_12(3), 
        ELK_RX_SER_WORD_12(2) => ELK_RX_SER_WORD_12(2), 
        ELK_RX_SER_WORD_12(1) => ELK_RX_SER_WORD_12(1), 
        ELK_RX_SER_WORD_12(0) => ELK_RX_SER_WORD_12(0), 
        BIT_OS_SEL_5_0 => BIT_OS_SEL_5_0, BIT_OS_SEL_6(2) => 
        BIT_OS_SEL_6(2), BIT_OS_SEL_6(1) => BIT_OS_SEL_6(1), 
        BIT_OS_SEL_4(2) => BIT_OS_SEL_4(2), BIT_OS_SEL_4(1) => 
        BIT_OS_SEL_4(1), BIT_OS_SEL_3_0 => BIT_OS_SEL_3_0, 
        CLK_40M_GL => CLK_40M_GL, CCC_160M_FXD => CCC_160M_FXD, 
        ELK_IN_R => \ELK_IN_R\, ELK_IN_F => \ELK_IN_F\, 
        MASTER_DCB_POR_B_i_0_i => MASTER_DCB_POR_B_i_0_i, 
        CCC_160M_ADJ => CCC_160M_ADJ);
    
    U_ELK1_CMD_TX : SER320M_3_34_12
      port map(ELK_TX_DAT(7) => \ELK_TX_DAT[7]\, ELK_TX_DAT(6)
         => \ELK_TX_DAT[6]\, ELK_TX_DAT(5) => \ELK_TX_DAT[5]\, 
        ELK_TX_DAT(4) => \ELK_TX_DAT[4]\, ELK_TX_DAT(3) => 
        \ELK_TX_DAT[3]\, ELK_TX_DAT(2) => \ELK_TX_DAT[2]\, 
        ELK_TX_DAT(1) => \ELK_TX_DAT[1]\, ELK_TX_DAT(0) => 
        \ELK_TX_DAT[0]\, MASTER_SALT_POR_B_i_0_i_15 => 
        MASTER_SALT_POR_B_i_0_i_15, MASTER_SALT_POR_B_i_0_i_10
         => MASTER_SALT_POR_B_i_0_i_10, MASTER_SALT_POR_B_i_0_i_0
         => MASTER_SALT_POR_B_i_0_i_0, MASTER_SALT_POR_B_i_0_i_8
         => MASTER_SALT_POR_B_i_0_i_8, ELK_OUT_R => ELK_OUT_R, 
        MASTER_SALT_POR_B_i_0_i_12 => MASTER_SALT_POR_B_i_0_i_12, 
        ELK_OUT_F => ELK_OUT_F, MASTER_SALT_POR_B_i_0_i_6 => 
        MASTER_SALT_POR_B_i_0_i_6, CCC_160M_FXD => CCC_160M_FXD, 
        CLK_40M_GL => CLK_40M_GL);
    
    U_DDR_ELK1 : DDR_BIDIR_LVDS_DUAL_CLK_12
      port map(DCB_SALT_SEL_c_i => DCB_SALT_SEL_c_i, ELK12_DAT_P
         => ELK12_DAT_P, ELK12_DAT_N => ELK12_DAT_N, ELK_OUT_R
         => ELK_OUT_R, ELK_OUT_F => ELK_OUT_F, CCC_160M_FXD => 
        CCC_160M_FXD, CCC_160M_ADJ => CCC_160M_ADJ, ELK_IN_DDR_R
         => ELK_IN_DDR_R, ELK_IN_DDR_F => ELK_IN_DDR_F);
    
    ELK_IN_F : DFN1C0
      port map(D => ELK_IN_DDR_F, CLK => CCC_160M_ADJ, CLR => 
        DEV_RST_B_c, Q => \ELK_IN_F\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    U_ELK1_SERDAT_SOURCE : SYNC_DAT_SEL_12
      port map(ELK_TX_DAT(7) => \ELK_TX_DAT[7]\, ELK_TX_DAT(6)
         => \ELK_TX_DAT[6]\, ELK_TX_DAT(5) => \ELK_TX_DAT[5]\, 
        ELK_TX_DAT(4) => \ELK_TX_DAT[4]\, ELK_TX_DAT(3) => 
        \ELK_TX_DAT[3]\, ELK_TX_DAT(2) => \ELK_TX_DAT[2]\, 
        ELK_TX_DAT(1) => \ELK_TX_DAT[1]\, ELK_TX_DAT(0) => 
        \ELK_TX_DAT[0]\, PATT_ELK_DAT_12(7) => PATT_ELK_DAT_12(7), 
        PATT_ELK_DAT_12(6) => PATT_ELK_DAT_12(6), 
        PATT_ELK_DAT_12(5) => PATT_ELK_DAT_12(5), 
        PATT_ELK_DAT_12(4) => PATT_ELK_DAT_12(4), 
        PATT_ELK_DAT_12(3) => PATT_ELK_DAT_12(3), 
        PATT_ELK_DAT_12(2) => PATT_ELK_DAT_12(2), 
        PATT_ELK_DAT_12(1) => PATT_ELK_DAT_12(1), 
        PATT_ELK_DAT_12(0) => PATT_ELK_DAT_12(0), OP_MODE_c_3_0
         => OP_MODE_c_3_0, OP_MODE_c_2_0 => OP_MODE_c_2_0, 
        MASTER_SALT_POR_B_i_0_i_2 => MASTER_SALT_POR_B_i_0_i_2, 
        CLK_40M_GL => CLK_40M_GL);
    
    ELK_IN_R : DFN1C0
      port map(D => ELK_IN_DDR_R, CLK => CCC_160M_ADJ, CLR => 
        DEV_RST_B_c, Q => \ELK_IN_R\);
    
    GND_i : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SLAVE_DES320S_1_17_11 is

    port( ELK_RX_SER_WORD_13     : out   std_logic_vector(7 downto 0);
          BIT_OS_SEL_4_0         : in    std_logic;
          BIT_OS_SEL_5_0         : in    std_logic;
          BIT_OS_SEL_6_0         : in    std_logic;
          BIT_OS_SEL_3           : in    std_logic_vector(2 downto 1);
          BIT_OS_SEL_2_0         : in    std_logic;
          CLK_40M_GL             : in    std_logic;
          CCC_160M_FXD           : in    std_logic;
          ELK_IN_R               : in    std_logic;
          ELK_IN_F               : in    std_logic;
          MASTER_DCB_POR_B_i_0_i : in    std_logic;
          CCC_160M_ADJ           : in    std_logic
        );

end SLAVE_DES320S_1_17_11;

architecture DEF_ARCH of SLAVE_DES320S_1_17_11 is 

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal N_17, \ARB_BYTE[0]_net_1\, \ARB_BYTE[4]_net_1\, N_18, 
        \ARB_BYTE[1]_net_1\, \ARB_BYTE[5]_net_1\, N_19, 
        \ARB_BYTE[2]_net_1\, \ARB_BYTE[6]_net_1\, N_20, 
        \ARB_BYTE[3]_net_1\, \ARB_BYTE[7]_net_1\, N_21, 
        \ARB_BYTE[8]_net_1\, N_22, \ARB_BYTE[9]_net_1\, N_23, 
        \ARB_BYTE[10]_net_1\, N_24, \ARB_BYTE[11]_net_1\, N_31, 
        \ARB_BYTE[12]_net_1\, N_32, \ARB_BYTE[13]_net_1\, N_33, 
        N_34, N_35, N_36, N_37, N_38, N_39, N_40, N_56, 
        \ARB_BYTE[14]_net_1\, N_64, \N_RECD_SER_WORD[0]\, 
        \N_RECD_SER_WORD[1]\, \N_RECD_SER_WORD[2]\, 
        \N_RECD_SER_WORD[3]\, \N_RECD_SER_WORD[4]\, 
        \N_RECD_SER_WORD[5]\, \N_RECD_SER_WORD[6]\, 
        \N_RECD_SER_WORD[7]\, \ADJ_SER_IN_F_0DEL\, 
        \ADJ_SER_IN_R_0DEL\, \ADJ_SER_IN_F_1DEL\, 
        \ADJ_SER_IN_R_1DEL\, \Q[0]_net_1\, \ADJ_Q[0]_net_1\, 
        \Q[1]_net_1\, \ADJ_Q[1]_net_1\, \Q[2]_net_1\, 
        \ADJ_Q[2]_net_1\, \Q[3]_net_1\, \ADJ_Q[3]_net_1\, 
        \Q[4]_net_1\, \ADJ_Q[4]_net_1\, \Q[5]_net_1\, 
        \ADJ_Q[5]_net_1\, \Q[6]_net_1\, \ADJ_Q[6]_net_1\, 
        \Q[7]_net_1\, \ADJ_Q[7]_net_1\, \Q[8]_net_1\, 
        \ADJ_Q[8]_net_1\, \Q[9]_net_1\, \ADJ_Q[9]_net_1\, 
        \Q[10]_net_1\, \ADJ_Q[10]_net_1\, \Q[11]_net_1\, 
        \ADJ_Q[11]_net_1\, \Q[12]_net_1\, \ADJ_Q[12]_net_1\, 
        \Q[13]_net_1\, \ADJ_Q[13]_net_1\, \Q[14]_net_1\, 
        \ADJ_Q[14]_net_1\, \ARB_WRD_40M_FIXED[0]_net_1\, 
        \ARB_WRD_40M_FIXED[1]_net_1\, 
        \ARB_WRD_40M_FIXED[2]_net_1\, 
        \ARB_WRD_40M_FIXED[3]_net_1\, 
        \ARB_WRD_40M_FIXED[4]_net_1\, 
        \ARB_WRD_40M_FIXED[5]_net_1\, 
        \ARB_WRD_40M_FIXED[6]_net_1\, 
        \ARB_WRD_40M_FIXED[7]_net_1\, 
        \ARB_WRD_40M_FIXED[8]_net_1\, 
        \ARB_WRD_40M_FIXED[9]_net_1\, 
        \ARB_WRD_40M_FIXED[10]_net_1\, 
        \ARB_WRD_40M_FIXED[11]_net_1\, 
        \ARB_WRD_40M_FIXED[12]_net_1\, 
        \ARB_WRD_40M_FIXED[13]_net_1\, 
        \ARB_WRD_40M_FIXED[14]_net_1\, \GND\, \VCC\ : std_logic;

begin 


    \RECD_SER_WORD_RNO[5]\ : MX2
      port map(A => N_38, B => N_39, S => BIT_OS_SEL_4_0, Y => 
        \N_RECD_SER_WORD[5]\);
    
    \ARB_WRD_40M_FIXED[9]\ : DFN1C0
      port map(D => \Q[9]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[9]_net_1\);
    
    \ADJ_Q[4]\ : DFN1C0
      port map(D => \ADJ_Q[2]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[4]_net_1\);
    
    \ARB_BYTE_RNIKUOM[12]\ : MX2
      port map(A => \ARB_BYTE[8]_net_1\, B => 
        \ARB_BYTE[12]_net_1\, S => BIT_OS_SEL_3(2), Y => N_31);
    
    \ARB_BYTE[6]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[6]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[6]_net_1\);
    
    ADJ_SER_IN_F_1DEL : DFN1C0
      port map(D => \ADJ_SER_IN_F_0DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_F_1DEL\);
    
    \ARB_BYTE[0]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[0]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[0]_net_1\);
    
    \Q[11]\ : DFN1C0
      port map(D => \ADJ_Q[11]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[11]_net_1\);
    
    \ADJ_Q[8]\ : DFN1C0
      port map(D => \ADJ_Q[6]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[8]_net_1\);
    
    \ADJ_Q[6]\ : DFN1C0
      port map(D => \ADJ_Q[4]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[6]_net_1\);
    
    \ADJ_Q[12]\ : DFN1C0
      port map(D => \ADJ_Q[10]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[12]_net_1\);
    
    \RECD_SER_WORD_RNO_1[0]\ : MX2
      port map(A => \ARB_BYTE[0]_net_1\, B => \ARB_BYTE[4]_net_1\, 
        S => BIT_OS_SEL_2_0, Y => N_17);
    
    \Q[1]\ : DFN1C0
      port map(D => \ADJ_Q[1]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[1]_net_1\);
    
    \ARB_BYTE[4]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[4]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[4]_net_1\);
    
    \ADJ_Q[2]\ : DFN1C0
      port map(D => \ADJ_Q[0]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[2]_net_1\);
    
    \RECD_SER_WORD_RNO_1[7]\ : MX2
      port map(A => \ARB_BYTE[10]_net_1\, B => 
        \ARB_BYTE[14]_net_1\, S => BIT_OS_SEL_6_0, Y => N_56);
    
    \RECD_SER_WORD[4]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[4]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_13(4));
    
    \Q[5]\ : DFN1C0
      port map(D => \ADJ_Q[5]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[5]_net_1\);
    
    \ADJ_Q[11]\ : DFN1C0
      port map(D => \ADJ_Q[9]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[11]_net_1\);
    
    \ARB_BYTE_RNIOLLR[3]\ : MX2
      port map(A => N_20, B => N_22, S => BIT_OS_SEL_3(1), Y => 
        N_36);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \ADJ_Q[3]\ : DFN1C0
      port map(D => \ADJ_Q[1]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[3]_net_1\);
    
    \Q[10]\ : DFN1C0
      port map(D => \ADJ_Q[10]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[10]_net_1\);
    
    \ARB_WRD_40M_FIXED[6]\ : DFN1C0
      port map(D => \Q[6]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[6]_net_1\);
    
    \ARB_WRD_40M_FIXED[1]\ : DFN1C0
      port map(D => \Q[1]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[1]_net_1\);
    
    \RECD_SER_WORD[3]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[3]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_13(3));
    
    \RECD_SER_WORD[0]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[0]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_13(0));
    
    \ARB_BYTE_RNIURVB[1]\ : MX2
      port map(A => \ARB_BYTE[1]_net_1\, B => \ARB_BYTE[5]_net_1\, 
        S => BIT_OS_SEL_2_0, Y => N_18);
    
    \ARB_BYTE_RNI773D[5]\ : MX2
      port map(A => \ARB_BYTE[5]_net_1\, B => \ARB_BYTE[9]_net_1\, 
        S => BIT_OS_SEL_3(2), Y => N_22);
    
    \ARB_BYTE_RNI0UVB[2]\ : MX2
      port map(A => \ARB_BYTE[2]_net_1\, B => \ARB_BYTE[6]_net_1\, 
        S => BIT_OS_SEL_2_0, Y => N_19);
    
    \RECD_SER_WORD_RNO[3]\ : MX2
      port map(A => N_36, B => N_37, S => BIT_OS_SEL_4_0, Y => 
        \N_RECD_SER_WORD[3]\);
    
    \Q[0]\ : DFN1C0
      port map(D => \ADJ_Q[0]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[0]_net_1\);
    
    \RECD_SER_WORD_RNO_0[7]\ : MX2
      port map(A => N_31, B => N_56, S => BIT_OS_SEL_5_0, Y => 
        N_64);
    
    \Q[7]\ : DFN1C0
      port map(D => \ADJ_Q[7]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[7]_net_1\);
    
    \ARB_BYTE[14]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[14]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[14]_net_1\);
    
    \ARB_WRD_40M_FIXED[2]\ : DFN1C0
      port map(D => \Q[2]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[2]_net_1\);
    
    \ARB_WRD_40M_FIXED[14]\ : DFN1C0
      port map(D => \Q[14]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[14]_net_1\);
    
    \RECD_SER_WORD_RNO[2]\ : MX2
      port map(A => N_35, B => N_36, S => BIT_OS_SEL_4_0, Y => 
        \N_RECD_SER_WORD[2]\);
    
    \ARB_BYTE[2]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[2]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[2]_net_1\);
    
    \ARB_BYTE_RNI333D[3]\ : MX2
      port map(A => \ARB_BYTE[3]_net_1\, B => \ARB_BYTE[7]_net_1\, 
        S => BIT_OS_SEL_3(2), Y => N_20);
    
    \ADJ_Q[7]\ : DFN1C0
      port map(D => \ADJ_Q[5]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[7]_net_1\);
    
    \ARB_BYTE[8]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[8]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[8]_net_1\);
    
    \RECD_SER_WORD[5]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[5]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_13(5));
    
    \ARB_BYTE[12]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[12]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[12]_net_1\);
    
    \ARB_BYTE_RNIM81F1[13]\ : MX2
      port map(A => N_24, B => N_32, S => BIT_OS_SEL_3(1), Y => 
        N_40);
    
    \RECD_SER_WORD[1]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[1]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_13(1));
    
    \ARB_BYTE_RNIJEIQ[2]\ : MX2
      port map(A => N_19, B => N_21, S => BIT_OS_SEL_3(1), Y => 
        N_35);
    
    \Q[3]\ : DFN1C0
      port map(D => \ADJ_Q[3]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[3]_net_1\);
    
    ADJ_SER_IN_F_0DEL : DFN1C0
      port map(D => ELK_IN_F, CLK => CCC_160M_ADJ, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_F_0DEL\);
    
    \RECD_SER_WORD_RNO[7]\ : MX2
      port map(A => N_40, B => N_64, S => BIT_OS_SEL_4_0, Y => 
        \N_RECD_SER_WORD[7]\);
    
    \RECD_SER_WORD_RNO[1]\ : MX2
      port map(A => N_34, B => N_35, S => BIT_OS_SEL_4_0, Y => 
        \N_RECD_SER_WORD[1]\);
    
    \ARB_WRD_40M_FIXED[4]\ : DFN1C0
      port map(D => \Q[4]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[4]_net_1\);
    
    \ARB_BYTE_RNI7FB51[5]\ : MX2
      port map(A => N_22, B => N_24, S => BIT_OS_SEL_3(1), Y => 
        N_38);
    
    \RECD_SER_WORD_RNO[0]\ : MX2
      port map(A => N_33, B => N_34, S => BIT_OS_SEL_4_0, Y => 
        \N_RECD_SER_WORD[0]\);
    
    \Q[6]\ : DFN1C0
      port map(D => \ADJ_Q[6]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[6]_net_1\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \ARB_WRD_40M_FIXED[8]\ : DFN1C0
      port map(D => \Q[8]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[8]_net_1\);
    
    \ARB_BYTE[11]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[11]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[11]_net_1\);
    
    \Q[9]\ : DFN1C0
      port map(D => \ADJ_Q[9]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[9]_net_1\);
    
    \Q[14]\ : DFN1C0
      port map(D => \ADJ_Q[14]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[14]_net_1\);
    
    ADJ_SER_IN_R_0DEL : DFN1C0
      port map(D => ELK_IN_R, CLK => CCC_160M_ADJ, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_R_0DEL\);
    
    \Q[13]\ : DFN1C0
      port map(D => \ADJ_Q[13]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[13]_net_1\);
    
    \ARB_BYTE[9]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[9]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[9]_net_1\);
    
    ADJ_SER_IN_R_1DEL : DFN1C0
      port map(D => \ADJ_SER_IN_R_0DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_R_1DEL\);
    
    \ARB_BYTE[10]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[10]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[10]_net_1\);
    
    \ADJ_Q[9]\ : DFN1C0
      port map(D => \ADJ_Q[7]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[9]_net_1\);
    
    \RECD_SER_WORD[7]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[7]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_13(7));
    
    \ARB_WRD_40M_FIXED[5]\ : DFN1C0
      port map(D => \Q[5]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[5]_net_1\);
    
    \ARB_WRD_40M_FIXED[12]\ : DFN1C0
      port map(D => \Q[12]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[12]_net_1\);
    
    \ARB_BYTE_RNIISOM[11]\ : MX2
      port map(A => \ARB_BYTE[7]_net_1\, B => 
        \ARB_BYTE[11]_net_1\, S => BIT_OS_SEL_3(2), Y => N_24);
    
    \ARB_BYTE_RNI3BB51[4]\ : MX2
      port map(A => N_21, B => N_23, S => BIT_OS_SEL_3(1), Y => 
        N_37);
    
    \ARB_WRD_40M_FIXED[11]\ : DFN1C0
      port map(D => \Q[11]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[11]_net_1\);
    
    \ARB_BYTE_RNIFAIQ[1]\ : MX2
      port map(A => N_18, B => N_20, S => BIT_OS_SEL_3(1), Y => 
        N_34);
    
    \ARB_WRD_40M_FIXED[0]\ : DFN1C0
      port map(D => \Q[0]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[0]_net_1\);
    
    \ADJ_Q[10]\ : DFN1C0
      port map(D => \ADJ_Q[8]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[10]_net_1\);
    
    \Q[2]\ : DFN1C0
      port map(D => \ADJ_Q[2]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[2]_net_1\);
    
    \ADJ_Q[1]\ : DFN1C0
      port map(D => \ADJ_SER_IN_F_1DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[1]_net_1\);
    
    \RECD_SER_WORD[6]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[6]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_13(6));
    
    \RECD_SER_WORD[2]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[2]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_13(2));
    
    \ADJ_Q[13]\ : DFN1C0
      port map(D => \ADJ_Q[11]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[13]_net_1\);
    
    \Q[8]\ : DFN1C0
      port map(D => \ADJ_Q[8]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[8]_net_1\);
    
    \ARB_BYTE[5]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[5]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[5]_net_1\);
    
    \ADJ_Q[14]\ : DFN1C0
      port map(D => \ADJ_Q[12]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[14]_net_1\);
    
    \RECD_SER_WORD_RNO[4]\ : MX2
      port map(A => N_37, B => N_38, S => BIT_OS_SEL_4_0, Y => 
        \N_RECD_SER_WORD[4]\);
    
    \Q[12]\ : DFN1C0
      port map(D => \ADJ_Q[12]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[12]_net_1\);
    
    \ARB_BYTE[13]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[13]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[13]_net_1\);
    
    \ARB_WRD_40M_FIXED[3]\ : DFN1C0
      port map(D => \Q[3]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[3]_net_1\);
    
    \ARB_BYTE[7]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[7]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[7]_net_1\);
    
    \RECD_SER_WORD_RNO_0[0]\ : MX2
      port map(A => N_17, B => N_19, S => BIT_OS_SEL_3(1), Y => 
        N_33);
    
    \ARB_BYTE_RNI553D[4]\ : MX2
      port map(A => \ARB_BYTE[4]_net_1\, B => \ARB_BYTE[8]_net_1\, 
        S => BIT_OS_SEL_3(2), Y => N_21);
    
    \ARB_BYTE_RNIGQOM[6]\ : MX2
      port map(A => \ARB_BYTE[6]_net_1\, B => 
        \ARB_BYTE[10]_net_1\, S => BIT_OS_SEL_3(2), Y => N_23);
    
    \Q[4]\ : DFN1C0
      port map(D => \ADJ_Q[4]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[4]_net_1\);
    
    \ARB_WRD_40M_FIXED[7]\ : DFN1C0
      port map(D => \Q[7]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[7]_net_1\);
    
    \RECD_SER_WORD_RNO[6]\ : MX2
      port map(A => N_39, B => N_40, S => BIT_OS_SEL_4_0, Y => 
        \N_RECD_SER_WORD[6]\);
    
    \ARB_BYTE[3]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[3]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[3]_net_1\);
    
    \ARB_BYTE_RNII41F1[6]\ : MX2
      port map(A => N_23, B => N_31, S => BIT_OS_SEL_3(1), Y => 
        N_39);
    
    \ADJ_Q[5]\ : DFN1C0
      port map(D => \ADJ_Q[3]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[5]_net_1\);
    
    \ARB_BYTE[1]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[1]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[1]_net_1\);
    
    \ARB_WRD_40M_FIXED[13]\ : DFN1C0
      port map(D => \Q[13]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[13]_net_1\);
    
    \ARB_BYTE_RNIM0PM[13]\ : MX2
      port map(A => \ARB_BYTE[9]_net_1\, B => 
        \ARB_BYTE[13]_net_1\, S => BIT_OS_SEL_3(2), Y => N_32);
    
    \ADJ_Q[0]\ : DFN1C0
      port map(D => \ADJ_SER_IN_R_1DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[0]_net_1\);
    
    \ARB_WRD_40M_FIXED[10]\ : DFN1C0
      port map(D => \Q[10]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[10]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SER320M_3_34_13 is

    port( ELK_TX_DAT                 : in    std_logic_vector(7 downto 0);
          MASTER_SALT_POR_B_i_0_i_16 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_9  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_1  : in    std_logic;
          ELK_OUT_R                  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_4  : in    std_logic;
          ELK_OUT_F                  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_6  : in    std_logic;
          CCC_160M_FXD               : in    std_logic;
          CLK_40M_GL                 : in    std_logic
        );

end SER320M_3_34_13;

architecture DEF_ARCH of SER320M_3_34_13 is 

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \N_SER_CMD_WORD_R[0]\, \START_RISE\, 
        \N_SER_CMD_WORD_F[0]\, \N_SER_CMD_WORD_R[3]\, 
        \SER_CMD_WORD_R[2]_net_1\, \N_SER_CMD_WORD_R[2]\, 
        \SER_CMD_WORD_R[1]_net_1\, \N_SER_CMD_WORD_R[1]\, 
        \SER_CMD_WORD_R[0]_net_1\, \N_SER_CMD_WORD_F[3]\, 
        \SER_CMD_WORD_F[2]_net_1\, \N_SER_CMD_WORD_F[2]\, 
        \SER_CMD_WORD_F[1]_net_1\, \N_SER_CMD_WORD_F[1]\, 
        \SER_CMD_WORD_F[0]_net_1\, N_START_RISE, 
        \CLK40M_GEN_DEL0\, \SER_OUT_FI\, \SER_OUT_RI\, 
        \SER_CMD_WORD_F[3]_net_1\, \SER_CMD_WORD_R[3]_net_1\, 
        \GND\, \VCC\ : std_logic;

begin 


    SER_OUT_FI : DFN1C0
      port map(D => \SER_CMD_WORD_F[3]_net_1\, CLK => 
        CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_1, Q => 
        \SER_OUT_FI\);
    
    \SER_CMD_WORD_F[3]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[3]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_1, Q => 
        \SER_CMD_WORD_F[3]_net_1\);
    
    \SER_CMD_WORD_R[1]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[1]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_16, Q => 
        \SER_CMD_WORD_R[1]_net_1\);
    
    \SER_CMD_WORD_R[2]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[2]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_16, Q => 
        \SER_CMD_WORD_R[2]_net_1\);
    
    \SER_CMD_WORD_R_RNO[3]\ : MX2
      port map(A => \SER_CMD_WORD_R[2]_net_1\, B => ELK_TX_DAT(7), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_R[3]\);
    
    \SER_CMD_WORD_R_RNO[0]\ : NOR2B
      port map(A => \START_RISE\, B => ELK_TX_DAT(1), Y => 
        \N_SER_CMD_WORD_R[0]\);
    
    \SER_CMD_WORD_F[0]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[0]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_1, Q => 
        \SER_CMD_WORD_F[0]_net_1\);
    
    \SER_CMD_WORD_R_RNO[1]\ : MX2
      port map(A => \SER_CMD_WORD_R[0]_net_1\, B => ELK_TX_DAT(3), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_R[1]\);
    
    \SER_CMD_WORD_F_RNO[2]\ : MX2
      port map(A => \SER_CMD_WORD_F[1]_net_1\, B => ELK_TX_DAT(4), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_F[2]\);
    
    \SER_CMD_WORD_F_RNO[3]\ : MX2
      port map(A => \SER_CMD_WORD_F[2]_net_1\, B => ELK_TX_DAT(6), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_F[3]\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    CLK40M_GEN_DEL0 : DFN1C0
      port map(D => CLK_40M_GL, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_6, Q => \CLK40M_GEN_DEL0\);
    
    SER_OUT_RI : DFN1C0
      port map(D => \SER_CMD_WORD_R[3]_net_1\, CLK => 
        CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_1, Q => 
        \SER_OUT_RI\);
    
    \SER_CMD_WORD_F[2]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[2]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_1, Q => 
        \SER_CMD_WORD_F[2]_net_1\);
    
    \SER_CMD_WORD_F_RNO[1]\ : MX2
      port map(A => \SER_CMD_WORD_F[0]_net_1\, B => ELK_TX_DAT(2), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_F[1]\);
    
    \SER_CMD_WORD_R[0]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[0]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_16, Q => 
        \SER_CMD_WORD_R[0]_net_1\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    START_RISE : DFN1C0
      port map(D => N_START_RISE, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_9, Q => \START_RISE\);
    
    \SER_CMD_WORD_R[3]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[3]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_16, Q => 
        \SER_CMD_WORD_R[3]_net_1\);
    
    \SER_CMD_WORD_F_RNO[0]\ : NOR2B
      port map(A => \START_RISE\, B => ELK_TX_DAT(0), Y => 
        \N_SER_CMD_WORD_F[0]\);
    
    SER_OUT_RDEL : DFN1C0
      port map(D => \SER_OUT_RI\, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_1, Q => ELK_OUT_R);
    
    \SER_CMD_WORD_F[1]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[1]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_1, Q => 
        \SER_CMD_WORD_F[1]_net_1\);
    
    START_RISE_RNO : NOR2B
      port map(A => \CLK40M_GEN_DEL0\, B => CLK_40M_GL, Y => 
        N_START_RISE);
    
    \SER_CMD_WORD_R_RNO[2]\ : MX2
      port map(A => \SER_CMD_WORD_R[1]_net_1\, B => ELK_TX_DAT(5), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_R[2]\);
    
    SER_OUT_FDEL : DFN1C0
      port map(D => \SER_OUT_FI\, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_4, Q => ELK_OUT_F);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity DDR_BIDIR_LVDS_DUAL_CLK_13 is

    port( DCB_SALT_SEL_c_i : in    std_logic;
          ELK13_DAT_P      : inout std_logic := 'Z';
          ELK13_DAT_N      : inout std_logic := 'Z';
          ELK_OUT_R        : in    std_logic;
          ELK_OUT_F        : in    std_logic;
          CCC_160M_FXD     : in    std_logic;
          CCC_160M_ADJ     : in    std_logic;
          ELK_IN_DDR_R     : out   std_logic;
          ELK_IN_DDR_F     : out   std_logic
        );

end DDR_BIDIR_LVDS_DUAL_CLK_13;

architecture DEF_ARCH of DDR_BIDIR_LVDS_DUAL_CLK_13 is 

  component DDR_REG
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          QR  : out   std_logic;
          QF  : out   std_logic
        );
  end component;

  component DDR_OUT
    port( DR  : in    std_logic := 'U';
          DF  : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component BIBUF_LVDS
    port( PADP : inout   std_logic;
          PADN : inout   std_logic;
          D    : in    std_logic := 'U';
          E    : in    std_logic := 'U';
          Y    : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal DDR_BIDIR_LVDS_DUAL_CLK_13_GND, BIBUF_LVDS_0_Y, 
        DDR_OUT_0_Q, \VCC\ : std_logic;

begin 


    DDR_REG_0 : DDR_REG
      port map(D => BIBUF_LVDS_0_Y, CLK => CCC_160M_ADJ, CLR => 
        DDR_BIDIR_LVDS_DUAL_CLK_13_GND, QR => ELK_IN_DDR_R, QF
         => ELK_IN_DDR_F);
    
    DDR_OUT_0 : DDR_OUT
      port map(DR => ELK_OUT_R, DF => ELK_OUT_F, CLK => 
        CCC_160M_FXD, CLR => DDR_BIDIR_LVDS_DUAL_CLK_13_GND, Q
         => DDR_OUT_0_Q);
    
    BIBUF_LVDS_0 : BIBUF_LVDS
      port map(PADP => ELK13_DAT_P, PADN => ELK13_DAT_N, D => 
        DDR_OUT_0_Q, E => DCB_SALT_SEL_c_i, Y => BIBUF_LVDS_0_Y);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    GND_i : GND
      port map(Y => DDR_BIDIR_LVDS_DUAL_CLK_13_GND);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SYNC_DAT_SEL_13 is

    port( ELK_TX_DAT                : out   std_logic_vector(7 downto 0);
          PATT_ELK_DAT_13           : in    std_logic_vector(7 downto 0);
          OP_MODE_c_0               : in    std_logic;
          OP_MODE_c_6_0             : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_4 : in    std_logic;
          CLK_40M_GL                : in    std_logic
        );

end SYNC_DAT_SEL_13;

architecture DEF_ARCH of SYNC_DAT_SEL_13 is 

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \N_SERDAT[0]\, \N_SERDAT[1]\, \N_SERDAT[2]\, 
        \N_SERDAT[3]\, \N_SERDAT[4]\, \N_SERDAT[5]\, 
        \N_SERDAT[6]\, \N_SERDAT[7]\, \GND\, \VCC\ : std_logic;

begin 


    \SERDAT_RNO[4]\ : NOR2A
      port map(A => PATT_ELK_DAT_13(4), B => OP_MODE_c_0, Y => 
        \N_SERDAT[4]\);
    
    \SERDAT_RNO[0]\ : NOR2A
      port map(A => PATT_ELK_DAT_13(0), B => OP_MODE_c_6_0, Y => 
        \N_SERDAT[0]\);
    
    \SERDAT[6]\ : DFN1C0
      port map(D => \N_SERDAT[6]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_4, Q => ELK_TX_DAT(6));
    
    \SERDAT[4]\ : DFN1C0
      port map(D => \N_SERDAT[4]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_4, Q => ELK_TX_DAT(4));
    
    \SERDAT_RNO[7]\ : OR2
      port map(A => PATT_ELK_DAT_13(7), B => OP_MODE_c_0, Y => 
        \N_SERDAT[7]\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \SERDAT_RNO[3]\ : OR2
      port map(A => PATT_ELK_DAT_13(3), B => OP_MODE_c_0, Y => 
        \N_SERDAT[3]\);
    
    \SERDAT_RNO[2]\ : OR2
      port map(A => PATT_ELK_DAT_13(2), B => OP_MODE_c_0, Y => 
        \N_SERDAT[2]\);
    
    \SERDAT[5]\ : DFN1C0
      port map(D => \N_SERDAT[5]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_4, Q => ELK_TX_DAT(5));
    
    \SERDAT[7]\ : DFN1C0
      port map(D => \N_SERDAT[7]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_4, Q => ELK_TX_DAT(7));
    
    GND_i : GND
      port map(Y => \GND\);
    
    \SERDAT_RNO[5]\ : NOR2A
      port map(A => PATT_ELK_DAT_13(5), B => OP_MODE_c_0, Y => 
        \N_SERDAT[5]\);
    
    \SERDAT[0]\ : DFN1C0
      port map(D => \N_SERDAT[0]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_4, Q => ELK_TX_DAT(0));
    
    \SERDAT_RNO[6]\ : NOR2A
      port map(A => PATT_ELK_DAT_13(6), B => OP_MODE_c_0, Y => 
        \N_SERDAT[6]\);
    
    \SERDAT[1]\ : DFN1C0
      port map(D => \N_SERDAT[1]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_4, Q => ELK_TX_DAT(1));
    
    \SERDAT_RNO[1]\ : OR2
      port map(A => PATT_ELK_DAT_13(1), B => OP_MODE_c_0, Y => 
        \N_SERDAT[1]\);
    
    \SERDAT[3]\ : DFN1C0
      port map(D => \N_SERDAT[3]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_4, Q => ELK_TX_DAT(3));
    
    \SERDAT[2]\ : DFN1C0
      port map(D => \N_SERDAT[2]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_4, Q => ELK_TX_DAT(2));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity ELINK_SLAVE_15_8 is

    port( BIT_OS_SEL_2_0             : in    std_logic;
          BIT_OS_SEL_3               : in    std_logic_vector(2 downto 1);
          BIT_OS_SEL_6_0             : in    std_logic;
          BIT_OS_SEL_5_0             : in    std_logic;
          BIT_OS_SEL_4_0             : in    std_logic;
          ELK_RX_SER_WORD_13         : out   std_logic_vector(7 downto 0);
          OP_MODE_c_6_0              : in    std_logic;
          OP_MODE_c_0                : in    std_logic;
          PATT_ELK_DAT_13            : in    std_logic_vector(7 downto 0);
          MASTER_DCB_POR_B_i_0_i     : in    std_logic;
          ELK13_DAT_N                : inout std_logic := 'Z';
          ELK13_DAT_P                : inout std_logic := 'Z';
          DCB_SALT_SEL_c_i           : in    std_logic;
          CCC_160M_FXD               : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_6  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_1  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_9  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_16 : in    std_logic;
          CLK_40M_GL                 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_4  : in    std_logic;
          DEV_RST_B_c                : in    std_logic;
          CCC_160M_ADJ               : in    std_logic
        );

end ELINK_SLAVE_15_8;

architecture DEF_ARCH of ELINK_SLAVE_15_8 is 

  component SLAVE_DES320S_1_17_11
    port( ELK_RX_SER_WORD_13     : out   std_logic_vector(7 downto 0);
          BIT_OS_SEL_4_0         : in    std_logic := 'U';
          BIT_OS_SEL_5_0         : in    std_logic := 'U';
          BIT_OS_SEL_6_0         : in    std_logic := 'U';
          BIT_OS_SEL_3           : in    std_logic_vector(2 downto 1) := (others => 'U');
          BIT_OS_SEL_2_0         : in    std_logic := 'U';
          CLK_40M_GL             : in    std_logic := 'U';
          CCC_160M_FXD           : in    std_logic := 'U';
          ELK_IN_R               : in    std_logic := 'U';
          ELK_IN_F               : in    std_logic := 'U';
          MASTER_DCB_POR_B_i_0_i : in    std_logic := 'U';
          CCC_160M_ADJ           : in    std_logic := 'U'
        );
  end component;

  component SER320M_3_34_13
    port( ELK_TX_DAT                 : in    std_logic_vector(7 downto 0) := (others => 'U');
          MASTER_SALT_POR_B_i_0_i_16 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_9  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_1  : in    std_logic := 'U';
          ELK_OUT_R                  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_4  : in    std_logic := 'U';
          ELK_OUT_F                  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_6  : in    std_logic := 'U';
          CCC_160M_FXD               : in    std_logic := 'U';
          CLK_40M_GL                 : in    std_logic := 'U'
        );
  end component;

  component DDR_BIDIR_LVDS_DUAL_CLK_13
    port( DCB_SALT_SEL_c_i : in    std_logic := 'U';
          ELK13_DAT_P      : inout   std_logic;
          ELK13_DAT_N      : inout   std_logic;
          ELK_OUT_R        : in    std_logic := 'U';
          ELK_OUT_F        : in    std_logic := 'U';
          CCC_160M_FXD     : in    std_logic := 'U';
          CCC_160M_ADJ     : in    std_logic := 'U';
          ELK_IN_DDR_R     : out   std_logic;
          ELK_IN_DDR_F     : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component SYNC_DAT_SEL_13
    port( ELK_TX_DAT                : out   std_logic_vector(7 downto 0);
          PATT_ELK_DAT_13           : in    std_logic_vector(7 downto 0) := (others => 'U');
          OP_MODE_c_0               : in    std_logic := 'U';
          OP_MODE_c_6_0             : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_4 : in    std_logic := 'U';
          CLK_40M_GL                : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \ELK_IN_F\, ELK_IN_DDR_F, \ELK_IN_R\, ELK_IN_DDR_R, 
        \ELK_TX_DAT[0]\, \ELK_TX_DAT[1]\, \ELK_TX_DAT[2]\, 
        \ELK_TX_DAT[3]\, \ELK_TX_DAT[4]\, \ELK_TX_DAT[5]\, 
        \ELK_TX_DAT[6]\, \ELK_TX_DAT[7]\, ELK_OUT_R, ELK_OUT_F, 
        \GND\, \VCC\ : std_logic;

    for all : SLAVE_DES320S_1_17_11
	Use entity work.SLAVE_DES320S_1_17_11(DEF_ARCH);
    for all : SER320M_3_34_13
	Use entity work.SER320M_3_34_13(DEF_ARCH);
    for all : DDR_BIDIR_LVDS_DUAL_CLK_13
	Use entity work.DDR_BIDIR_LVDS_DUAL_CLK_13(DEF_ARCH);
    for all : SYNC_DAT_SEL_13
	Use entity work.SYNC_DAT_SEL_13(DEF_ARCH);
begin 


    U_SLAVE_1ELK : SLAVE_DES320S_1_17_11
      port map(ELK_RX_SER_WORD_13(7) => ELK_RX_SER_WORD_13(7), 
        ELK_RX_SER_WORD_13(6) => ELK_RX_SER_WORD_13(6), 
        ELK_RX_SER_WORD_13(5) => ELK_RX_SER_WORD_13(5), 
        ELK_RX_SER_WORD_13(4) => ELK_RX_SER_WORD_13(4), 
        ELK_RX_SER_WORD_13(3) => ELK_RX_SER_WORD_13(3), 
        ELK_RX_SER_WORD_13(2) => ELK_RX_SER_WORD_13(2), 
        ELK_RX_SER_WORD_13(1) => ELK_RX_SER_WORD_13(1), 
        ELK_RX_SER_WORD_13(0) => ELK_RX_SER_WORD_13(0), 
        BIT_OS_SEL_4_0 => BIT_OS_SEL_4_0, BIT_OS_SEL_5_0 => 
        BIT_OS_SEL_5_0, BIT_OS_SEL_6_0 => BIT_OS_SEL_6_0, 
        BIT_OS_SEL_3(2) => BIT_OS_SEL_3(2), BIT_OS_SEL_3(1) => 
        BIT_OS_SEL_3(1), BIT_OS_SEL_2_0 => BIT_OS_SEL_2_0, 
        CLK_40M_GL => CLK_40M_GL, CCC_160M_FXD => CCC_160M_FXD, 
        ELK_IN_R => \ELK_IN_R\, ELK_IN_F => \ELK_IN_F\, 
        MASTER_DCB_POR_B_i_0_i => MASTER_DCB_POR_B_i_0_i, 
        CCC_160M_ADJ => CCC_160M_ADJ);
    
    U_ELK1_CMD_TX : SER320M_3_34_13
      port map(ELK_TX_DAT(7) => \ELK_TX_DAT[7]\, ELK_TX_DAT(6)
         => \ELK_TX_DAT[6]\, ELK_TX_DAT(5) => \ELK_TX_DAT[5]\, 
        ELK_TX_DAT(4) => \ELK_TX_DAT[4]\, ELK_TX_DAT(3) => 
        \ELK_TX_DAT[3]\, ELK_TX_DAT(2) => \ELK_TX_DAT[2]\, 
        ELK_TX_DAT(1) => \ELK_TX_DAT[1]\, ELK_TX_DAT(0) => 
        \ELK_TX_DAT[0]\, MASTER_SALT_POR_B_i_0_i_16 => 
        MASTER_SALT_POR_B_i_0_i_16, MASTER_SALT_POR_B_i_0_i_9 => 
        MASTER_SALT_POR_B_i_0_i_9, MASTER_SALT_POR_B_i_0_i_1 => 
        MASTER_SALT_POR_B_i_0_i_1, ELK_OUT_R => ELK_OUT_R, 
        MASTER_SALT_POR_B_i_0_i_4 => MASTER_SALT_POR_B_i_0_i_4, 
        ELK_OUT_F => ELK_OUT_F, MASTER_SALT_POR_B_i_0_i_6 => 
        MASTER_SALT_POR_B_i_0_i_6, CCC_160M_FXD => CCC_160M_FXD, 
        CLK_40M_GL => CLK_40M_GL);
    
    U_DDR_ELK1 : DDR_BIDIR_LVDS_DUAL_CLK_13
      port map(DCB_SALT_SEL_c_i => DCB_SALT_SEL_c_i, ELK13_DAT_P
         => ELK13_DAT_P, ELK13_DAT_N => ELK13_DAT_N, ELK_OUT_R
         => ELK_OUT_R, ELK_OUT_F => ELK_OUT_F, CCC_160M_FXD => 
        CCC_160M_FXD, CCC_160M_ADJ => CCC_160M_ADJ, ELK_IN_DDR_R
         => ELK_IN_DDR_R, ELK_IN_DDR_F => ELK_IN_DDR_F);
    
    ELK_IN_F : DFN1C0
      port map(D => ELK_IN_DDR_F, CLK => CCC_160M_ADJ, CLR => 
        DEV_RST_B_c, Q => \ELK_IN_F\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    U_ELK1_SERDAT_SOURCE : SYNC_DAT_SEL_13
      port map(ELK_TX_DAT(7) => \ELK_TX_DAT[7]\, ELK_TX_DAT(6)
         => \ELK_TX_DAT[6]\, ELK_TX_DAT(5) => \ELK_TX_DAT[5]\, 
        ELK_TX_DAT(4) => \ELK_TX_DAT[4]\, ELK_TX_DAT(3) => 
        \ELK_TX_DAT[3]\, ELK_TX_DAT(2) => \ELK_TX_DAT[2]\, 
        ELK_TX_DAT(1) => \ELK_TX_DAT[1]\, ELK_TX_DAT(0) => 
        \ELK_TX_DAT[0]\, PATT_ELK_DAT_13(7) => PATT_ELK_DAT_13(7), 
        PATT_ELK_DAT_13(6) => PATT_ELK_DAT_13(6), 
        PATT_ELK_DAT_13(5) => PATT_ELK_DAT_13(5), 
        PATT_ELK_DAT_13(4) => PATT_ELK_DAT_13(4), 
        PATT_ELK_DAT_13(3) => PATT_ELK_DAT_13(3), 
        PATT_ELK_DAT_13(2) => PATT_ELK_DAT_13(2), 
        PATT_ELK_DAT_13(1) => PATT_ELK_DAT_13(1), 
        PATT_ELK_DAT_13(0) => PATT_ELK_DAT_13(0), OP_MODE_c_0 => 
        OP_MODE_c_0, OP_MODE_c_6_0 => OP_MODE_c_6_0, 
        MASTER_SALT_POR_B_i_0_i_4 => MASTER_SALT_POR_B_i_0_i_4, 
        CLK_40M_GL => CLK_40M_GL);
    
    ELK_IN_R : DFN1C0
      port map(D => ELK_IN_DDR_R, CLK => CCC_160M_ADJ, CLR => 
        DEV_RST_B_c, Q => \ELK_IN_R\);
    
    GND_i : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SYNC_DAT_SEL_0 is

    port( ELK0_TX_DAT                : out   std_logic_vector(7 downto 0);
          PATT_ELK_DAT_0             : in    std_logic_vector(7 downto 0);
          OP_MODE_c_4_0              : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_10 : in    std_logic;
          CLK_40M_GL                 : in    std_logic
        );

end SYNC_DAT_SEL_0;

architecture DEF_ARCH of SYNC_DAT_SEL_0 is 

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \N_SERDAT[0]\, \N_SERDAT[1]\, \N_SERDAT[2]\, 
        \N_SERDAT[3]\, \N_SERDAT[4]\, \N_SERDAT[5]\, 
        \N_SERDAT[6]\, \N_SERDAT[7]\, \GND\, \VCC\ : std_logic;

begin 


    \SERDAT_RNO[4]\ : NOR2A
      port map(A => PATT_ELK_DAT_0(4), B => OP_MODE_c_4_0, Y => 
        \N_SERDAT[4]\);
    
    \SERDAT_RNO[0]\ : NOR2A
      port map(A => PATT_ELK_DAT_0(0), B => OP_MODE_c_4_0, Y => 
        \N_SERDAT[0]\);
    
    \SERDAT[6]\ : DFN1C0
      port map(D => \N_SERDAT[6]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_10, Q => ELK0_TX_DAT(6));
    
    \SERDAT[4]\ : DFN1C0
      port map(D => \N_SERDAT[4]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_10, Q => ELK0_TX_DAT(4));
    
    \SERDAT_RNO[7]\ : OR2
      port map(A => PATT_ELK_DAT_0(7), B => OP_MODE_c_4_0, Y => 
        \N_SERDAT[7]\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \SERDAT_RNO[3]\ : OR2
      port map(A => PATT_ELK_DAT_0(3), B => OP_MODE_c_4_0, Y => 
        \N_SERDAT[3]\);
    
    \SERDAT_RNO[2]\ : OR2
      port map(A => PATT_ELK_DAT_0(2), B => OP_MODE_c_4_0, Y => 
        \N_SERDAT[2]\);
    
    \SERDAT[5]\ : DFN1C0
      port map(D => \N_SERDAT[5]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_10, Q => ELK0_TX_DAT(5));
    
    \SERDAT[7]\ : DFN1C0
      port map(D => \N_SERDAT[7]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_10, Q => ELK0_TX_DAT(7));
    
    GND_i : GND
      port map(Y => \GND\);
    
    \SERDAT_RNO[5]\ : NOR2A
      port map(A => PATT_ELK_DAT_0(5), B => OP_MODE_c_4_0, Y => 
        \N_SERDAT[5]\);
    
    \SERDAT[0]\ : DFN1C0
      port map(D => \N_SERDAT[0]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_10, Q => ELK0_TX_DAT(0));
    
    \SERDAT_RNO[6]\ : NOR2A
      port map(A => PATT_ELK_DAT_0(6), B => OP_MODE_c_4_0, Y => 
        \N_SERDAT[6]\);
    
    \SERDAT[1]\ : DFN1C0
      port map(D => \N_SERDAT[1]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_10, Q => ELK0_TX_DAT(1));
    
    \SERDAT_RNO[1]\ : OR2
      port map(A => PATT_ELK_DAT_0(1), B => OP_MODE_c_4_0, Y => 
        \N_SERDAT[1]\);
    
    \SERDAT[3]\ : DFN1C0
      port map(D => \N_SERDAT[3]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_10, Q => ELK0_TX_DAT(3));
    
    \SERDAT[2]\ : DFN1C0
      port map(D => \N_SERDAT[2]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_10, Q => ELK0_TX_DAT(2));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity USB_EXEC is

    port( P_MASTER_POR_B_c_24    : in    std_logic;
          P_MASTER_POR_B_c_28    : in    std_logic;
          P_MASTER_POR_B_c_27    : in    std_logic;
          P_MASTER_POR_B_c_34_0  : in    std_logic;
          P_USB_MASTER_EN_c      : out   std_logic;
          P_MASTER_POR_B_c_29    : in    std_logic;
          P_MASTER_POR_B_c_32_0  : in    std_logic;
          CLK_40M_GL             : in    std_logic;
          P_MASTER_POR_B_c_23    : in    std_logic;
          P_USB_MASTER_EN_c_0    : out   std_logic;
          P_USB_MASTER_EN_c_1    : out   std_logic;
          P_USB_MASTER_EN_c_2    : out   std_logic;
          P_USB_MASTER_EN_c_3    : out   std_logic;
          P_USB_MASTER_EN_c_4    : out   std_logic;
          P_USB_MASTER_EN_c_5    : out   std_logic;
          P_USB_MASTER_EN_c_6    : out   std_logic;
          P_USB_MASTER_EN_c_7    : out   std_logic;
          P_USB_MASTER_EN_c_8    : out   std_logic;
          P_USB_MASTER_EN_c_9    : out   std_logic;
          P_USB_MASTER_EN_c_10   : out   std_logic;
          P_USB_MASTER_EN_c_11   : out   std_logic;
          P_USB_MASTER_EN_c_12   : out   std_logic;
          P_USB_MASTER_EN_c_13   : out   std_logic;
          P_USB_MASTER_EN_c_14   : out   std_logic;
          P_USB_MASTER_EN_c_15   : out   std_logic;
          P_USB_MASTER_EN_c_16   : out   std_logic;
          P_USB_MASTER_EN_c_17   : out   std_logic;
          P_USB_MASTER_EN_c_18   : out   std_logic;
          P_USB_MASTER_EN_c_19   : out   std_logic;
          P_USB_MASTER_EN_c_20   : out   std_logic;
          P_USB_MASTER_EN_c_21   : out   std_logic;
          P_MASTER_POR_B_c_0     : in    std_logic;
          P_USB_MASTER_EN_c_22   : out   std_logic;
          P_USB_MASTER_EN_c_22_0 : out   std_logic;
          P_USB_MASTER_EN_c_2_0  : out   std_logic;
          P_MASTER_POR_B_c_0_0   : in    std_logic;
          P_USB_MASTER_EN_c_1_0  : out   std_logic;
          P_MASTER_POR_B_c_22_0  : in    std_logic;
          CLK60MHZ               : in    std_logic
        );

end USB_EXEC;

architecture DEF_ARCH of USB_EXEC is 

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component MX2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component DFN1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OA1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component AO1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \USB_EN_60M_1S_0\, \USB_EN_60M_S\, \USB_EN_60M_1S\, 
        T_CNT60M_18_0, \T_CNT60M[6]_net_1\, T_CNT60M_c5, 
        un8_cnt_en_60m2s_2, \T_CNT60M[4]_net_1\, 
        \T_CNT60M[7]_net_1\, un8_cnt_en_60m2s_1, 
        \T_CNT60M[5]_net_1\, N_T_CNT60M_0_sqmuxa, T_CNT60M_c3, 
        \CNT_EN_60M2S\, N_T_CNT60M_1_sqmuxa, N_49, 
        \T_CNT60M[1]_net_1\, N_51, \T_CNT60M[2]_net_1\, 
        T_CNT60M_c2, T_CNT60M_c1, N_53, \T_CNT60M[3]_net_1\, N_55, 
        T_CNT60M_c4, N_57, N_59, N_61, T_CNT60M_n0, 
        \T_CNT60M[0]_net_1\, T_CNT60M_n1, T_CNT60M_n2, 
        T_CNT60M_n3, T_CNT60M_n4, T_CNT60M_n5, T_CNT60M_n6, 
        T_CNT60M_n7, \TEST_SM_RNO[3]_net_1\, \TEST_SM_i_0[2]\, 
        \TEST_SM[3]_net_1\, \TERMCNT_FG40M2S\, 
        \TEST_SM_RNO[2]_net_1\, \TEST_SM[1]_net_1\, 
        \TEST_SM_ns[1]\, \TEST_SM[0]_net_1\, N_CNT_EN_40M, 
        \TEST_SM_ns[4]\, \TEST_SM[4]_net_1\, \CNT_EN_60M1S\, 
        \CNT_EN_60M0S\, \TERMCNT_FG40M0S\, \TERMCNT_FG60M\, 
        \TERMCNT_FG40M1S\, \USB_EN_40M\, \CNT_EN_40M\, 
        USB_EXEC_GND, \VCC\ : std_logic;

begin 


    \T_CNT60M_RNIVI6H[5]\ : NOR2B
      port map(A => \T_CNT60M[5]_net_1\, B => \T_CNT60M[6]_net_1\, 
        Y => un8_cnt_en_60m2s_1);
    
    \TEST_SM_RNO[4]\ : AO1
      port map(A => \TERMCNT_FG40M2S\, B => \TEST_SM[3]_net_1\, C
         => \TEST_SM[4]_net_1\, Y => \TEST_SM_ns[4]\);
    
    \TEST_SM_RNO[2]\ : AO1C
      port map(A => \TEST_SM[1]_net_1\, B => \TEST_SM_i_0[2]\, C
         => \TERMCNT_FG40M2S\, Y => \TEST_SM_RNO[2]_net_1\);
    
    \T_CNT60M_RNO_0[1]\ : MX2
      port map(A => \CNT_EN_60M2S\, B => \T_CNT60M[1]_net_1\, S
         => N_T_CNT60M_1_sqmuxa, Y => N_49);
    
    \T_CNT60M_RNO[2]\ : AX1C
      port map(A => N_T_CNT60M_1_sqmuxa, B => T_CNT60M_c1, C => 
        N_51, Y => T_CNT60M_n2);
    
    CNT_EN_60M2S_RNI1R172 : AOI1B
      port map(A => un8_cnt_en_60m2s_2, B => T_CNT60M_c3, C => 
        \CNT_EN_60M2S\, Y => N_T_CNT60M_1_sqmuxa);
    
    \T_CNT60M_RNO_0[7]\ : NOR2B
      port map(A => \T_CNT60M[6]_net_1\, B => T_CNT60M_c5, Y => 
        T_CNT60M_18_0);
    
    \T_CNT60M[5]\ : DFN1C0
      port map(D => T_CNT60M_n5, CLK => CLK60MHZ, CLR => 
        P_MASTER_POR_B_c_28, Q => \T_CNT60M[5]_net_1\);
    
    USB_EN_60M_2S_13 : DFN1C0
      port map(D => \USB_EN_60M_1S_0\, CLK => CLK60MHZ, CLR => 
        P_MASTER_POR_B_c_0, Q => P_USB_MASTER_EN_c_13);
    
    \TEST_SM_RNO[1]\ : MX2B
      port map(A => \TEST_SM[0]_net_1\, B => \TERMCNT_FG40M2S\, S
         => \TEST_SM[1]_net_1\, Y => \TEST_SM_ns[1]\);
    
    CNT_EN_40M : DFN1C0
      port map(D => N_CNT_EN_40M, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_23, Q => \CNT_EN_40M\);
    
    \T_CNT60M_RNIL86H[1]\ : NOR2B
      port map(A => \T_CNT60M[1]_net_1\, B => \T_CNT60M[0]_net_1\, 
        Y => T_CNT60M_c1);
    
    \T_CNT60M_RNO_0[6]\ : MX2
      port map(A => \CNT_EN_60M2S\, B => \T_CNT60M[6]_net_1\, S
         => N_T_CNT60M_1_sqmuxa, Y => N_59);
    
    TERMCNT_FG60M : DFN1C0
      port map(D => N_T_CNT60M_0_sqmuxa, CLK => CLK60MHZ, CLR => 
        P_MASTER_POR_B_c_27, Q => \TERMCNT_FG60M\);
    
    \T_CNT60M_RNO_0[4]\ : MX2
      port map(A => \CNT_EN_60M2S\, B => \T_CNT60M[4]_net_1\, S
         => N_T_CNT60M_1_sqmuxa, Y => N_55);
    
    USB_EN_60M_2S_8 : DFN1C0
      port map(D => \USB_EN_60M_1S\, CLK => CLK60MHZ, CLR => 
        P_MASTER_POR_B_c_0_0, Q => P_USB_MASTER_EN_c_8);
    
    USB_EN_60M_2S_17 : DFN1C0
      port map(D => \USB_EN_60M_1S_0\, CLK => CLK60MHZ, CLR => 
        P_MASTER_POR_B_c_0, Q => P_USB_MASTER_EN_c_17);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    USB_EN_60M_2S_7 : DFN1C0
      port map(D => \USB_EN_60M_1S\, CLK => CLK60MHZ, CLR => 
        P_MASTER_POR_B_c_0_0, Q => P_USB_MASTER_EN_c_7);
    
    USB_EN_60M_2S_16 : DFN1C0
      port map(D => \USB_EN_60M_1S_0\, CLK => CLK60MHZ, CLR => 
        P_MASTER_POR_B_c_0, Q => P_USB_MASTER_EN_c_16);
    
    CNT_EN_60M0S : DFN1C0
      port map(D => \CNT_EN_40M\, CLK => CLK60MHZ, CLR => 
        P_MASTER_POR_B_c_23, Q => \CNT_EN_60M0S\);
    
    USB_EN_60M_2S_18 : DFN1C0
      port map(D => \USB_EN_60M_1S_0\, CLK => CLK60MHZ, CLR => 
        P_MASTER_POR_B_c_0, Q => P_USB_MASTER_EN_c_18);
    
    \T_CNT60M_RNO[5]\ : AX1C
      port map(A => N_T_CNT60M_1_sqmuxa, B => T_CNT60M_c4, C => 
        N_57, Y => T_CNT60M_n5);
    
    \T_CNT60M_RNO[4]\ : AX1C
      port map(A => N_T_CNT60M_1_sqmuxa, B => T_CNT60M_c3, C => 
        N_55, Y => T_CNT60M_n4);
    
    USB_EN_60M_2S_2 : DFN1C0
      port map(D => \USB_EN_60M_1S\, CLK => CLK60MHZ, CLR => 
        P_MASTER_POR_B_c_0_0, Q => P_USB_MASTER_EN_c_2);
    
    \T_CNT60M[1]\ : DFN1C0
      port map(D => T_CNT60M_n1, CLK => CLK60MHZ, CLR => 
        P_MASTER_POR_B_c_28, Q => \T_CNT60M[1]_net_1\);
    
    USB_EN_60M_2S_6 : DFN1C0
      port map(D => \USB_EN_60M_1S\, CLK => CLK60MHZ, CLR => 
        P_MASTER_POR_B_c_0_0, Q => P_USB_MASTER_EN_c_6);
    
    USB_EN_60M_2S_1_0 : DFN1C0
      port map(D => \USB_EN_60M_1S_0\, CLK => CLK60MHZ, CLR => 
        P_MASTER_POR_B_c_0_0, Q => P_USB_MASTER_EN_c_1_0);
    
    \T_CNT60M[7]\ : DFN1C0
      port map(D => T_CNT60M_n7, CLK => CLK60MHZ, CLR => 
        P_MASTER_POR_B_c_29, Q => \T_CNT60M[7]_net_1\);
    
    TERMCNT_FG40M1S : DFN1C0
      port map(D => \TERMCNT_FG40M0S\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_32_0, Q => \TERMCNT_FG40M1S\);
    
    USB_EN_60M_2S_10 : DFN1C0
      port map(D => \USB_EN_60M_1S\, CLK => CLK60MHZ, CLR => 
        P_MASTER_POR_B_c_0, Q => P_USB_MASTER_EN_c_10);
    
    \T_CNT60M_RNO_1[7]\ : MX2
      port map(A => \CNT_EN_60M2S\, B => \T_CNT60M[7]_net_1\, S
         => N_T_CNT60M_1_sqmuxa, Y => N_61);
    
    \T_CNT60M_RNO[0]\ : MX2B
      port map(A => \CNT_EN_60M2S\, B => \T_CNT60M[0]_net_1\, S
         => N_T_CNT60M_1_sqmuxa, Y => T_CNT60M_n0);
    
    \T_CNT60M_RNIELC21[3]\ : NOR2B
      port map(A => \T_CNT60M[3]_net_1\, B => T_CNT60M_c2, Y => 
        T_CNT60M_c3);
    
    \TEST_SM[1]\ : DFN1C0
      port map(D => \TEST_SM_ns[1]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_24, Q => \TEST_SM[1]_net_1\);
    
    USB_EN_60M_2S_19 : DFN1C0
      port map(D => \USB_EN_60M_1S_0\, CLK => CLK60MHZ, CLR => 
        P_MASTER_POR_B_c_0, Q => P_USB_MASTER_EN_c_19);
    
    \T_CNT60M_RNO_0[3]\ : MX2
      port map(A => \CNT_EN_60M2S\, B => \T_CNT60M[3]_net_1\, S
         => N_T_CNT60M_1_sqmuxa, Y => N_53);
    
    \T_CNT60M_RNIB6JJ1[5]\ : NOR2B
      port map(A => T_CNT60M_c4, B => \T_CNT60M[5]_net_1\, Y => 
        T_CNT60M_c5);
    
    \T_CNT60M[6]\ : DFN1C0
      port map(D => T_CNT60M_n6, CLK => CLK60MHZ, CLR => 
        P_MASTER_POR_B_c_28, Q => \T_CNT60M[6]_net_1\);
    
    \TEST_SM[0]\ : DFN1P0
      port map(D => USB_EXEC_GND, CLK => CLK_40M_GL, PRE => 
        P_MASTER_POR_B_c_24, Q => \TEST_SM[0]_net_1\);
    
    USB_EN_60M_2S_22 : DFN1C0
      port map(D => \USB_EN_60M_1S_0\, CLK => CLK60MHZ, CLR => 
        P_MASTER_POR_B_c_0, Q => P_USB_MASTER_EN_c_22);
    
    \TEST_SM_RNO[3]\ : OA1C
      port map(A => \TEST_SM_i_0[2]\, B => \TEST_SM[3]_net_1\, C
         => \TERMCNT_FG40M2S\, Y => \TEST_SM_RNO[3]_net_1\);
    
    \T_CNT60M[2]\ : DFN1C0
      port map(D => T_CNT60M_n2, CLK => CLK60MHZ, CLR => 
        P_MASTER_POR_B_c_28, Q => \T_CNT60M[2]_net_1\);
    
    USB_EN_40M : DFN1C0
      port map(D => \TEST_SM[4]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_29, Q => \USB_EN_40M\);
    
    USB_EN_60M_2S_22_0 : DFN1C0
      port map(D => \USB_EN_60M_1S_0\, CLK => CLK60MHZ, CLR => 
        P_MASTER_POR_B_c_0_0, Q => P_USB_MASTER_EN_c_22_0);
    
    USB_EN_60M_1S : DFN1C0
      port map(D => \USB_EN_60M_S\, CLK => CLK60MHZ, CLR => 
        P_MASTER_POR_B_c_22_0, Q => \USB_EN_60M_1S\);
    
    \T_CNT60M_RNO[6]\ : AX1C
      port map(A => N_T_CNT60M_1_sqmuxa, B => T_CNT60M_c5, C => 
        N_59, Y => T_CNT60M_n6);
    
    \T_CNT60M_RNO[3]\ : AX1C
      port map(A => N_T_CNT60M_1_sqmuxa, B => T_CNT60M_c2, C => 
        N_53, Y => T_CNT60M_n3);
    
    USB_EN_60M_2S_21 : DFN1C0
      port map(D => \USB_EN_60M_1S_0\, CLK => CLK60MHZ, CLR => 
        P_MASTER_POR_B_c_0, Q => P_USB_MASTER_EN_c_21);
    
    USB_EN_60M_2S_3 : DFN1C0
      port map(D => \USB_EN_60M_1S\, CLK => CLK60MHZ, CLR => 
        P_MASTER_POR_B_c_0_0, Q => P_USB_MASTER_EN_c_3);
    
    \T_CNT60M[4]\ : DFN1C0
      port map(D => T_CNT60M_n4, CLK => CLK60MHZ, CLR => 
        P_MASTER_POR_B_c_28, Q => \T_CNT60M[4]_net_1\);
    
    GND_i : GND
      port map(Y => USB_EXEC_GND);
    
    TERMCNT_FG40M0S : DFN1C0
      port map(D => \TERMCNT_FG60M\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_32_0, Q => \TERMCNT_FG40M0S\);
    
    USB_EN_60M_2S_9 : DFN1C0
      port map(D => \USB_EN_60M_1S\, CLK => CLK60MHZ, CLR => 
        P_MASTER_POR_B_c_0_0, Q => P_USB_MASTER_EN_c_9);
    
    USB_EN_60M_2S_0 : DFN1C0
      port map(D => \USB_EN_60M_1S\, CLK => CLK60MHZ, CLR => 
        P_MASTER_POR_B_c_0_0, Q => P_USB_MASTER_EN_c_0);
    
    \T_CNT60M_RNICTVA1[4]\ : NOR2B
      port map(A => \T_CNT60M[4]_net_1\, B => T_CNT60M_c3, Y => 
        T_CNT60M_c4);
    
    CNT_EN_40M_RNO : AO1A
      port map(A => \TERMCNT_FG40M2S\, B => \TEST_SM[1]_net_1\, C
         => \TEST_SM[3]_net_1\, Y => N_CNT_EN_40M);
    
    USB_EN_60M_2S_15 : DFN1C0
      port map(D => \USB_EN_60M_1S_0\, CLK => CLK60MHZ, CLR => 
        P_MASTER_POR_B_c_0, Q => P_USB_MASTER_EN_c_15);
    
    \TEST_SM[2]\ : DFN1P0
      port map(D => \TEST_SM_RNO[2]_net_1\, CLK => CLK_40M_GL, 
        PRE => P_MASTER_POR_B_c_24, Q => \TEST_SM_i_0[2]\);
    
    USB_EN_60M_2S_5 : DFN1C0
      port map(D => \USB_EN_60M_1S\, CLK => CLK60MHZ, CLR => 
        P_MASTER_POR_B_c_0_0, Q => P_USB_MASTER_EN_c_5);
    
    \T_CNT60M_RNO_0[2]\ : MX2
      port map(A => \CNT_EN_60M2S\, B => \T_CNT60M[2]_net_1\, S
         => N_T_CNT60M_1_sqmuxa, Y => N_51);
    
    \TEST_SM[3]\ : DFN1C0
      port map(D => \TEST_SM_RNO[3]_net_1\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_24, Q => \TEST_SM[3]_net_1\);
    
    TERMCNT_FG60M_RNO : NOR3C
      port map(A => T_CNT60M_c3, B => un8_cnt_en_60m2s_2, C => 
        \CNT_EN_60M2S\, Y => N_T_CNT60M_0_sqmuxa);
    
    USB_EN_60M_S : DFN1C0
      port map(D => \USB_EN_40M\, CLK => CLK60MHZ, CLR => 
        P_MASTER_POR_B_c_34_0, Q => \USB_EN_60M_S\);
    
    USB_EN_60M_2S_1 : DFN1C0
      port map(D => \USB_EN_60M_1S\, CLK => CLK60MHZ, CLR => 
        P_MASTER_POR_B_c_0_0, Q => P_USB_MASTER_EN_c_1);
    
    USB_EN_60M_1S_0 : DFN1C0
      port map(D => \USB_EN_60M_S\, CLK => CLK60MHZ, CLR => 
        P_MASTER_POR_B_c_22_0, Q => \USB_EN_60M_1S_0\);
    
    CNT_EN_60M2S : DFN1C0
      port map(D => \CNT_EN_60M1S\, CLK => CLK60MHZ, CLR => 
        P_MASTER_POR_B_c_23, Q => \CNT_EN_60M2S\);
    
    \TEST_SM[4]\ : DFN1C0
      port map(D => \TEST_SM_ns[4]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_24, Q => \TEST_SM[4]_net_1\);
    
    USB_EN_60M_2S_4 : DFN1C0
      port map(D => \USB_EN_60M_1S\, CLK => CLK60MHZ, CLR => 
        P_MASTER_POR_B_c_0_0, Q => P_USB_MASTER_EN_c_4);
    
    USB_EN_60M_2S_2_0 : DFN1C0
      port map(D => \USB_EN_60M_1S_0\, CLK => CLK60MHZ, CLR => 
        P_MASTER_POR_B_c_0_0, Q => P_USB_MASTER_EN_c_2_0);
    
    \T_CNT60M_RNO[1]\ : AX1C
      port map(A => N_T_CNT60M_1_sqmuxa, B => \T_CNT60M[0]_net_1\, 
        C => N_49, Y => T_CNT60M_n1);
    
    \T_CNT60M_RNO_0[5]\ : MX2
      port map(A => \CNT_EN_60M2S\, B => \T_CNT60M[5]_net_1\, S
         => N_T_CNT60M_1_sqmuxa, Y => N_57);
    
    TERMCNT_FG40M2S : DFN1C0
      port map(D => \TERMCNT_FG40M1S\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_32_0, Q => \TERMCNT_FG40M2S\);
    
    USB_EN_60M_2S_12 : DFN1C0
      port map(D => \USB_EN_60M_1S_0\, CLK => CLK60MHZ, CLR => 
        P_MASTER_POR_B_c_0, Q => P_USB_MASTER_EN_c_12);
    
    \T_CNT60M_RNO[7]\ : AX1C
      port map(A => N_T_CNT60M_1_sqmuxa, B => T_CNT60M_18_0, C
         => N_61, Y => T_CNT60M_n7);
    
    \T_CNT60M[0]\ : DFN1C0
      port map(D => T_CNT60M_n0, CLK => CLK60MHZ, CLR => 
        P_MASTER_POR_B_c_28, Q => \T_CNT60M[0]_net_1\);
    
    USB_EN_60M_2S_14 : DFN1C0
      port map(D => \USB_EN_60M_1S_0\, CLK => CLK60MHZ, CLR => 
        P_MASTER_POR_B_c_0, Q => P_USB_MASTER_EN_c_14);
    
    USB_EN_60M_2S_11 : DFN1C0
      port map(D => \USB_EN_60M_1S\, CLK => CLK60MHZ, CLR => 
        P_MASTER_POR_B_c_0, Q => P_USB_MASTER_EN_c_11);
    
    \T_CNT60M_RNIHEPP[2]\ : NOR2B
      port map(A => \T_CNT60M[2]_net_1\, B => T_CNT60M_c1, Y => 
        T_CNT60M_c2);
    
    \T_CNT60M_RNIU5D21[7]\ : NOR3C
      port map(A => \T_CNT60M[4]_net_1\, B => \T_CNT60M[7]_net_1\, 
        C => un8_cnt_en_60m2s_1, Y => un8_cnt_en_60m2s_2);
    
    CNT_EN_60M1S : DFN1C0
      port map(D => \CNT_EN_60M0S\, CLK => CLK60MHZ, CLR => 
        P_MASTER_POR_B_c_23, Q => \CNT_EN_60M1S\);
    
    USB_EN_60M_2S_20 : DFN1C0
      port map(D => \USB_EN_60M_1S_0\, CLK => CLK60MHZ, CLR => 
        P_MASTER_POR_B_c_0, Q => P_USB_MASTER_EN_c_20);
    
    \T_CNT60M[3]\ : DFN1C0
      port map(D => T_CNT60M_n3, CLK => CLK60MHZ, CLR => 
        P_MASTER_POR_B_c_28, Q => \T_CNT60M[3]_net_1\);
    
    USB_EN_60M_2S : DFN1C0
      port map(D => \USB_EN_60M_1S\, CLK => CLK60MHZ, CLR => 
        P_MASTER_POR_B_c_22_0, Q => P_USB_MASTER_EN_c);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity EXEC_MODE_CNTL is

    port( CLK60MHZ                   : in    std_logic;
          P_USB_MASTER_EN_c_1_0      : out   std_logic;
          P_USB_MASTER_EN_c_2_0      : out   std_logic;
          P_USB_MASTER_EN_c_22_0     : out   std_logic;
          P_USB_MASTER_EN_c_22       : out   std_logic;
          P_USB_MASTER_EN_c_21       : out   std_logic;
          P_USB_MASTER_EN_c_20       : out   std_logic;
          P_USB_MASTER_EN_c_19       : out   std_logic;
          P_USB_MASTER_EN_c_18       : out   std_logic;
          P_USB_MASTER_EN_c_17       : out   std_logic;
          P_USB_MASTER_EN_c_16       : out   std_logic;
          P_USB_MASTER_EN_c_15       : out   std_logic;
          P_USB_MASTER_EN_c_14       : out   std_logic;
          P_USB_MASTER_EN_c_13       : out   std_logic;
          P_USB_MASTER_EN_c_12       : out   std_logic;
          P_USB_MASTER_EN_c_11       : out   std_logic;
          P_USB_MASTER_EN_c_10       : out   std_logic;
          P_USB_MASTER_EN_c_9        : out   std_logic;
          P_USB_MASTER_EN_c_8        : out   std_logic;
          P_USB_MASTER_EN_c_7        : out   std_logic;
          P_USB_MASTER_EN_c_6        : out   std_logic;
          P_USB_MASTER_EN_c_5        : out   std_logic;
          P_USB_MASTER_EN_c_4        : out   std_logic;
          P_USB_MASTER_EN_c_3        : out   std_logic;
          P_USB_MASTER_EN_c_2        : out   std_logic;
          P_USB_MASTER_EN_c_1        : out   std_logic;
          P_USB_MASTER_EN_c_0        : out   std_logic;
          P_USB_MASTER_EN_c          : out   std_logic;
          P_MASTER_POR_B_c           : out   std_logic;
          CCC_MAIN_LOCK              : in    std_logic;
          DCB_SALT_SEL_c             : in    std_logic;
          DEV_RST_B_c_1              : in    std_logic;
          MASTER_SALT_POR_B_i_0_i    : out   std_logic;
          MASTER_DCB_POR_B_i_0_i     : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_0  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_1  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_2  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_3  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_4  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_5  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_6  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_7  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_8  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_9  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_10 : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_11 : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_12 : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_13 : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_14 : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_15 : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_16 : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_17 : out   std_logic;
          P_MASTER_POR_B_c_1         : out   std_logic;
          P_MASTER_POR_B_c_2         : out   std_logic;
          P_MASTER_POR_B_c_3         : out   std_logic;
          P_MASTER_POR_B_c_4         : out   std_logic;
          P_MASTER_POR_B_c_5         : out   std_logic;
          P_MASTER_POR_B_c_6         : out   std_logic;
          P_MASTER_POR_B_c_7         : out   std_logic;
          P_MASTER_POR_B_c_8         : out   std_logic;
          P_MASTER_POR_B_c_9         : out   std_logic;
          P_MASTER_POR_B_c_10        : out   std_logic;
          P_MASTER_POR_B_c_11        : out   std_logic;
          P_MASTER_POR_B_c_12        : out   std_logic;
          P_MASTER_POR_B_c_13        : out   std_logic;
          P_MASTER_POR_B_c_14        : out   std_logic;
          P_MASTER_POR_B_c_15        : out   std_logic;
          P_MASTER_POR_B_c_16        : out   std_logic;
          P_MASTER_POR_B_c_17        : out   std_logic;
          P_MASTER_POR_B_c_18        : out   std_logic;
          P_MASTER_POR_B_c_19        : out   std_logic;
          P_MASTER_POR_B_c_20        : out   std_logic;
          P_MASTER_POR_B_c_21        : out   std_logic;
          P_MASTER_POR_B_c_22        : out   std_logic;
          P_MASTER_POR_B_c_23        : out   std_logic;
          P_MASTER_POR_B_c_24        : out   std_logic;
          P_MASTER_POR_B_c_25        : out   std_logic;
          P_MASTER_POR_B_c_26        : out   std_logic;
          P_MASTER_POR_B_c_27        : out   std_logic;
          P_MASTER_POR_B_c_28        : out   std_logic;
          P_MASTER_POR_B_c_29        : out   std_logic;
          P_MASTER_POR_B_c_30        : out   std_logic;
          P_MASTER_POR_B_c_31        : out   std_logic;
          P_MASTER_POR_B_c_32        : out   std_logic;
          P_MASTER_POR_B_c_33        : out   std_logic;
          P_MASTER_POR_B_c_34        : out   std_logic;
          P_MASTER_POR_B_c_34_0      : out   std_logic;
          P_MASTER_POR_B_c_32_0      : out   std_logic;
          P_MASTER_POR_B_c_31_0      : out   std_logic;
          P_MASTER_POR_B_c_27_0      : out   std_logic;
          P_MASTER_POR_B_c_27_1      : out   std_logic;
          P_MASTER_POR_B_c_24_0      : out   std_logic;
          P_MASTER_POR_B_c_22_0      : out   std_logic;
          P_MASTER_POR_B_c_17_0      : out   std_logic;
          P_MASTER_POR_B_c_16_0      : out   std_logic;
          DEV_RST_B_c                : in    std_logic;
          CCC_160M_FXD               : in    std_logic;
          CLK_40M_GL                 : in    std_logic;
          P_MASTER_POR_B_c_0_0       : out   std_logic
        );

end EXEC_MODE_CNTL;

architecture DEF_ARCH of EXEC_MODE_CNTL is 

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFI1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          QN  : out   std_logic
        );
  end component;

  component DFI1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          QN  : out   std_logic
        );
  end component;

  component XA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E0C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component OA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XNOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component USB_EXEC
    port( P_MASTER_POR_B_c_24    : in    std_logic := 'U';
          P_MASTER_POR_B_c_28    : in    std_logic := 'U';
          P_MASTER_POR_B_c_27    : in    std_logic := 'U';
          P_MASTER_POR_B_c_34_0  : in    std_logic := 'U';
          P_USB_MASTER_EN_c      : out   std_logic;
          P_MASTER_POR_B_c_29    : in    std_logic := 'U';
          P_MASTER_POR_B_c_32_0  : in    std_logic := 'U';
          CLK_40M_GL             : in    std_logic := 'U';
          P_MASTER_POR_B_c_23    : in    std_logic := 'U';
          P_USB_MASTER_EN_c_0    : out   std_logic;
          P_USB_MASTER_EN_c_1    : out   std_logic;
          P_USB_MASTER_EN_c_2    : out   std_logic;
          P_USB_MASTER_EN_c_3    : out   std_logic;
          P_USB_MASTER_EN_c_4    : out   std_logic;
          P_USB_MASTER_EN_c_5    : out   std_logic;
          P_USB_MASTER_EN_c_6    : out   std_logic;
          P_USB_MASTER_EN_c_7    : out   std_logic;
          P_USB_MASTER_EN_c_8    : out   std_logic;
          P_USB_MASTER_EN_c_9    : out   std_logic;
          P_USB_MASTER_EN_c_10   : out   std_logic;
          P_USB_MASTER_EN_c_11   : out   std_logic;
          P_USB_MASTER_EN_c_12   : out   std_logic;
          P_USB_MASTER_EN_c_13   : out   std_logic;
          P_USB_MASTER_EN_c_14   : out   std_logic;
          P_USB_MASTER_EN_c_15   : out   std_logic;
          P_USB_MASTER_EN_c_16   : out   std_logic;
          P_USB_MASTER_EN_c_17   : out   std_logic;
          P_USB_MASTER_EN_c_18   : out   std_logic;
          P_USB_MASTER_EN_c_19   : out   std_logic;
          P_USB_MASTER_EN_c_20   : out   std_logic;
          P_USB_MASTER_EN_c_21   : out   std_logic;
          P_MASTER_POR_B_c_0     : in    std_logic := 'U';
          P_USB_MASTER_EN_c_22   : out   std_logic;
          P_USB_MASTER_EN_c_22_0 : out   std_logic;
          P_USB_MASTER_EN_c_2_0  : out   std_logic;
          P_MASTER_POR_B_c_0_0   : in    std_logic := 'U';
          P_USB_MASTER_EN_c_1_0  : out   std_logic;
          P_MASTER_POR_B_c_22_0  : in    std_logic := 'U';
          CLK60MHZ               : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component OA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \P_MASTER_POR_B_c_0_0\, SYNC_BRD_RST_BI_i_0_i_2, 
        N_PRESCALE_2_sqmuxa, N_PRESCALE_2_sqmuxa_1, 
        un1_CCC_1_LOCK_STAT_1D_i_i_a2_0_5, 
        un1_CCC_1_LOCK_STAT_1D_i_i_a2_0_4, N_PRESCALE_2_sqmuxa_0, 
        DEV_RST_1B_i, SYNC_BRD_RST_BI_i_0_i_1, 
        SYNC_BRD_RST_BI_i_0_i_0, \P_MASTER_POR_B_c_22_0\, 
        \P_MASTER_POR_B_c_32_0\, \P_MASTER_POR_B_c_34_0\, 
        \P_MASTER_POR_B_c_29\, \P_MASTER_POR_B_c_28\, 
        \P_MASTER_POR_B_c_27\, \P_MASTER_POR_B_c_24\, 
        \P_MASTER_POR_B_c_23\, P_MASTER_POR_B_c_0, N_MPOR_SALT_B, 
        SYNC_BRD_RST_BI_i_0_i, \MPOR_DCB_B\, N_MPOR_DCB_B, 
        \DEV_RST_0B\, \DEL_CNT[4]_net_1\, \DEL_CNT[5]_net_1\, 
        un1_CCC_1_LOCK_STAT_1D_i_i_a2_0_3, \DEL_CNT[1]_net_1\, 
        \DEL_CNT[7]_net_1\, un1_CCC_1_LOCK_STAT_1D_i_i_a2_0_1, 
        \DEL_CNT[6]_net_1\, \CCC_1_LOCK_STAT_1D\, 
        \DEL_CNT[3]_net_1\, \DEL_CNT[2]_net_1\, PRESCALE_n2_i_0, 
        \PRESCALE[2]_net_1\, N_42, PRESCALE_n1_i_0, 
        \PRESCALE[0]_net_1\, \PRESCALE[1]_net_1\, 
        DEL_CNTlde_i_o2_0, \PRESCALE[3]_net_1\, N_17, N_47, N_92, 
        N_19, N_41, N_21, N_39, N_23, N_38, N_25, N_37, N_27, 
        \DEL_CNT[0]_net_1\, N_84, N_11, N_9, N_81_i, N_99, N_61, 
        N_15, N_31, N_63_i, N_7, N_82_i, \CCC_1_LOCK_STAT_0D\, 
        EXEC_MODE_CNTL_VCC, \GND\ : std_logic;

    for all : USB_EXEC
	Use entity work.USB_EXEC(DEF_ARCH);
begin 

    P_MASTER_POR_B_c_23 <= \P_MASTER_POR_B_c_23\;
    P_MASTER_POR_B_c_24 <= \P_MASTER_POR_B_c_24\;
    P_MASTER_POR_B_c_27 <= \P_MASTER_POR_B_c_27\;
    P_MASTER_POR_B_c_28 <= \P_MASTER_POR_B_c_28\;
    P_MASTER_POR_B_c_29 <= \P_MASTER_POR_B_c_29\;
    P_MASTER_POR_B_c_34_0 <= \P_MASTER_POR_B_c_34_0\;
    P_MASTER_POR_B_c_32_0 <= \P_MASTER_POR_B_c_32_0\;
    P_MASTER_POR_B_c_22_0 <= \P_MASTER_POR_B_c_22_0\;
    P_MASTER_POR_B_c_0_0 <= \P_MASTER_POR_B_c_0_0\;

    MPOR_B_22_0 : DFN1C0
      port map(D => N_PRESCALE_2_sqmuxa_0, CLK => CLK_40M_GL, CLR
         => SYNC_BRD_RST_BI_i_0_i_0, Q => \P_MASTER_POR_B_c_22_0\);
    
    MPOR_DCB_B_RNIPFG8 : CLKINT
      port map(A => \MPOR_DCB_B\, Y => MASTER_DCB_POR_B_i_0_i);
    
    SYNC_BRD_RST_BI_0 : DFI1P0
      port map(D => DEV_RST_1B_i, CLK => CCC_160M_FXD, PRE => 
        DEV_RST_B_c, QN => SYNC_BRD_RST_BI_i_0_i_0);
    
    MPOR_B_22 : DFN1C0
      port map(D => N_PRESCALE_2_sqmuxa_1, CLK => CLK_40M_GL, CLR
         => SYNC_BRD_RST_BI_i_0_i_1, Q => P_MASTER_POR_B_c_22);
    
    DEV_RST_1B : DFI1C0
      port map(D => \DEV_RST_0B\, CLK => CCC_160M_FXD, CLR => 
        DEV_RST_B_c_1, QN => DEV_RST_1B_i);
    
    MPOR_B_31_0 : DFN1C0
      port map(D => N_PRESCALE_2_sqmuxa_0, CLK => CLK_40M_GL, CLR
         => SYNC_BRD_RST_BI_i_0_i_0, Q => P_MASTER_POR_B_c_31_0);
    
    MPOR_SALT_B_9 : DFI1P0
      port map(D => N_MPOR_SALT_B, CLK => CLK_40M_GL, PRE => 
        SYNC_BRD_RST_BI_i_0_i_2, QN => MASTER_SALT_POR_B_i_0_i_9);
    
    \DEL_CNT_RNO[2]\ : XA1A
      port map(A => \DEL_CNT[2]_net_1\, B => N_37, C => 
        \CCC_1_LOCK_STAT_1D\, Y => N_25);
    
    MPOR_B_32_0 : DFN1C0
      port map(D => N_PRESCALE_2_sqmuxa_0, CLK => CLK_40M_GL, CLR
         => SYNC_BRD_RST_BI_i_0_i_0, Q => \P_MASTER_POR_B_c_32_0\);
    
    MPOR_B_10 : DFN1C0
      port map(D => N_PRESCALE_2_sqmuxa_1, CLK => CLK_40M_GL, CLR
         => SYNC_BRD_RST_BI_i_0_i_1, Q => P_MASTER_POR_B_c_10);
    
    MPOR_B_0_0 : DFN1C0
      port map(D => N_PRESCALE_2_sqmuxa, CLK => CLK_40M_GL, CLR
         => SYNC_BRD_RST_BI_i_0_i_2, Q => \P_MASTER_POR_B_c_0_0\);
    
    MPOR_B_32 : DFN1C0
      port map(D => N_PRESCALE_2_sqmuxa_0, CLK => CLK_40M_GL, CLR
         => SYNC_BRD_RST_BI_i_0_i_0, Q => P_MASTER_POR_B_c_32);
    
    MPOR_B_24 : DFN1C0
      port map(D => N_PRESCALE_2_sqmuxa_1, CLK => CLK_40M_GL, CLR
         => SYNC_BRD_RST_BI_i_0_i_0, Q => \P_MASTER_POR_B_c_24\);
    
    MPOR_B_23 : DFN1C0
      port map(D => N_PRESCALE_2_sqmuxa_1, CLK => CLK_40M_GL, CLR
         => SYNC_BRD_RST_BI_i_0_i_1, Q => \P_MASTER_POR_B_c_23\);
    
    CCC_1_LOCK_STAT_0D : DFN1C0
      port map(D => CCC_MAIN_LOCK, CLK => CLK_40M_GL, CLR => 
        SYNC_BRD_RST_BI_i_0_i, Q => \CCC_1_LOCK_STAT_0D\);
    
    MPOR_B_27_1 : DFN1C0
      port map(D => N_PRESCALE_2_sqmuxa_0, CLK => CLK_40M_GL, CLR
         => SYNC_BRD_RST_BI_i_0_i_0, Q => P_MASTER_POR_B_c_27_1);
    
    \DEL_CNT[1]\ : DFN1E0C0
      port map(D => N_27, CLK => CLK_40M_GL, CLR => 
        SYNC_BRD_RST_BI_i_0_i, E => N_31, Q => \DEL_CNT[1]_net_1\);
    
    MPOR_SALT_B_6 : DFI1P0
      port map(D => N_MPOR_SALT_B, CLK => CLK_40M_GL, PRE => 
        SYNC_BRD_RST_BI_i_0_i_2, QN => MASTER_SALT_POR_B_i_0_i_6);
    
    MPOR_SALT_B_13 : DFI1P0
      port map(D => N_MPOR_SALT_B, CLK => CLK_40M_GL, PRE => 
        SYNC_BRD_RST_BI_i_0_i_2, QN => MASTER_SALT_POR_B_i_0_i_13);
    
    \DEL_CNT_RNIMTCH1[4]\ : OR2A
      port map(A => N_PRESCALE_2_sqmuxa, B => DCB_SALT_SEL_c, Y
         => N_MPOR_SALT_B);
    
    \PRESCALE_RNO[0]\ : NOR3B
      port map(A => \CCC_1_LOCK_STAT_1D\, B => N_84, C => 
        \PRESCALE[0]_net_1\, Y => N_82_i);
    
    \PRESCALE_RNO_0[3]\ : AX1A
      port map(A => N_42, B => \PRESCALE[2]_net_1\, C => 
        \PRESCALE[3]_net_1\, Y => N_63_i);
    
    MPOR_B_34 : DFN1C0
      port map(D => N_PRESCALE_2_sqmuxa_0, CLK => CLK_40M_GL, CLR
         => SYNC_BRD_RST_BI_i_0_i_0, Q => P_MASTER_POR_B_c_34);
    
    MPOR_B_33 : DFN1C0
      port map(D => N_PRESCALE_2_sqmuxa_0, CLK => CLK_40M_GL, CLR
         => SYNC_BRD_RST_BI_i_0_i_0, Q => P_MASTER_POR_B_c_33);
    
    \DEL_CNT[3]\ : DFN1E0C0
      port map(D => N_23, CLK => CLK_40M_GL, CLR => 
        SYNC_BRD_RST_BI_i_0_i, E => N_31, Q => \DEL_CNT[3]_net_1\);
    
    SYNC_BRD_RST_BI : DFI1P0
      port map(D => DEV_RST_1B_i, CLK => CCC_160M_FXD, PRE => 
        DEV_RST_B_c, QN => SYNC_BRD_RST_BI_i_0_i);
    
    MPOR_SALT_B_2 : DFI1P0
      port map(D => N_MPOR_SALT_B, CLK => CLK_40M_GL, PRE => 
        SYNC_BRD_RST_BI_i_0_i_2, QN => MASTER_SALT_POR_B_i_0_i_2);
    
    MPOR_B_20 : DFN1C0
      port map(D => N_PRESCALE_2_sqmuxa_1, CLK => CLK_40M_GL, CLR
         => SYNC_BRD_RST_BI_i_0_i_1, Q => P_MASTER_POR_B_c_20);
    
    MPOR_SALT_B_12 : DFI1P0
      port map(D => N_MPOR_SALT_B, CLK => CLK_40M_GL, PRE => 
        SYNC_BRD_RST_BI_i_0_i_2, QN => MASTER_SALT_POR_B_i_0_i_12);
    
    VCC_i : VCC
      port map(Y => EXEC_MODE_CNTL_VCC);
    
    MPOR_SALT_B_14 : DFI1P0
      port map(D => N_MPOR_SALT_B, CLK => CLK_40M_GL, PRE => 
        SYNC_BRD_RST_BI_i_0_i_2, QN => MASTER_SALT_POR_B_i_0_i_14);
    
    CCC_1_LOCK_STAT_1D_RNICAH41 : OA1
      port map(A => N_61, B => DEL_CNTlde_i_o2_0, C => 
        \CCC_1_LOCK_STAT_1D\, Y => N_99);
    
    MPOR_DCB_B_RNO : OR2B
      port map(A => N_PRESCALE_2_sqmuxa, B => DCB_SALT_SEL_c, Y
         => N_MPOR_DCB_B);
    
    MPOR_B_15 : DFN1C0
      port map(D => N_PRESCALE_2_sqmuxa_1, CLK => CLK_40M_GL, CLR
         => SYNC_BRD_RST_BI_i_0_i_1, Q => P_MASTER_POR_B_c_15);
    
    \DEL_CNT_RNIPJUG[7]\ : NOR3C
      port map(A => \DEL_CNT[1]_net_1\, B => \DEL_CNT[7]_net_1\, 
        C => un1_CCC_1_LOCK_STAT_1D_i_i_a2_0_1, Y => 
        un1_CCC_1_LOCK_STAT_1D_i_i_a2_0_4);
    
    \PRESCALE[3]\ : DFN1E0C0
      port map(D => N_7, CLK => CLK_40M_GL, CLR => 
        SYNC_BRD_RST_BI_i_0_i, E => N_PRESCALE_2_sqmuxa, Q => 
        \PRESCALE[3]_net_1\);
    
    MPOR_B_11 : DFN1C0
      port map(D => N_PRESCALE_2_sqmuxa_1, CLK => CLK_40M_GL, CLR
         => SYNC_BRD_RST_BI_i_0_i_1, Q => P_MASTER_POR_B_c_11);
    
    MPOR_B_16 : DFN1C0
      port map(D => N_PRESCALE_2_sqmuxa_1, CLK => CLK_40M_GL, CLR
         => SYNC_BRD_RST_BI_i_0_i_1, Q => P_MASTER_POR_B_c_16);
    
    \PRESCALE_RNO[1]\ : NOR3B
      port map(A => \CCC_1_LOCK_STAT_1D\, B => N_84, C => 
        PRESCALE_n1_i_0, Y => N_11);
    
    MPOR_B_30 : DFN1C0
      port map(D => N_PRESCALE_2_sqmuxa_0, CLK => CLK_40M_GL, CLR
         => SYNC_BRD_RST_BI_i_0_i_0, Q => P_MASTER_POR_B_c_30);
    
    \DEL_CNT_RNO_0[6]\ : OA1C
      port map(A => \DEL_CNT[5]_net_1\, B => N_41, C => 
        \DEL_CNT[6]_net_1\, Y => N_92);
    
    MPOR_SALT_B_5 : DFI1P0
      port map(D => N_MPOR_SALT_B, CLK => CLK_40M_GL, PRE => 
        SYNC_BRD_RST_BI_i_0_i_2, QN => MASTER_SALT_POR_B_i_0_i_5);
    
    MPOR_SALT_B_16 : DFI1P0
      port map(D => N_MPOR_SALT_B, CLK => CLK_40M_GL, PRE => 
        SYNC_BRD_RST_BI_i_0_i_2, QN => MASTER_SALT_POR_B_i_0_i_16);
    
    \DEL_CNT_RNI74F8[0]\ : OR2B
      port map(A => \DEL_CNT[1]_net_1\, B => \DEL_CNT[0]_net_1\, 
        Y => N_37);
    
    \PRESCALE_RNO[2]\ : NOR3B
      port map(A => \CCC_1_LOCK_STAT_1D\, B => N_84, C => 
        PRESCALE_n2_i_0, Y => N_9);
    
    \DEL_CNT_RNIAJAL[4]\ : NOR3C
      port map(A => \DEL_CNT[4]_net_1\, B => \DEL_CNT[5]_net_1\, 
        C => un1_CCC_1_LOCK_STAT_1D_i_i_a2_0_3, Y => 
        un1_CCC_1_LOCK_STAT_1D_i_i_a2_0_5);
    
    \DEL_CNT_RNI37961_1[4]\ : NOR2B
      port map(A => un1_CCC_1_LOCK_STAT_1D_i_i_a2_0_5, B => 
        un1_CCC_1_LOCK_STAT_1D_i_i_a2_0_4, Y => 
        N_PRESCALE_2_sqmuxa);
    
    \PRESCALE_RNO_0[1]\ : XNOR2
      port map(A => \PRESCALE[0]_net_1\, B => \PRESCALE[1]_net_1\, 
        Y => PRESCALE_n1_i_0);
    
    \DEL_CNT_RNI37961_0[4]\ : NOR2B
      port map(A => un1_CCC_1_LOCK_STAT_1D_i_i_a2_0_5, B => 
        un1_CCC_1_LOCK_STAT_1D_i_i_a2_0_4, Y => 
        N_PRESCALE_2_sqmuxa_1);
    
    MPOR_B_25 : DFN1C0
      port map(D => N_PRESCALE_2_sqmuxa_1, CLK => CLK_40M_GL, CLR
         => SYNC_BRD_RST_BI_i_0_i_0, Q => P_MASTER_POR_B_c_25);
    
    \PRESCALE[2]\ : DFN1E0C0
      port map(D => N_9, CLK => CLK_40M_GL, CLR => 
        SYNC_BRD_RST_BI_i_0_i, E => N_PRESCALE_2_sqmuxa, Q => 
        \PRESCALE[2]_net_1\);
    
    MPOR_SALT_B_15 : DFI1P0
      port map(D => N_MPOR_SALT_B, CLK => CLK_40M_GL, PRE => 
        SYNC_BRD_RST_BI_i_0_i_2, QN => MASTER_SALT_POR_B_i_0_i_15);
    
    MPOR_B_21 : DFN1C0
      port map(D => N_PRESCALE_2_sqmuxa_1, CLK => CLK_40M_GL, CLR
         => SYNC_BRD_RST_BI_i_0_i_1, Q => P_MASTER_POR_B_c_21);
    
    MPOR_SALT_B_8 : DFI1P0
      port map(D => N_MPOR_SALT_B, CLK => CLK_40M_GL, PRE => 
        SYNC_BRD_RST_BI_i_0_i_2, QN => MASTER_SALT_POR_B_i_0_i_8);
    
    MPOR_B_26 : DFN1C0
      port map(D => N_PRESCALE_2_sqmuxa_0, CLK => CLK_40M_GL, CLR
         => SYNC_BRD_RST_BI_i_0_i_0, Q => P_MASTER_POR_B_c_26);
    
    \DEL_CNT_RNO[1]\ : XA1
      port map(A => \DEL_CNT[0]_net_1\, B => \DEL_CNT[1]_net_1\, 
        C => \CCC_1_LOCK_STAT_1D\, Y => N_27);
    
    \PRESCALE_RNIJRUD_0[0]\ : OR2
      port map(A => \PRESCALE[1]_net_1\, B => \PRESCALE[0]_net_1\, 
        Y => N_61);
    
    \DEL_CNT_RNO[0]\ : NOR2A
      port map(A => \CCC_1_LOCK_STAT_1D\, B => \DEL_CNT[0]_net_1\, 
        Y => N_81_i);
    
    \DEL_CNT_RNI926L[4]\ : OR2A
      port map(A => \DEL_CNT[4]_net_1\, B => N_39, Y => N_41);
    
    MPOR_B_9 : DFN1C0
      port map(D => N_PRESCALE_2_sqmuxa_1, CLK => CLK_40M_GL, CLR
         => SYNC_BRD_RST_BI_i_0_i_1, Q => P_MASTER_POR_B_c_9);
    
    MPOR_B_31 : DFN1C0
      port map(D => N_PRESCALE_2_sqmuxa_0, CLK => CLK_40M_GL, CLR
         => SYNC_BRD_RST_BI_i_0_i_0, Q => P_MASTER_POR_B_c_31);
    
    MPOR_B_17 : DFN1C0
      port map(D => N_PRESCALE_2_sqmuxa_1, CLK => CLK_40M_GL, CLR
         => SYNC_BRD_RST_BI_i_0_i_1, Q => P_MASTER_POR_B_c_17);
    
    \PRESCALE_RNO_0[2]\ : XOR2
      port map(A => \PRESCALE[2]_net_1\, B => N_42, Y => 
        PRESCALE_n2_i_0);
    
    \DEL_CNT_RNI37961[4]\ : NOR2B
      port map(A => un1_CCC_1_LOCK_STAT_1D_i_i_a2_0_5, B => 
        un1_CCC_1_LOCK_STAT_1D_i_i_a2_0_4, Y => 
        N_PRESCALE_2_sqmuxa_0);
    
    \DEL_CNT[0]\ : DFN1E0C0
      port map(D => N_81_i, CLK => CLK_40M_GL, CLR => 
        SYNC_BRD_RST_BI_i_0_i, E => N_31, Q => \DEL_CNT[0]_net_1\);
    
    MPOR_B_6 : DFN1C0
      port map(D => N_PRESCALE_2_sqmuxa, CLK => CLK_40M_GL, CLR
         => SYNC_BRD_RST_BI_i_0_i_1, Q => P_MASTER_POR_B_c_6);
    
    MPOR_B_1 : DFN1C0
      port map(D => N_PRESCALE_2_sqmuxa, CLK => CLK_40M_GL, CLR
         => SYNC_BRD_RST_BI_i_0_i_2, Q => P_MASTER_POR_B_c_1);
    
    MPOR_B_5 : DFN1C0
      port map(D => N_PRESCALE_2_sqmuxa, CLK => CLK_40M_GL, CLR
         => SYNC_BRD_RST_BI_i_0_i_1, Q => P_MASTER_POR_B_c_5);
    
    MPOR_B_27_0 : DFN1C0
      port map(D => N_PRESCALE_2_sqmuxa_0, CLK => CLK_40M_GL, CLR
         => SYNC_BRD_RST_BI_i_0_i_0, Q => P_MASTER_POR_B_c_27_0);
    
    \DEL_CNT_RNISNMC[2]\ : OR2A
      port map(A => \DEL_CNT[2]_net_1\, B => N_37, Y => N_38);
    
    \PRESCALE[0]\ : DFN1E0C0
      port map(D => N_82_i, CLK => CLK_40M_GL, CLR => 
        SYNC_BRD_RST_BI_i_0_i, E => N_PRESCALE_2_sqmuxa, Q => 
        \PRESCALE[0]_net_1\);
    
    MPOR_B_4 : DFN1C0
      port map(D => N_PRESCALE_2_sqmuxa, CLK => CLK_40M_GL, CLR
         => SYNC_BRD_RST_BI_i_0_i_1, Q => P_MASTER_POR_B_c_4);
    
    \DEL_CNT[2]\ : DFN1E0C0
      port map(D => N_25, CLK => CLK_40M_GL, CLR => 
        SYNC_BRD_RST_BI_i_0_i, E => N_31, Q => \DEL_CNT[2]_net_1\);
    
    MPOR_B_8 : DFN1C0
      port map(D => N_PRESCALE_2_sqmuxa_1, CLK => CLK_40M_GL, CLR
         => SYNC_BRD_RST_BI_i_0_i_1, Q => P_MASTER_POR_B_c_8);
    
    MPOR_B_27 : DFN1C0
      port map(D => N_PRESCALE_2_sqmuxa_0, CLK => CLK_40M_GL, CLR
         => SYNC_BRD_RST_BI_i_0_i_0, Q => \P_MASTER_POR_B_c_27\);
    
    MPOR_B_0 : DFN1C0
      port map(D => N_PRESCALE_2_sqmuxa, CLK => CLK_40M_GL, CLR
         => SYNC_BRD_RST_BI_i_0_i_2, Q => P_MASTER_POR_B_c_0);
    
    USB_MASTER_EN : USB_EXEC
      port map(P_MASTER_POR_B_c_24 => \P_MASTER_POR_B_c_24\, 
        P_MASTER_POR_B_c_28 => \P_MASTER_POR_B_c_28\, 
        P_MASTER_POR_B_c_27 => \P_MASTER_POR_B_c_27\, 
        P_MASTER_POR_B_c_34_0 => \P_MASTER_POR_B_c_34_0\, 
        P_USB_MASTER_EN_c => P_USB_MASTER_EN_c, 
        P_MASTER_POR_B_c_29 => \P_MASTER_POR_B_c_29\, 
        P_MASTER_POR_B_c_32_0 => \P_MASTER_POR_B_c_32_0\, 
        CLK_40M_GL => CLK_40M_GL, P_MASTER_POR_B_c_23 => 
        \P_MASTER_POR_B_c_23\, P_USB_MASTER_EN_c_0 => 
        P_USB_MASTER_EN_c_0, P_USB_MASTER_EN_c_1 => 
        P_USB_MASTER_EN_c_1, P_USB_MASTER_EN_c_2 => 
        P_USB_MASTER_EN_c_2, P_USB_MASTER_EN_c_3 => 
        P_USB_MASTER_EN_c_3, P_USB_MASTER_EN_c_4 => 
        P_USB_MASTER_EN_c_4, P_USB_MASTER_EN_c_5 => 
        P_USB_MASTER_EN_c_5, P_USB_MASTER_EN_c_6 => 
        P_USB_MASTER_EN_c_6, P_USB_MASTER_EN_c_7 => 
        P_USB_MASTER_EN_c_7, P_USB_MASTER_EN_c_8 => 
        P_USB_MASTER_EN_c_8, P_USB_MASTER_EN_c_9 => 
        P_USB_MASTER_EN_c_9, P_USB_MASTER_EN_c_10 => 
        P_USB_MASTER_EN_c_10, P_USB_MASTER_EN_c_11 => 
        P_USB_MASTER_EN_c_11, P_USB_MASTER_EN_c_12 => 
        P_USB_MASTER_EN_c_12, P_USB_MASTER_EN_c_13 => 
        P_USB_MASTER_EN_c_13, P_USB_MASTER_EN_c_14 => 
        P_USB_MASTER_EN_c_14, P_USB_MASTER_EN_c_15 => 
        P_USB_MASTER_EN_c_15, P_USB_MASTER_EN_c_16 => 
        P_USB_MASTER_EN_c_16, P_USB_MASTER_EN_c_17 => 
        P_USB_MASTER_EN_c_17, P_USB_MASTER_EN_c_18 => 
        P_USB_MASTER_EN_c_18, P_USB_MASTER_EN_c_19 => 
        P_USB_MASTER_EN_c_19, P_USB_MASTER_EN_c_20 => 
        P_USB_MASTER_EN_c_20, P_USB_MASTER_EN_c_21 => 
        P_USB_MASTER_EN_c_21, P_MASTER_POR_B_c_0 => 
        P_MASTER_POR_B_c_0, P_USB_MASTER_EN_c_22 => 
        P_USB_MASTER_EN_c_22, P_USB_MASTER_EN_c_22_0 => 
        P_USB_MASTER_EN_c_22_0, P_USB_MASTER_EN_c_2_0 => 
        P_USB_MASTER_EN_c_2_0, P_MASTER_POR_B_c_0_0 => 
        \P_MASTER_POR_B_c_0_0\, P_USB_MASTER_EN_c_1_0 => 
        P_USB_MASTER_EN_c_1_0, P_MASTER_POR_B_c_22_0 => 
        \P_MASTER_POR_B_c_22_0\, CLK60MHZ => CLK60MHZ);
    
    \PRESCALE_RNINVUD[3]\ : OR2
      port map(A => \PRESCALE[3]_net_1\, B => \PRESCALE[2]_net_1\, 
        Y => DEL_CNTlde_i_o2_0);
    
    MPOR_SALT_B_0 : DFI1P0
      port map(D => N_MPOR_SALT_B, CLK => CLK_40M_GL, PRE => 
        SYNC_BRD_RST_BI_i_0_i, QN => MASTER_SALT_POR_B_i_0_i_0);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \DEL_CNT_RNIICUG[3]\ : OR2A
      port map(A => \DEL_CNT[3]_net_1\, B => N_38, Y => N_39);
    
    CCC_1_LOCK_STAT_1D : DFN1C0
      port map(D => \CCC_1_LOCK_STAT_0D\, CLK => CLK_40M_GL, CLR
         => SYNC_BRD_RST_BI_i_0_i, Q => \CCC_1_LOCK_STAT_1D\);
    
    MPOR_SALT_B_3 : DFI1P0
      port map(D => N_MPOR_SALT_B, CLK => CLK_40M_GL, PRE => 
        SYNC_BRD_RST_BI_i_0_i_2, QN => MASTER_SALT_POR_B_i_0_i_3);
    
    MPOR_B_7 : DFN1C0
      port map(D => N_PRESCALE_2_sqmuxa, CLK => CLK_40M_GL, CLR
         => SYNC_BRD_RST_BI_i_0_i_1, Q => P_MASTER_POR_B_c_7);
    
    \DEL_CNT[6]\ : DFN1E0C0
      port map(D => N_17, CLK => CLK_40M_GL, CLR => 
        SYNC_BRD_RST_BI_i_0_i, E => N_31, Q => \DEL_CNT[6]_net_1\);
    
    SYNC_BRD_RST_BI_2 : DFI1P0
      port map(D => DEV_RST_1B_i, CLK => CCC_160M_FXD, PRE => 
        DEV_RST_B_c, QN => SYNC_BRD_RST_BI_i_0_i_2);
    
    MPOR_SALT_B_4 : DFI1P0
      port map(D => N_MPOR_SALT_B, CLK => CLK_40M_GL, PRE => 
        SYNC_BRD_RST_BI_i_0_i_2, QN => MASTER_SALT_POR_B_i_0_i_4);
    
    MPOR_B_2 : DFN1C0
      port map(D => N_PRESCALE_2_sqmuxa, CLK => CLK_40M_GL, CLR
         => SYNC_BRD_RST_BI_i_0_i_2, Q => P_MASTER_POR_B_c_2);
    
    \DEL_CNT[4]\ : DFN1E0C0
      port map(D => N_21, CLK => CLK_40M_GL, CLR => 
        SYNC_BRD_RST_BI_i_0_i, E => N_31, Q => \DEL_CNT[4]_net_1\);
    
    \PRESCALE_RNO[3]\ : NOR3B
      port map(A => \CCC_1_LOCK_STAT_1D\, B => N_84, C => N_63_i, 
        Y => N_7);
    
    MPOR_B_24_0 : DFN1C0
      port map(D => N_PRESCALE_2_sqmuxa_0, CLK => CLK_40M_GL, CLR
         => SYNC_BRD_RST_BI_i_0_i_0, Q => P_MASTER_POR_B_c_24_0);
    
    MPOR_B_3 : DFN1C0
      port map(D => N_PRESCALE_2_sqmuxa, CLK => CLK_40M_GL, CLR
         => SYNC_BRD_RST_BI_i_0_i_2, Q => P_MASTER_POR_B_c_3);
    
    \DEL_CNT_RNO[7]\ : OA1A
      port map(A => N_47, B => \DEL_CNT[7]_net_1\, C => 
        \CCC_1_LOCK_STAT_1D\, Y => N_15);
    
    MPOR_SALT_B_17 : DFI1P0
      port map(D => N_MPOR_SALT_B, CLK => CLK_40M_GL, PRE => 
        SYNC_BRD_RST_BI_i_0_i_2, QN => MASTER_SALT_POR_B_i_0_i_17);
    
    \DEL_CNT_RNIB8F8[2]\ : NOR2B
      port map(A => \DEL_CNT[3]_net_1\, B => \DEL_CNT[2]_net_1\, 
        Y => un1_CCC_1_LOCK_STAT_1D_i_i_a2_0_1);
    
    MPOR_B_34_0 : DFN1C0
      port map(D => N_PRESCALE_2_sqmuxa_0, CLK => CLK_40M_GL, CLR
         => SYNC_BRD_RST_BI_i_0_i_0, Q => \P_MASTER_POR_B_c_34_0\);
    
    SYNC_BRD_RST_BI_1 : DFI1P0
      port map(D => DEV_RST_1B_i, CLK => CCC_160M_FXD, PRE => 
        DEV_RST_B_c, QN => SYNC_BRD_RST_BI_i_0_i_1);
    
    \PRESCALE[1]\ : DFN1E0C0
      port map(D => N_11, CLK => CLK_40M_GL, CLR => 
        SYNC_BRD_RST_BI_i_0_i, E => N_PRESCALE_2_sqmuxa, Q => 
        \PRESCALE[1]_net_1\);
    
    MPOR_B_17_0 : DFN1C0
      port map(D => N_PRESCALE_2_sqmuxa_0, CLK => CLK_40M_GL, CLR
         => SYNC_BRD_RST_BI_i_0_i_0, Q => P_MASTER_POR_B_c_17_0);
    
    MPOR_B_16_0 : DFN1C0
      port map(D => N_PRESCALE_2_sqmuxa_0, CLK => CLK_40M_GL, CLR
         => SYNC_BRD_RST_BI_i_0_i_0, Q => P_MASTER_POR_B_c_16_0);
    
    CCC_1_LOCK_STAT_1D_RNIFHQA2 : OR2
      port map(A => N_99, B => N_PRESCALE_2_sqmuxa, Y => N_31);
    
    MPOR_B_19 : DFN1C0
      port map(D => N_PRESCALE_2_sqmuxa_1, CLK => CLK_40M_GL, CLR
         => SYNC_BRD_RST_BI_i_0_i_1, Q => P_MASTER_POR_B_c_19);
    
    \DEL_CNT_RNIR6RC[6]\ : NOR2B
      port map(A => \DEL_CNT[6]_net_1\, B => \CCC_1_LOCK_STAT_1D\, 
        Y => un1_CCC_1_LOCK_STAT_1D_i_i_a2_0_3);
    
    MPOR_B_18 : DFN1C0
      port map(D => N_PRESCALE_2_sqmuxa_1, CLK => CLK_40M_GL, CLR
         => SYNC_BRD_RST_BI_i_0_i_1, Q => P_MASTER_POR_B_c_18);
    
    DEV_RST_0B : DFN1C0
      port map(D => EXEC_MODE_CNTL_VCC, CLK => CCC_160M_FXD, CLR
         => DEV_RST_B_c_1, Q => \DEV_RST_0B\);
    
    MPOR_SALT_B_11 : DFI1P0
      port map(D => N_MPOR_SALT_B, CLK => CLK_40M_GL, PRE => 
        SYNC_BRD_RST_BI_i_0_i_2, QN => MASTER_SALT_POR_B_i_0_i_11);
    
    \DEL_CNT_RNIQGLT[6]\ : OR3B
      port map(A => \DEL_CNT[5]_net_1\, B => \DEL_CNT[6]_net_1\, 
        C => N_41, Y => N_47);
    
    \PRESCALE_RNIJRUD[0]\ : OR2B
      port map(A => \PRESCALE[1]_net_1\, B => \PRESCALE[0]_net_1\, 
        Y => N_42);
    
    MPOR_B_29 : DFN1C0
      port map(D => N_PRESCALE_2_sqmuxa_0, CLK => CLK_40M_GL, CLR
         => SYNC_BRD_RST_BI_i_0_i_0, Q => \P_MASTER_POR_B_c_29\);
    
    MPOR_SALT_B_7 : DFI1P0
      port map(D => N_MPOR_SALT_B, CLK => CLK_40M_GL, PRE => 
        SYNC_BRD_RST_BI_i_0_i_2, QN => MASTER_SALT_POR_B_i_0_i_7);
    
    MPOR_SALT_B_10 : DFI1P0
      port map(D => N_MPOR_SALT_B, CLK => CLK_40M_GL, PRE => 
        SYNC_BRD_RST_BI_i_0_i_2, QN => MASTER_SALT_POR_B_i_0_i_10);
    
    \PRESCALE_RNI1EUK[3]\ : OR3C
      port map(A => \PRESCALE[1]_net_1\, B => \PRESCALE[3]_net_1\, 
        C => \PRESCALE[2]_net_1\, Y => N_84);
    
    MPOR_SALT_B : DFI1P0
      port map(D => N_MPOR_SALT_B, CLK => CLK_40M_GL, PRE => 
        SYNC_BRD_RST_BI_i_0_i, QN => MASTER_SALT_POR_B_i_0_i);
    
    MPOR_B_28 : DFN1C0
      port map(D => N_PRESCALE_2_sqmuxa_0, CLK => CLK_40M_GL, CLR
         => SYNC_BRD_RST_BI_i_0_i_0, Q => \P_MASTER_POR_B_c_28\);
    
    MPOR_DCB_B : DFI1P0
      port map(D => N_MPOR_DCB_B, CLK => CLK_40M_GL, PRE => 
        SYNC_BRD_RST_BI_i_0_i, QN => \MPOR_DCB_B\);
    
    MPOR_B_12 : DFN1C0
      port map(D => N_PRESCALE_2_sqmuxa_1, CLK => CLK_40M_GL, CLR
         => SYNC_BRD_RST_BI_i_0_i_1, Q => P_MASTER_POR_B_c_12);
    
    \DEL_CNT_RNO[3]\ : XA1A
      port map(A => \DEL_CNT[3]_net_1\, B => N_38, C => 
        \CCC_1_LOCK_STAT_1D\, Y => N_23);
    
    \DEL_CNT[7]\ : DFN1E0C0
      port map(D => N_15, CLK => CLK_40M_GL, CLR => 
        SYNC_BRD_RST_BI_i_0_i, E => N_31, Q => \DEL_CNT[7]_net_1\);
    
    MPOR_SALT_B_1 : DFI1P0
      port map(D => N_MPOR_SALT_B, CLK => CLK_40M_GL, PRE => 
        SYNC_BRD_RST_BI_i_0_i, QN => MASTER_SALT_POR_B_i_0_i_1);
    
    \DEL_CNT_RNO[5]\ : XA1A
      port map(A => \DEL_CNT[5]_net_1\, B => N_41, C => 
        \CCC_1_LOCK_STAT_1D\, Y => N_19);
    
    \DEL_CNT_RNO[6]\ : NOR3B
      port map(A => \CCC_1_LOCK_STAT_1D\, B => N_47, C => N_92, Y
         => N_17);
    
    \DEL_CNT[5]\ : DFN1E0C0
      port map(D => N_19, CLK => CLK_40M_GL, CLR => 
        SYNC_BRD_RST_BI_i_0_i, E => N_31, Q => \DEL_CNT[5]_net_1\);
    
    \DEL_CNT_RNO[4]\ : XA1A
      port map(A => \DEL_CNT[4]_net_1\, B => N_39, C => 
        \CCC_1_LOCK_STAT_1D\, Y => N_21);
    
    MPOR_B_14 : DFN1C0
      port map(D => N_PRESCALE_2_sqmuxa_1, CLK => CLK_40M_GL, CLR
         => SYNC_BRD_RST_BI_i_0_i_1, Q => P_MASTER_POR_B_c_14);
    
    MPOR_B_13 : DFN1C0
      port map(D => N_PRESCALE_2_sqmuxa_1, CLK => CLK_40M_GL, CLR
         => SYNC_BRD_RST_BI_i_0_i_1, Q => P_MASTER_POR_B_c_13);
    
    MPOR_B : DFN1C0
      port map(D => N_PRESCALE_2_sqmuxa, CLK => CLK_40M_GL, CLR
         => SYNC_BRD_RST_BI_i_0_i, Q => P_MASTER_POR_B_c);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SLAVE_DES320S_1_17_5 is

    port( ELK_RX_SER_WORD_7      : out   std_logic_vector(7 downto 0);
          BIT_OS_SEL_0           : in    std_logic;
          BIT_OS_SEL_5_2         : in    std_logic;
          BIT_OS_SEL_5_0         : in    std_logic;
          BIT_OS_SEL_6           : in    std_logic_vector(2 downto 1);
          BIT_OS_SEL_4           : in    std_logic_vector(2 downto 1);
          CLK_40M_GL             : in    std_logic;
          CCC_160M_FXD           : in    std_logic;
          ELK_IN_R               : in    std_logic;
          ELK_IN_F               : in    std_logic;
          MASTER_DCB_POR_B_i_0_i : in    std_logic;
          CCC_160M_ADJ           : in    std_logic
        );

end SLAVE_DES320S_1_17_5;

architecture DEF_ARCH of SLAVE_DES320S_1_17_5 is 

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal N_17, \ARB_BYTE[0]_net_1\, \ARB_BYTE[4]_net_1\, N_18, 
        \ARB_BYTE[1]_net_1\, \ARB_BYTE[5]_net_1\, N_19, 
        \ARB_BYTE[2]_net_1\, \ARB_BYTE[6]_net_1\, N_20, 
        \ARB_BYTE[3]_net_1\, \ARB_BYTE[7]_net_1\, N_21, 
        \ARB_BYTE[8]_net_1\, N_22, \ARB_BYTE[9]_net_1\, N_23, 
        \ARB_BYTE[10]_net_1\, N_24, \ARB_BYTE[11]_net_1\, N_31, 
        \ARB_BYTE[12]_net_1\, N_32, \ARB_BYTE[13]_net_1\, N_33, 
        N_34, N_35, N_36, N_37, N_38, N_39, N_40, N_56, 
        \ARB_BYTE[14]_net_1\, N_64, \N_RECD_SER_WORD[0]\, 
        \N_RECD_SER_WORD[1]\, \N_RECD_SER_WORD[2]\, 
        \N_RECD_SER_WORD[3]\, \N_RECD_SER_WORD[4]\, 
        \N_RECD_SER_WORD[5]\, \N_RECD_SER_WORD[6]\, 
        \N_RECD_SER_WORD[7]\, \ADJ_SER_IN_F_0DEL\, 
        \ADJ_SER_IN_R_0DEL\, \ADJ_SER_IN_F_1DEL\, 
        \ADJ_SER_IN_R_1DEL\, \Q[0]_net_1\, \ADJ_Q[0]_net_1\, 
        \Q[1]_net_1\, \ADJ_Q[1]_net_1\, \Q[2]_net_1\, 
        \ADJ_Q[2]_net_1\, \Q[3]_net_1\, \ADJ_Q[3]_net_1\, 
        \Q[4]_net_1\, \ADJ_Q[4]_net_1\, \Q[5]_net_1\, 
        \ADJ_Q[5]_net_1\, \Q[6]_net_1\, \ADJ_Q[6]_net_1\, 
        \Q[7]_net_1\, \ADJ_Q[7]_net_1\, \Q[8]_net_1\, 
        \ADJ_Q[8]_net_1\, \Q[9]_net_1\, \ADJ_Q[9]_net_1\, 
        \Q[10]_net_1\, \ADJ_Q[10]_net_1\, \Q[11]_net_1\, 
        \ADJ_Q[11]_net_1\, \Q[12]_net_1\, \ADJ_Q[12]_net_1\, 
        \Q[13]_net_1\, \ADJ_Q[13]_net_1\, \Q[14]_net_1\, 
        \ADJ_Q[14]_net_1\, \ARB_WRD_40M_FIXED[0]_net_1\, 
        \ARB_WRD_40M_FIXED[1]_net_1\, 
        \ARB_WRD_40M_FIXED[2]_net_1\, 
        \ARB_WRD_40M_FIXED[3]_net_1\, 
        \ARB_WRD_40M_FIXED[4]_net_1\, 
        \ARB_WRD_40M_FIXED[5]_net_1\, 
        \ARB_WRD_40M_FIXED[6]_net_1\, 
        \ARB_WRD_40M_FIXED[7]_net_1\, 
        \ARB_WRD_40M_FIXED[8]_net_1\, 
        \ARB_WRD_40M_FIXED[9]_net_1\, 
        \ARB_WRD_40M_FIXED[10]_net_1\, 
        \ARB_WRD_40M_FIXED[11]_net_1\, 
        \ARB_WRD_40M_FIXED[12]_net_1\, 
        \ARB_WRD_40M_FIXED[13]_net_1\, 
        \ARB_WRD_40M_FIXED[14]_net_1\, \GND\, \VCC\ : std_logic;

begin 


    \RECD_SER_WORD_RNO[5]\ : MX2
      port map(A => N_38, B => N_39, S => BIT_OS_SEL_5_0, Y => 
        \N_RECD_SER_WORD[5]\);
    
    \ARB_WRD_40M_FIXED[9]\ : DFN1C0
      port map(D => \Q[9]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[9]_net_1\);
    
    \ADJ_Q[4]\ : DFN1C0
      port map(D => \ADJ_Q[2]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[4]_net_1\);
    
    \ARB_BYTE[6]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[6]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[6]_net_1\);
    
    ADJ_SER_IN_F_1DEL : DFN1C0
      port map(D => \ADJ_SER_IN_F_0DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_F_1DEL\);
    
    \ARB_BYTE[0]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[0]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[0]_net_1\);
    
    \Q[11]\ : DFN1C0
      port map(D => \ADJ_Q[11]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[11]_net_1\);
    
    \ADJ_Q[8]\ : DFN1C0
      port map(D => \ADJ_Q[6]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[8]_net_1\);
    
    \ARB_BYTE_RNINJO11[10]\ : MX2
      port map(A => \ARB_BYTE[6]_net_1\, B => 
        \ARB_BYTE[10]_net_1\, S => BIT_OS_SEL_4(2), Y => N_23);
    
    \ADJ_Q[6]\ : DFN1C0
      port map(D => \ADJ_Q[4]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[6]_net_1\);
    
    \ADJ_Q[12]\ : DFN1C0
      port map(D => \ADJ_Q[10]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[12]_net_1\);
    
    \RECD_SER_WORD_RNO_1[0]\ : MX2
      port map(A => \ARB_BYTE[0]_net_1\, B => \ARB_BYTE[4]_net_1\, 
        S => BIT_OS_SEL_4(2), Y => N_17);
    
    \Q[1]\ : DFN1C0
      port map(D => \ADJ_Q[1]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[1]_net_1\);
    
    \ARB_BYTE[4]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[4]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[4]_net_1\);
    
    \ADJ_Q[2]\ : DFN1C0
      port map(D => \ADJ_Q[0]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[2]_net_1\);
    
    \RECD_SER_WORD_RNO_1[7]\ : MX2
      port map(A => \ARB_BYTE[10]_net_1\, B => 
        \ARB_BYTE[14]_net_1\, S => BIT_OS_SEL_6(2), Y => N_56);
    
    \RECD_SER_WORD[4]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[4]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_7(4));
    
    \Q[5]\ : DFN1C0
      port map(D => \ADJ_Q[5]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[5]_net_1\);
    
    \ADJ_Q[11]\ : DFN1C0
      port map(D => \ADJ_Q[9]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[11]_net_1\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \ARB_BYTE_RNIPLO11[11]\ : MX2
      port map(A => \ARB_BYTE[7]_net_1\, B => 
        \ARB_BYTE[11]_net_1\, S => BIT_OS_SEL_4(2), Y => N_24);
    
    \ADJ_Q[3]\ : DFN1C0
      port map(D => \ADJ_Q[1]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[3]_net_1\);
    
    \Q[10]\ : DFN1C0
      port map(D => \ADJ_Q[10]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[10]_net_1\);
    
    \ARB_BYTE_RNIEDH21[5]\ : MX2
      port map(A => \ARB_BYTE[5]_net_1\, B => \ARB_BYTE[9]_net_1\, 
        S => BIT_OS_SEL_4(2), Y => N_22);
    
    \ARB_WRD_40M_FIXED[6]\ : DFN1C0
      port map(D => \Q[6]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[6]_net_1\);
    
    \ARB_WRD_40M_FIXED[1]\ : DFN1C0
      port map(D => \Q[1]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[1]_net_1\);
    
    \ARB_BYTE_RNIRNO11[12]\ : MX2
      port map(A => \ARB_BYTE[8]_net_1\, B => 
        \ARB_BYTE[12]_net_1\, S => BIT_OS_SEL_4(2), Y => N_31);
    
    \RECD_SER_WORD[3]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[3]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_7(3));
    
    \RECD_SER_WORD[0]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[0]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_7(0));
    
    \RECD_SER_WORD_RNO[3]\ : MX2
      port map(A => N_36, B => N_37, S => BIT_OS_SEL_5_0, Y => 
        \N_RECD_SER_WORD[3]\);
    
    \Q[0]\ : DFN1C0
      port map(D => \ADJ_Q[0]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[0]_net_1\);
    
    \RECD_SER_WORD_RNO_0[7]\ : MX2
      port map(A => N_31, B => N_56, S => BIT_OS_SEL_6(1), Y => 
        N_64);
    
    \Q[7]\ : DFN1C0
      port map(D => \ADJ_Q[7]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[7]_net_1\);
    
    \ARB_BYTE[14]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[14]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[14]_net_1\);
    
    \ARB_WRD_40M_FIXED[2]\ : DFN1C0
      port map(D => \Q[2]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[2]_net_1\);
    
    \ARB_WRD_40M_FIXED[14]\ : DFN1C0
      port map(D => \Q[14]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[14]_net_1\);
    
    \RECD_SER_WORD_RNO[2]\ : MX2
      port map(A => N_35, B => N_36, S => BIT_OS_SEL_5_0, Y => 
        \N_RECD_SER_WORD[2]\);
    
    \ARB_BYTE_RNIVSK72[1]\ : MX2
      port map(A => N_18, B => N_20, S => BIT_OS_SEL_4(1), Y => 
        N_34);
    
    \ARB_BYTE[2]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[2]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[2]_net_1\);
    
    \ADJ_Q[7]\ : DFN1C0
      port map(D => \ADJ_Q[5]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[7]_net_1\);
    
    \ARB_BYTE[8]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[8]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[8]_net_1\);
    
    \ARB_BYTE_RNICBH21[4]\ : MX2
      port map(A => \ARB_BYTE[4]_net_1\, B => \ARB_BYTE[8]_net_1\, 
        S => BIT_OS_SEL_4(2), Y => N_21);
    
    \RECD_SER_WORD[5]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[5]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_7(5));
    
    \ARB_BYTE[12]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[12]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[12]_net_1\);
    
    \RECD_SER_WORD[1]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[1]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_7(1));
    
    \Q[3]\ : DFN1C0
      port map(D => \ADJ_Q[3]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[3]_net_1\);
    
    ADJ_SER_IN_F_0DEL : DFN1C0
      port map(D => ELK_IN_F, CLK => CCC_160M_ADJ, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_F_0DEL\);
    
    \RECD_SER_WORD_RNO[7]\ : MX2
      port map(A => N_40, B => N_64, S => BIT_OS_SEL_0, Y => 
        \N_RECD_SER_WORD[7]\);
    
    \RECD_SER_WORD_RNO[1]\ : MX2
      port map(A => N_34, B => N_35, S => BIT_OS_SEL_5_0, Y => 
        \N_RECD_SER_WORD[1]\);
    
    \ARB_WRD_40M_FIXED[4]\ : DFN1C0
      port map(D => \Q[4]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[4]_net_1\);
    
    \ARB_BYTE_RNIIDS62[10]\ : MX2
      port map(A => N_21, B => N_23, S => BIT_OS_SEL_4(1), Y => 
        N_37);
    
    \RECD_SER_WORD_RNO[0]\ : MX2
      port map(A => N_33, B => N_34, S => BIT_OS_SEL_5_0, Y => 
        \N_RECD_SER_WORD[0]\);
    
    \Q[6]\ : DFN1C0
      port map(D => \ADJ_Q[6]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[6]_net_1\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \ARB_WRD_40M_FIXED[8]\ : DFN1C0
      port map(D => \Q[8]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[8]_net_1\);
    
    \ARB_BYTE[11]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[11]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[11]_net_1\);
    
    \Q[9]\ : DFN1C0
      port map(D => \ADJ_Q[9]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[9]_net_1\);
    
    \ARB_BYTE_RNIUSR21[13]\ : MX2
      port map(A => \ARB_BYTE[9]_net_1\, B => 
        \ARB_BYTE[13]_net_1\, S => BIT_OS_SEL_5_2, Y => N_32);
    
    \Q[14]\ : DFN1C0
      port map(D => \ADJ_Q[14]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[14]_net_1\);
    
    \ARB_BYTE_RNI1Q362[10]\ : MX2
      port map(A => N_23, B => N_31, S => BIT_OS_SEL_4(1), Y => 
        N_39);
    
    ADJ_SER_IN_R_0DEL : DFN1C0
      port map(D => ELK_IN_R, CLK => CCC_160M_ADJ, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_R_0DEL\);
    
    \Q[13]\ : DFN1C0
      port map(D => \ADJ_Q[13]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[13]_net_1\);
    
    \ARB_BYTE[9]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[9]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[9]_net_1\);
    
    ADJ_SER_IN_R_1DEL : DFN1C0
      port map(D => \ADJ_SER_IN_R_0DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_R_1DEL\);
    
    \ARB_BYTE[10]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[10]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[10]_net_1\);
    
    \ADJ_Q[9]\ : DFN1C0
      port map(D => \ADJ_Q[7]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[9]_net_1\);
    
    \RECD_SER_WORD[7]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[7]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_7(7));
    
    \ARB_WRD_40M_FIXED[5]\ : DFN1C0
      port map(D => \Q[5]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[5]_net_1\);
    
    \ARB_WRD_40M_FIXED[12]\ : DFN1C0
      port map(D => \Q[12]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[12]_net_1\);
    
    \ARB_WRD_40M_FIXED[11]\ : DFN1C0
      port map(D => \Q[11]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[11]_net_1\);
    
    \ARB_BYTE_RNI75L72[3]\ : MX2
      port map(A => N_20, B => N_22, S => BIT_OS_SEL_4(1), Y => 
        N_36);
    
    \ARB_WRD_40M_FIXED[0]\ : DFN1C0
      port map(D => \Q[0]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[0]_net_1\);
    
    \ADJ_Q[10]\ : DFN1C0
      port map(D => \ADJ_Q[8]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[10]_net_1\);
    
    \Q[2]\ : DFN1C0
      port map(D => \ADJ_Q[2]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[2]_net_1\);
    
    \ADJ_Q[1]\ : DFN1C0
      port map(D => \ADJ_SER_IN_F_1DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[1]_net_1\);
    
    \RECD_SER_WORD[6]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[6]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_7(6));
    
    \RECD_SER_WORD[2]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[2]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_7(2));
    
    \ADJ_Q[13]\ : DFN1C0
      port map(D => \ADJ_Q[11]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[13]_net_1\);
    
    \Q[8]\ : DFN1C0
      port map(D => \ADJ_Q[8]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[8]_net_1\);
    
    \ARB_BYTE[5]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[5]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[5]_net_1\);
    
    \ADJ_Q[14]\ : DFN1C0
      port map(D => \ADJ_Q[12]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[14]_net_1\);
    
    \RECD_SER_WORD_RNO[4]\ : MX2
      port map(A => N_37, B => N_38, S => BIT_OS_SEL_5_0, Y => 
        \N_RECD_SER_WORD[4]\);
    
    \Q[12]\ : DFN1C0
      port map(D => \ADJ_Q[12]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[12]_net_1\);
    
    \ARB_BYTE_RNI87H21[2]\ : MX2
      port map(A => \ARB_BYTE[2]_net_1\, B => \ARB_BYTE[6]_net_1\, 
        S => BIT_OS_SEL_4(2), Y => N_19);
    
    \ARB_BYTE[13]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[13]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[13]_net_1\);
    
    \ARB_WRD_40M_FIXED[3]\ : DFN1C0
      port map(D => \Q[3]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[3]_net_1\);
    
    \ARB_BYTE[7]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[7]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[7]_net_1\);
    
    \RECD_SER_WORD_RNO_0[0]\ : MX2
      port map(A => N_17, B => N_19, S => BIT_OS_SEL_4(1), Y => 
        N_33);
    
    \ARB_BYTE_RNIA9H21[3]\ : MX2
      port map(A => \ARB_BYTE[3]_net_1\, B => \ARB_BYTE[7]_net_1\, 
        S => BIT_OS_SEL_4(2), Y => N_20);
    
    \Q[4]\ : DFN1C0
      port map(D => \ADJ_Q[4]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[4]_net_1\);
    
    \ARB_WRD_40M_FIXED[7]\ : DFN1C0
      port map(D => \Q[7]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[7]_net_1\);
    
    \RECD_SER_WORD_RNO[6]\ : MX2
      port map(A => N_39, B => N_40, S => BIT_OS_SEL_5_0, Y => 
        \N_RECD_SER_WORD[6]\);
    
    \ARB_BYTE[3]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[3]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[3]_net_1\);
    
    \ARB_BYTE_RNI65H21[1]\ : MX2
      port map(A => \ARB_BYTE[1]_net_1\, B => \ARB_BYTE[5]_net_1\, 
        S => BIT_OS_SEL_4(2), Y => N_18);
    
    \ARB_BYTE_RNI61772[13]\ : MX2
      port map(A => N_24, B => N_32, S => BIT_OS_SEL_4(1), Y => 
        N_40);
    
    \ADJ_Q[5]\ : DFN1C0
      port map(D => \ADJ_Q[3]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[5]_net_1\);
    
    \ARB_BYTE[1]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[1]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[1]_net_1\);
    
    \ARB_WRD_40M_FIXED[13]\ : DFN1C0
      port map(D => \Q[13]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[13]_net_1\);
    
    \ADJ_Q[0]\ : DFN1C0
      port map(D => \ADJ_SER_IN_R_1DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[0]_net_1\);
    
    \ARB_BYTE_RNIMHS62[11]\ : MX2
      port map(A => N_22, B => N_24, S => BIT_OS_SEL_4(1), Y => 
        N_38);
    
    \ARB_WRD_40M_FIXED[10]\ : DFN1C0
      port map(D => \Q[10]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[10]_net_1\);
    
    \ARB_BYTE_RNI31L72[2]\ : MX2
      port map(A => N_19, B => N_21, S => BIT_OS_SEL_4(1), Y => 
        N_35);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SER320M_3_34_7 is

    port( ELK_TX_DAT                 : in    std_logic_vector(7 downto 0);
          MASTER_SALT_POR_B_i_0_i_10 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_14 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_13 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_2  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_8  : in    std_logic;
          ELK_OUT_R                  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_12 : in    std_logic;
          ELK_OUT_F                  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_11 : in    std_logic;
          CCC_160M_FXD               : in    std_logic;
          CLK_40M_GL                 : in    std_logic
        );

end SER320M_3_34_7;

architecture DEF_ARCH of SER320M_3_34_7 is 

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \N_SER_CMD_WORD_R[0]\, \START_RISE\, 
        \N_SER_CMD_WORD_F[0]\, \N_SER_CMD_WORD_R[3]\, 
        \SER_CMD_WORD_R[2]_net_1\, \N_SER_CMD_WORD_R[2]\, 
        \SER_CMD_WORD_R[1]_net_1\, \N_SER_CMD_WORD_R[1]\, 
        \SER_CMD_WORD_R[0]_net_1\, \N_SER_CMD_WORD_F[3]\, 
        \SER_CMD_WORD_F[2]_net_1\, \N_SER_CMD_WORD_F[2]\, 
        \SER_CMD_WORD_F[1]_net_1\, \N_SER_CMD_WORD_F[1]\, 
        \SER_CMD_WORD_F[0]_net_1\, N_START_RISE, 
        \CLK40M_GEN_DEL0\, \SER_OUT_FI\, \SER_OUT_RI\, 
        \SER_CMD_WORD_F[3]_net_1\, \SER_CMD_WORD_R[3]_net_1\, 
        \GND\, \VCC\ : std_logic;

begin 


    SER_OUT_FI : DFN1C0
      port map(D => \SER_CMD_WORD_F[3]_net_1\, CLK => 
        CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_13, Q => 
        \SER_OUT_FI\);
    
    \SER_CMD_WORD_F[3]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[3]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_14, Q => 
        \SER_CMD_WORD_F[3]_net_1\);
    
    \SER_CMD_WORD_R[1]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[1]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_10, Q => 
        \SER_CMD_WORD_R[1]_net_1\);
    
    \SER_CMD_WORD_R[2]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[2]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_11, Q => 
        \SER_CMD_WORD_R[2]_net_1\);
    
    \SER_CMD_WORD_R_RNO[3]\ : MX2
      port map(A => \SER_CMD_WORD_R[2]_net_1\, B => ELK_TX_DAT(7), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_R[3]\);
    
    \SER_CMD_WORD_R_RNO[0]\ : NOR2B
      port map(A => \START_RISE\, B => ELK_TX_DAT(1), Y => 
        \N_SER_CMD_WORD_R[0]\);
    
    \SER_CMD_WORD_F[0]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[0]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_14, Q => 
        \SER_CMD_WORD_F[0]_net_1\);
    
    \SER_CMD_WORD_R_RNO[1]\ : MX2
      port map(A => \SER_CMD_WORD_R[0]_net_1\, B => ELK_TX_DAT(3), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_R[1]\);
    
    \SER_CMD_WORD_F_RNO[2]\ : MX2
      port map(A => \SER_CMD_WORD_F[1]_net_1\, B => ELK_TX_DAT(4), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_F[2]\);
    
    \SER_CMD_WORD_F_RNO[3]\ : MX2
      port map(A => \SER_CMD_WORD_F[2]_net_1\, B => ELK_TX_DAT(6), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_F[3]\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    CLK40M_GEN_DEL0 : DFN1C0
      port map(D => CLK_40M_GL, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_11, Q => \CLK40M_GEN_DEL0\);
    
    SER_OUT_RI : DFN1C0
      port map(D => \SER_CMD_WORD_R[3]_net_1\, CLK => 
        CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_13, Q => 
        \SER_OUT_RI\);
    
    \SER_CMD_WORD_F[2]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[2]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_14, Q => 
        \SER_CMD_WORD_F[2]_net_1\);
    
    \SER_CMD_WORD_F_RNO[1]\ : MX2
      port map(A => \SER_CMD_WORD_F[0]_net_1\, B => ELK_TX_DAT(2), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_F[1]\);
    
    \SER_CMD_WORD_R[0]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[0]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_10, Q => 
        \SER_CMD_WORD_R[0]_net_1\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    START_RISE : DFN1C0
      port map(D => N_START_RISE, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_2, Q => \START_RISE\);
    
    \SER_CMD_WORD_R[3]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[3]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_11, Q => 
        \SER_CMD_WORD_R[3]_net_1\);
    
    \SER_CMD_WORD_F_RNO[0]\ : NOR2B
      port map(A => \START_RISE\, B => ELK_TX_DAT(0), Y => 
        \N_SER_CMD_WORD_F[0]\);
    
    SER_OUT_RDEL : DFN1C0
      port map(D => \SER_OUT_RI\, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_8, Q => ELK_OUT_R);
    
    \SER_CMD_WORD_F[1]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[1]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_14, Q => 
        \SER_CMD_WORD_F[1]_net_1\);
    
    START_RISE_RNO : NOR2B
      port map(A => \CLK40M_GEN_DEL0\, B => CLK_40M_GL, Y => 
        N_START_RISE);
    
    \SER_CMD_WORD_R_RNO[2]\ : MX2
      port map(A => \SER_CMD_WORD_R[1]_net_1\, B => ELK_TX_DAT(5), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_R[2]\);
    
    SER_OUT_FDEL : DFN1C0
      port map(D => \SER_OUT_FI\, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_12, Q => ELK_OUT_F);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity DDR_BIDIR_LVDS_DUAL_CLK_7 is

    port( DCB_SALT_SEL_c_i : in    std_logic;
          ELK7_DAT_P       : inout std_logic := 'Z';
          ELK7_DAT_N       : inout std_logic := 'Z';
          ELK_OUT_R        : in    std_logic;
          ELK_OUT_F        : in    std_logic;
          CCC_160M_FXD     : in    std_logic;
          CCC_160M_ADJ     : in    std_logic;
          ELK_IN_DDR_R     : out   std_logic;
          ELK_IN_DDR_F     : out   std_logic
        );

end DDR_BIDIR_LVDS_DUAL_CLK_7;

architecture DEF_ARCH of DDR_BIDIR_LVDS_DUAL_CLK_7 is 

  component DDR_REG
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          QR  : out   std_logic;
          QF  : out   std_logic
        );
  end component;

  component DDR_OUT
    port( DR  : in    std_logic := 'U';
          DF  : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component BIBUF_LVDS
    port( PADP : inout   std_logic;
          PADN : inout   std_logic;
          D    : in    std_logic := 'U';
          E    : in    std_logic := 'U';
          Y    : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal DDR_BIDIR_LVDS_DUAL_CLK_7_GND, BIBUF_LVDS_0_Y, 
        DDR_OUT_0_Q, \VCC\ : std_logic;

begin 


    DDR_REG_0 : DDR_REG
      port map(D => BIBUF_LVDS_0_Y, CLK => CCC_160M_ADJ, CLR => 
        DDR_BIDIR_LVDS_DUAL_CLK_7_GND, QR => ELK_IN_DDR_R, QF => 
        ELK_IN_DDR_F);
    
    DDR_OUT_0 : DDR_OUT
      port map(DR => ELK_OUT_R, DF => ELK_OUT_F, CLK => 
        CCC_160M_FXD, CLR => DDR_BIDIR_LVDS_DUAL_CLK_7_GND, Q => 
        DDR_OUT_0_Q);
    
    BIBUF_LVDS_0 : BIBUF_LVDS
      port map(PADP => ELK7_DAT_P, PADN => ELK7_DAT_N, D => 
        DDR_OUT_0_Q, E => DCB_SALT_SEL_c_i, Y => BIBUF_LVDS_0_Y);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    GND_i : GND
      port map(Y => DDR_BIDIR_LVDS_DUAL_CLK_7_GND);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SYNC_DAT_SEL_7 is

    port( ELK_TX_DAT                : out   std_logic_vector(7 downto 0);
          PATT_ELK_DAT_7            : in    std_logic_vector(7 downto 0);
          OP_MODE_c_4_0             : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_3 : in    std_logic;
          CLK_40M_GL                : in    std_logic
        );

end SYNC_DAT_SEL_7;

architecture DEF_ARCH of SYNC_DAT_SEL_7 is 

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \N_SERDAT[0]\, \N_SERDAT[1]\, \N_SERDAT[2]\, 
        \N_SERDAT[3]\, \N_SERDAT[4]\, \N_SERDAT[5]\, 
        \N_SERDAT[6]\, \N_SERDAT[7]\, \GND\, \VCC\ : std_logic;

begin 


    \SERDAT_RNO[4]\ : NOR2A
      port map(A => PATT_ELK_DAT_7(4), B => OP_MODE_c_4_0, Y => 
        \N_SERDAT[4]\);
    
    \SERDAT_RNO[0]\ : NOR2A
      port map(A => PATT_ELK_DAT_7(0), B => OP_MODE_c_4_0, Y => 
        \N_SERDAT[0]\);
    
    \SERDAT[6]\ : DFN1C0
      port map(D => \N_SERDAT[6]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_3, Q => ELK_TX_DAT(6));
    
    \SERDAT[4]\ : DFN1C0
      port map(D => \N_SERDAT[4]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_3, Q => ELK_TX_DAT(4));
    
    \SERDAT_RNO[7]\ : OR2
      port map(A => PATT_ELK_DAT_7(7), B => OP_MODE_c_4_0, Y => 
        \N_SERDAT[7]\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \SERDAT_RNO[3]\ : OR2
      port map(A => PATT_ELK_DAT_7(3), B => OP_MODE_c_4_0, Y => 
        \N_SERDAT[3]\);
    
    \SERDAT_RNO[2]\ : OR2
      port map(A => PATT_ELK_DAT_7(2), B => OP_MODE_c_4_0, Y => 
        \N_SERDAT[2]\);
    
    \SERDAT[5]\ : DFN1C0
      port map(D => \N_SERDAT[5]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_3, Q => ELK_TX_DAT(5));
    
    \SERDAT[7]\ : DFN1C0
      port map(D => \N_SERDAT[7]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_3, Q => ELK_TX_DAT(7));
    
    GND_i : GND
      port map(Y => \GND\);
    
    \SERDAT_RNO[5]\ : NOR2A
      port map(A => PATT_ELK_DAT_7(5), B => OP_MODE_c_4_0, Y => 
        \N_SERDAT[5]\);
    
    \SERDAT[0]\ : DFN1C0
      port map(D => \N_SERDAT[0]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_3, Q => ELK_TX_DAT(0));
    
    \SERDAT_RNO[6]\ : NOR2A
      port map(A => PATT_ELK_DAT_7(6), B => OP_MODE_c_4_0, Y => 
        \N_SERDAT[6]\);
    
    \SERDAT[1]\ : DFN1C0
      port map(D => \N_SERDAT[1]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_3, Q => ELK_TX_DAT(1));
    
    \SERDAT_RNO[1]\ : OR2
      port map(A => PATT_ELK_DAT_7(1), B => OP_MODE_c_4_0, Y => 
        \N_SERDAT[1]\);
    
    \SERDAT[3]\ : DFN1C0
      port map(D => \N_SERDAT[3]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_3, Q => ELK_TX_DAT(3));
    
    \SERDAT[2]\ : DFN1C0
      port map(D => \N_SERDAT[2]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_3, Q => ELK_TX_DAT(2));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity ELINK_SLAVE_15_2 is

    port( BIT_OS_SEL_4               : in    std_logic_vector(2 downto 1);
          BIT_OS_SEL_6               : in    std_logic_vector(2 downto 1);
          BIT_OS_SEL_5_2             : in    std_logic;
          BIT_OS_SEL_5_0             : in    std_logic;
          BIT_OS_SEL_0               : in    std_logic;
          ELK_RX_SER_WORD_7          : out   std_logic_vector(7 downto 0);
          OP_MODE_c_4_0              : in    std_logic;
          PATT_ELK_DAT_7             : in    std_logic_vector(7 downto 0);
          MASTER_DCB_POR_B_i_0_i     : in    std_logic;
          ELK7_DAT_N                 : inout std_logic := 'Z';
          ELK7_DAT_P                 : inout std_logic := 'Z';
          DCB_SALT_SEL_c_i           : in    std_logic;
          CCC_160M_FXD               : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_11 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_12 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_8  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_2  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_13 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_14 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_10 : in    std_logic;
          CLK_40M_GL                 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_3  : in    std_logic;
          DEV_RST_B_c_1              : in    std_logic;
          CCC_160M_ADJ               : in    std_logic
        );

end ELINK_SLAVE_15_2;

architecture DEF_ARCH of ELINK_SLAVE_15_2 is 

  component SLAVE_DES320S_1_17_5
    port( ELK_RX_SER_WORD_7      : out   std_logic_vector(7 downto 0);
          BIT_OS_SEL_0           : in    std_logic := 'U';
          BIT_OS_SEL_5_2         : in    std_logic := 'U';
          BIT_OS_SEL_5_0         : in    std_logic := 'U';
          BIT_OS_SEL_6           : in    std_logic_vector(2 downto 1) := (others => 'U');
          BIT_OS_SEL_4           : in    std_logic_vector(2 downto 1) := (others => 'U');
          CLK_40M_GL             : in    std_logic := 'U';
          CCC_160M_FXD           : in    std_logic := 'U';
          ELK_IN_R               : in    std_logic := 'U';
          ELK_IN_F               : in    std_logic := 'U';
          MASTER_DCB_POR_B_i_0_i : in    std_logic := 'U';
          CCC_160M_ADJ           : in    std_logic := 'U'
        );
  end component;

  component SER320M_3_34_7
    port( ELK_TX_DAT                 : in    std_logic_vector(7 downto 0) := (others => 'U');
          MASTER_SALT_POR_B_i_0_i_10 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_14 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_13 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_2  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_8  : in    std_logic := 'U';
          ELK_OUT_R                  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_12 : in    std_logic := 'U';
          ELK_OUT_F                  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_11 : in    std_logic := 'U';
          CCC_160M_FXD               : in    std_logic := 'U';
          CLK_40M_GL                 : in    std_logic := 'U'
        );
  end component;

  component DDR_BIDIR_LVDS_DUAL_CLK_7
    port( DCB_SALT_SEL_c_i : in    std_logic := 'U';
          ELK7_DAT_P       : inout   std_logic;
          ELK7_DAT_N       : inout   std_logic;
          ELK_OUT_R        : in    std_logic := 'U';
          ELK_OUT_F        : in    std_logic := 'U';
          CCC_160M_FXD     : in    std_logic := 'U';
          CCC_160M_ADJ     : in    std_logic := 'U';
          ELK_IN_DDR_R     : out   std_logic;
          ELK_IN_DDR_F     : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component SYNC_DAT_SEL_7
    port( ELK_TX_DAT                : out   std_logic_vector(7 downto 0);
          PATT_ELK_DAT_7            : in    std_logic_vector(7 downto 0) := (others => 'U');
          OP_MODE_c_4_0             : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_3 : in    std_logic := 'U';
          CLK_40M_GL                : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \ELK_IN_F\, ELK_IN_DDR_F, \ELK_IN_R\, ELK_IN_DDR_R, 
        \ELK_TX_DAT[0]\, \ELK_TX_DAT[1]\, \ELK_TX_DAT[2]\, 
        \ELK_TX_DAT[3]\, \ELK_TX_DAT[4]\, \ELK_TX_DAT[5]\, 
        \ELK_TX_DAT[6]\, \ELK_TX_DAT[7]\, ELK_OUT_R, ELK_OUT_F, 
        \GND\, \VCC\ : std_logic;

    for all : SLAVE_DES320S_1_17_5
	Use entity work.SLAVE_DES320S_1_17_5(DEF_ARCH);
    for all : SER320M_3_34_7
	Use entity work.SER320M_3_34_7(DEF_ARCH);
    for all : DDR_BIDIR_LVDS_DUAL_CLK_7
	Use entity work.DDR_BIDIR_LVDS_DUAL_CLK_7(DEF_ARCH);
    for all : SYNC_DAT_SEL_7
	Use entity work.SYNC_DAT_SEL_7(DEF_ARCH);
begin 


    U_SLAVE_1ELK : SLAVE_DES320S_1_17_5
      port map(ELK_RX_SER_WORD_7(7) => ELK_RX_SER_WORD_7(7), 
        ELK_RX_SER_WORD_7(6) => ELK_RX_SER_WORD_7(6), 
        ELK_RX_SER_WORD_7(5) => ELK_RX_SER_WORD_7(5), 
        ELK_RX_SER_WORD_7(4) => ELK_RX_SER_WORD_7(4), 
        ELK_RX_SER_WORD_7(3) => ELK_RX_SER_WORD_7(3), 
        ELK_RX_SER_WORD_7(2) => ELK_RX_SER_WORD_7(2), 
        ELK_RX_SER_WORD_7(1) => ELK_RX_SER_WORD_7(1), 
        ELK_RX_SER_WORD_7(0) => ELK_RX_SER_WORD_7(0), 
        BIT_OS_SEL_0 => BIT_OS_SEL_0, BIT_OS_SEL_5_2 => 
        BIT_OS_SEL_5_2, BIT_OS_SEL_5_0 => BIT_OS_SEL_5_0, 
        BIT_OS_SEL_6(2) => BIT_OS_SEL_6(2), BIT_OS_SEL_6(1) => 
        BIT_OS_SEL_6(1), BIT_OS_SEL_4(2) => BIT_OS_SEL_4(2), 
        BIT_OS_SEL_4(1) => BIT_OS_SEL_4(1), CLK_40M_GL => 
        CLK_40M_GL, CCC_160M_FXD => CCC_160M_FXD, ELK_IN_R => 
        \ELK_IN_R\, ELK_IN_F => \ELK_IN_F\, 
        MASTER_DCB_POR_B_i_0_i => MASTER_DCB_POR_B_i_0_i, 
        CCC_160M_ADJ => CCC_160M_ADJ);
    
    U_ELK1_CMD_TX : SER320M_3_34_7
      port map(ELK_TX_DAT(7) => \ELK_TX_DAT[7]\, ELK_TX_DAT(6)
         => \ELK_TX_DAT[6]\, ELK_TX_DAT(5) => \ELK_TX_DAT[5]\, 
        ELK_TX_DAT(4) => \ELK_TX_DAT[4]\, ELK_TX_DAT(3) => 
        \ELK_TX_DAT[3]\, ELK_TX_DAT(2) => \ELK_TX_DAT[2]\, 
        ELK_TX_DAT(1) => \ELK_TX_DAT[1]\, ELK_TX_DAT(0) => 
        \ELK_TX_DAT[0]\, MASTER_SALT_POR_B_i_0_i_10 => 
        MASTER_SALT_POR_B_i_0_i_10, MASTER_SALT_POR_B_i_0_i_14
         => MASTER_SALT_POR_B_i_0_i_14, 
        MASTER_SALT_POR_B_i_0_i_13 => MASTER_SALT_POR_B_i_0_i_13, 
        MASTER_SALT_POR_B_i_0_i_2 => MASTER_SALT_POR_B_i_0_i_2, 
        MASTER_SALT_POR_B_i_0_i_8 => MASTER_SALT_POR_B_i_0_i_8, 
        ELK_OUT_R => ELK_OUT_R, MASTER_SALT_POR_B_i_0_i_12 => 
        MASTER_SALT_POR_B_i_0_i_12, ELK_OUT_F => ELK_OUT_F, 
        MASTER_SALT_POR_B_i_0_i_11 => MASTER_SALT_POR_B_i_0_i_11, 
        CCC_160M_FXD => CCC_160M_FXD, CLK_40M_GL => CLK_40M_GL);
    
    U_DDR_ELK1 : DDR_BIDIR_LVDS_DUAL_CLK_7
      port map(DCB_SALT_SEL_c_i => DCB_SALT_SEL_c_i, ELK7_DAT_P
         => ELK7_DAT_P, ELK7_DAT_N => ELK7_DAT_N, ELK_OUT_R => 
        ELK_OUT_R, ELK_OUT_F => ELK_OUT_F, CCC_160M_FXD => 
        CCC_160M_FXD, CCC_160M_ADJ => CCC_160M_ADJ, ELK_IN_DDR_R
         => ELK_IN_DDR_R, ELK_IN_DDR_F => ELK_IN_DDR_F);
    
    ELK_IN_F : DFN1C0
      port map(D => ELK_IN_DDR_F, CLK => CCC_160M_ADJ, CLR => 
        DEV_RST_B_c_1, Q => \ELK_IN_F\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    U_ELK1_SERDAT_SOURCE : SYNC_DAT_SEL_7
      port map(ELK_TX_DAT(7) => \ELK_TX_DAT[7]\, ELK_TX_DAT(6)
         => \ELK_TX_DAT[6]\, ELK_TX_DAT(5) => \ELK_TX_DAT[5]\, 
        ELK_TX_DAT(4) => \ELK_TX_DAT[4]\, ELK_TX_DAT(3) => 
        \ELK_TX_DAT[3]\, ELK_TX_DAT(2) => \ELK_TX_DAT[2]\, 
        ELK_TX_DAT(1) => \ELK_TX_DAT[1]\, ELK_TX_DAT(0) => 
        \ELK_TX_DAT[0]\, PATT_ELK_DAT_7(7) => PATT_ELK_DAT_7(7), 
        PATT_ELK_DAT_7(6) => PATT_ELK_DAT_7(6), PATT_ELK_DAT_7(5)
         => PATT_ELK_DAT_7(5), PATT_ELK_DAT_7(4) => 
        PATT_ELK_DAT_7(4), PATT_ELK_DAT_7(3) => PATT_ELK_DAT_7(3), 
        PATT_ELK_DAT_7(2) => PATT_ELK_DAT_7(2), PATT_ELK_DAT_7(1)
         => PATT_ELK_DAT_7(1), PATT_ELK_DAT_7(0) => 
        PATT_ELK_DAT_7(0), OP_MODE_c_4_0 => OP_MODE_c_4_0, 
        MASTER_SALT_POR_B_i_0_i_3 => MASTER_SALT_POR_B_i_0_i_3, 
        CLK_40M_GL => CLK_40M_GL);
    
    ELK_IN_R : DFN1C0
      port map(D => ELK_IN_DDR_R, CLK => CCC_160M_ADJ, CLR => 
        DEV_RST_B_c_1, Q => \ELK_IN_R\);
    
    GND_i : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SLAVE_DES320S_1_17_12 is

    port( ELK_RX_SER_WORD_14     : out   std_logic_vector(7 downto 0);
          BIT_OS_SEL_4           : in    std_logic_vector(1 downto 0);
          BIT_OS_SEL_3_0         : in    std_logic;
          BIT_OS_SEL_5_0         : in    std_logic;
          BIT_OS_SEL_2           : in    std_logic_vector(2 downto 1);
          CLK_40M_GL             : in    std_logic;
          CCC_160M_FXD           : in    std_logic;
          ELK_IN_R               : in    std_logic;
          ELK_IN_F               : in    std_logic;
          MASTER_DCB_POR_B_i_0_i : in    std_logic;
          CCC_160M_ADJ           : in    std_logic
        );

end SLAVE_DES320S_1_17_12;

architecture DEF_ARCH of SLAVE_DES320S_1_17_12 is 

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal N_17, \ARB_BYTE[0]_net_1\, \ARB_BYTE[4]_net_1\, N_18, 
        \ARB_BYTE[1]_net_1\, \ARB_BYTE[5]_net_1\, N_19, 
        \ARB_BYTE[2]_net_1\, \ARB_BYTE[6]_net_1\, N_20, 
        \ARB_BYTE[3]_net_1\, \ARB_BYTE[7]_net_1\, N_21, 
        \ARB_BYTE[8]_net_1\, N_22, \ARB_BYTE[9]_net_1\, N_23, 
        \ARB_BYTE[10]_net_1\, N_24, \ARB_BYTE[11]_net_1\, N_31, 
        \ARB_BYTE[12]_net_1\, N_32, \ARB_BYTE[13]_net_1\, N_33, 
        N_34, N_35, N_36, N_37, N_38, N_39, N_40, N_56, 
        \ARB_BYTE[14]_net_1\, N_64, \N_RECD_SER_WORD[0]\, 
        \N_RECD_SER_WORD[1]\, \N_RECD_SER_WORD[2]\, 
        \N_RECD_SER_WORD[3]\, \N_RECD_SER_WORD[4]\, 
        \N_RECD_SER_WORD[5]\, \N_RECD_SER_WORD[6]\, 
        \N_RECD_SER_WORD[7]\, \ADJ_SER_IN_F_0DEL\, 
        \ADJ_SER_IN_R_0DEL\, \ADJ_SER_IN_F_1DEL\, 
        \ADJ_SER_IN_R_1DEL\, \Q[0]_net_1\, \ADJ_Q[0]_net_1\, 
        \Q[1]_net_1\, \ADJ_Q[1]_net_1\, \Q[2]_net_1\, 
        \ADJ_Q[2]_net_1\, \Q[3]_net_1\, \ADJ_Q[3]_net_1\, 
        \Q[4]_net_1\, \ADJ_Q[4]_net_1\, \Q[5]_net_1\, 
        \ADJ_Q[5]_net_1\, \Q[6]_net_1\, \ADJ_Q[6]_net_1\, 
        \Q[7]_net_1\, \ADJ_Q[7]_net_1\, \Q[8]_net_1\, 
        \ADJ_Q[8]_net_1\, \Q[9]_net_1\, \ADJ_Q[9]_net_1\, 
        \Q[10]_net_1\, \ADJ_Q[10]_net_1\, \Q[11]_net_1\, 
        \ADJ_Q[11]_net_1\, \Q[12]_net_1\, \ADJ_Q[12]_net_1\, 
        \Q[13]_net_1\, \ADJ_Q[13]_net_1\, \Q[14]_net_1\, 
        \ADJ_Q[14]_net_1\, \ARB_WRD_40M_FIXED[0]_net_1\, 
        \ARB_WRD_40M_FIXED[1]_net_1\, 
        \ARB_WRD_40M_FIXED[2]_net_1\, 
        \ARB_WRD_40M_FIXED[3]_net_1\, 
        \ARB_WRD_40M_FIXED[4]_net_1\, 
        \ARB_WRD_40M_FIXED[5]_net_1\, 
        \ARB_WRD_40M_FIXED[6]_net_1\, 
        \ARB_WRD_40M_FIXED[7]_net_1\, 
        \ARB_WRD_40M_FIXED[8]_net_1\, 
        \ARB_WRD_40M_FIXED[9]_net_1\, 
        \ARB_WRD_40M_FIXED[10]_net_1\, 
        \ARB_WRD_40M_FIXED[11]_net_1\, 
        \ARB_WRD_40M_FIXED[12]_net_1\, 
        \ARB_WRD_40M_FIXED[13]_net_1\, 
        \ARB_WRD_40M_FIXED[14]_net_1\, \GND\, \VCC\ : std_logic;

begin 


    \RECD_SER_WORD_RNO[5]\ : MX2
      port map(A => N_38, B => N_39, S => BIT_OS_SEL_4(0), Y => 
        \N_RECD_SER_WORD[5]\);
    
    \ARB_WRD_40M_FIXED[9]\ : DFN1C0
      port map(D => \Q[9]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[9]_net_1\);
    
    \ARB_BYTE_RNI0KLR[1]\ : MX2
      port map(A => \ARB_BYTE[1]_net_1\, B => \ARB_BYTE[5]_net_1\, 
        S => BIT_OS_SEL_2(2), Y => N_18);
    
    \ADJ_Q[4]\ : DFN1C0
      port map(D => \ADJ_Q[2]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[4]_net_1\);
    
    \ARB_BYTE[6]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[6]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[6]_net_1\);
    
    ADJ_SER_IN_F_1DEL : DFN1C0
      port map(D => \ADJ_SER_IN_F_0DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_F_1DEL\);
    
    \ARB_BYTE[0]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[0]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[0]_net_1\);
    
    \Q[11]\ : DFN1C0
      port map(D => \ADJ_Q[11]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[11]_net_1\);
    
    \ADJ_Q[8]\ : DFN1C0
      port map(D => \ADJ_Q[6]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[8]_net_1\);
    
    \ADJ_Q[6]\ : DFN1C0
      port map(D => \ADJ_Q[4]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[6]_net_1\);
    
    \ARB_BYTE_RNI6QLR[4]\ : MX2
      port map(A => \ARB_BYTE[4]_net_1\, B => \ARB_BYTE[8]_net_1\, 
        S => BIT_OS_SEL_2(2), Y => N_21);
    
    \ADJ_Q[12]\ : DFN1C0
      port map(D => \ADJ_Q[10]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[12]_net_1\);
    
    \RECD_SER_WORD_RNO_1[0]\ : MX2
      port map(A => \ARB_BYTE[0]_net_1\, B => \ARB_BYTE[4]_net_1\, 
        S => BIT_OS_SEL_2(2), Y => N_17);
    
    \Q[1]\ : DFN1C0
      port map(D => \ADJ_Q[1]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[1]_net_1\);
    
    \ARB_BYTE[4]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[4]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[4]_net_1\);
    
    \ADJ_Q[2]\ : DFN1C0
      port map(D => \ADJ_Q[0]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[2]_net_1\);
    
    \RECD_SER_WORD_RNO_1[7]\ : MX2
      port map(A => \ARB_BYTE[10]_net_1\, B => 
        \ARB_BYTE[14]_net_1\, S => BIT_OS_SEL_5_0, Y => N_56);
    
    \RECD_SER_WORD[4]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[4]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_14(4));
    
    \Q[5]\ : DFN1C0
      port map(D => \ADJ_Q[5]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[5]_net_1\);
    
    \ADJ_Q[11]\ : DFN1C0
      port map(D => \ADJ_Q[9]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[11]_net_1\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \ADJ_Q[3]\ : DFN1C0
      port map(D => \ADJ_Q[1]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[3]_net_1\);
    
    \Q[10]\ : DFN1C0
      port map(D => \ADJ_Q[10]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[10]_net_1\);
    
    \ARB_WRD_40M_FIXED[6]\ : DFN1C0
      port map(D => \Q[6]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[6]_net_1\);
    
    \ARB_WRD_40M_FIXED[1]\ : DFN1C0
      port map(D => \Q[1]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[1]_net_1\);
    
    \RECD_SER_WORD[3]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[3]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_14(3));
    
    \RECD_SER_WORD[0]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[0]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_14(0));
    
    \ARB_BYTE_RNINM7G[13]\ : MX2
      port map(A => \ARB_BYTE[9]_net_1\, B => 
        \ARB_BYTE[13]_net_1\, S => BIT_OS_SEL_2(2), Y => N_32);
    
    \RECD_SER_WORD_RNO[3]\ : MX2
      port map(A => N_36, B => N_37, S => BIT_OS_SEL_4(0), Y => 
        \N_RECD_SER_WORD[3]\);
    
    \Q[0]\ : DFN1C0
      port map(D => \ADJ_Q[0]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[0]_net_1\);
    
    \RECD_SER_WORD_RNO_0[7]\ : MX2
      port map(A => N_31, B => N_56, S => BIT_OS_SEL_4(1), Y => 
        N_64);
    
    \Q[7]\ : DFN1C0
      port map(D => \ADJ_Q[7]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[7]_net_1\);
    
    \ARB_BYTE[14]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[14]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[14]_net_1\);
    
    \ARB_WRD_40M_FIXED[2]\ : DFN1C0
      port map(D => \Q[2]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[2]_net_1\);
    
    \ARB_WRD_40M_FIXED[14]\ : DFN1C0
      port map(D => \Q[14]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[14]_net_1\);
    
    \RECD_SER_WORD_RNO[2]\ : MX2
      port map(A => N_35, B => N_36, S => BIT_OS_SEL_4(0), Y => 
        \N_RECD_SER_WORD[2]\);
    
    \ARB_BYTE[2]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[2]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[2]_net_1\);
    
    \ARB_BYTE_RNILONN1[2]\ : MX2
      port map(A => N_19, B => N_21, S => BIT_OS_SEL_2(1), Y => 
        N_35);
    
    \ADJ_Q[7]\ : DFN1C0
      port map(D => \ADJ_Q[5]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[7]_net_1\);
    
    \ARB_BYTE[8]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[8]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[8]_net_1\);
    
    \ARB_BYTE_RNIHG7G[10]\ : MX2
      port map(A => \ARB_BYTE[6]_net_1\, B => 
        \ARB_BYTE[10]_net_1\, S => BIT_OS_SEL_2(2), Y => N_23);
    
    \RECD_SER_WORD[5]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[5]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_14(5));
    
    \ARB_BYTE[12]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[12]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[12]_net_1\);
    
    \RECD_SER_WORD[1]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[1]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_14(1));
    
    \Q[3]\ : DFN1C0
      port map(D => \ADJ_Q[3]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[3]_net_1\);
    
    ADJ_SER_IN_F_0DEL : DFN1C0
      port map(D => ELK_IN_F, CLK => CCC_160M_ADJ, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_F_0DEL\);
    
    \RECD_SER_WORD_RNO[7]\ : MX2
      port map(A => N_40, B => N_64, S => BIT_OS_SEL_4(0), Y => 
        \N_RECD_SER_WORD[7]\);
    
    \RECD_SER_WORD_RNO[1]\ : MX2
      port map(A => N_34, B => N_35, S => BIT_OS_SEL_4(0), Y => 
        \N_RECD_SER_WORD[1]\);
    
    \ARB_WRD_40M_FIXED[4]\ : DFN1C0
      port map(D => \Q[4]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[4]_net_1\);
    
    \RECD_SER_WORD_RNO[0]\ : MX2
      port map(A => N_33, B => N_34, S => BIT_OS_SEL_3_0, Y => 
        \N_RECD_SER_WORD[0]\);
    
    \Q[6]\ : DFN1C0
      port map(D => \ADJ_Q[6]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[6]_net_1\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \ARB_WRD_40M_FIXED[8]\ : DFN1C0
      port map(D => \Q[8]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[8]_net_1\);
    
    \ARB_BYTE[11]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[11]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[11]_net_1\);
    
    \Q[9]\ : DFN1C0
      port map(D => \ADJ_Q[9]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[9]_net_1\);
    
    \ARB_BYTE_RNINHR01[13]\ : MX2
      port map(A => N_24, B => N_32, S => BIT_OS_SEL_2(1), Y => 
        N_40);
    
    \Q[14]\ : DFN1C0
      port map(D => \ADJ_Q[14]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[14]_net_1\);
    
    ADJ_SER_IN_R_0DEL : DFN1C0
      port map(D => ELK_IN_R, CLK => CCC_160M_ADJ, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_R_0DEL\);
    
    \Q[13]\ : DFN1C0
      port map(D => \ADJ_Q[13]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[13]_net_1\);
    
    \ARB_BYTE[9]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[9]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[9]_net_1\);
    
    ADJ_SER_IN_R_1DEL : DFN1C0
      port map(D => \ADJ_SER_IN_R_0DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_R_1DEL\);
    
    \ARB_BYTE[10]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[10]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[10]_net_1\);
    
    \ADJ_Q[9]\ : DFN1C0
      port map(D => \ADJ_Q[7]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[9]_net_1\);
    
    \RECD_SER_WORD[7]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[7]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_14(7));
    
    \ARB_WRD_40M_FIXED[5]\ : DFN1C0
      port map(D => \Q[5]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[5]_net_1\);
    
    \ARB_WRD_40M_FIXED[12]\ : DFN1C0
      port map(D => \Q[12]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[12]_net_1\);
    
    \ARB_WRD_40M_FIXED[11]\ : DFN1C0
      port map(D => \Q[11]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[11]_net_1\);
    
    \ARB_BYTE_RNILK7G[12]\ : MX2
      port map(A => \ARB_BYTE[8]_net_1\, B => 
        \ARB_BYTE[12]_net_1\, S => BIT_OS_SEL_2(2), Y => N_31);
    
    \ARB_WRD_40M_FIXED[0]\ : DFN1C0
      port map(D => \Q[0]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[0]_net_1\);
    
    \ADJ_Q[10]\ : DFN1C0
      port map(D => \ADJ_Q[8]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[10]_net_1\);
    
    \Q[2]\ : DFN1C0
      port map(D => \ADJ_Q[2]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[2]_net_1\);
    
    \ARB_BYTE_RNIJI7G[11]\ : MX2
      port map(A => \ARB_BYTE[7]_net_1\, B => 
        \ARB_BYTE[11]_net_1\, S => BIT_OS_SEL_2(2), Y => N_24);
    
    \ARB_BYTE_RNI4J9C1[10]\ : MX2
      port map(A => N_21, B => N_23, S => BIT_OS_SEL_2(1), Y => 
        N_37);
    
    \ARB_BYTE_RNI2MLR[2]\ : MX2
      port map(A => \ARB_BYTE[2]_net_1\, B => \ARB_BYTE[6]_net_1\, 
        S => BIT_OS_SEL_2(2), Y => N_19);
    
    \ADJ_Q[1]\ : DFN1C0
      port map(D => \ADJ_SER_IN_F_1DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[1]_net_1\);
    
    \RECD_SER_WORD[6]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[6]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_14(6));
    
    \RECD_SER_WORD[2]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[2]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_14(2));
    
    \ADJ_Q[13]\ : DFN1C0
      port map(D => \ADJ_Q[11]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[13]_net_1\);
    
    \Q[8]\ : DFN1C0
      port map(D => \ADJ_Q[8]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[8]_net_1\);
    
    \ARB_BYTE[5]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[5]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[5]_net_1\);
    
    \ARB_BYTE_RNI8N9C1[11]\ : MX2
      port map(A => N_22, B => N_24, S => BIT_OS_SEL_2(1), Y => 
        N_38);
    
    \ADJ_Q[14]\ : DFN1C0
      port map(D => \ADJ_Q[12]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[14]_net_1\);
    
    \RECD_SER_WORD_RNO[4]\ : MX2
      port map(A => N_37, B => N_38, S => BIT_OS_SEL_4(0), Y => 
        \N_RECD_SER_WORD[4]\);
    
    \Q[12]\ : DFN1C0
      port map(D => \ADJ_Q[12]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[12]_net_1\);
    
    \ARB_BYTE[13]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[13]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[13]_net_1\);
    
    \ARB_WRD_40M_FIXED[3]\ : DFN1C0
      port map(D => \Q[3]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[3]_net_1\);
    
    \ARB_BYTE[7]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[7]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[7]_net_1\);
    
    \RECD_SER_WORD_RNO_0[0]\ : MX2
      port map(A => N_17, B => N_19, S => BIT_OS_SEL_2(1), Y => 
        N_33);
    
    \Q[4]\ : DFN1C0
      port map(D => \ADJ_Q[4]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[4]_net_1\);
    
    \ARB_WRD_40M_FIXED[7]\ : DFN1C0
      port map(D => \Q[7]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[7]_net_1\);
    
    \RECD_SER_WORD_RNO[6]\ : MX2
      port map(A => N_39, B => N_40, S => BIT_OS_SEL_4(0), Y => 
        \N_RECD_SER_WORD[6]\);
    
    \ARB_BYTE_RNIJDR01[10]\ : MX2
      port map(A => N_23, B => N_31, S => BIT_OS_SEL_2(1), Y => 
        N_39);
    
    \ARB_BYTE_RNIHKNN1[1]\ : MX2
      port map(A => N_18, B => N_20, S => BIT_OS_SEL_2(1), Y => 
        N_34);
    
    \ARB_BYTE_RNIPSNN1[3]\ : MX2
      port map(A => N_20, B => N_22, S => BIT_OS_SEL_2(1), Y => 
        N_36);
    
    \ARB_BYTE[3]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[3]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[3]_net_1\);
    
    \ADJ_Q[5]\ : DFN1C0
      port map(D => \ADJ_Q[3]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[5]_net_1\);
    
    \ARB_BYTE_RNI4OLR[3]\ : MX2
      port map(A => \ARB_BYTE[3]_net_1\, B => \ARB_BYTE[7]_net_1\, 
        S => BIT_OS_SEL_2(2), Y => N_20);
    
    \ARB_BYTE[1]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[1]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[1]_net_1\);
    
    \ARB_WRD_40M_FIXED[13]\ : DFN1C0
      port map(D => \Q[13]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[13]_net_1\);
    
    \ADJ_Q[0]\ : DFN1C0
      port map(D => \ADJ_SER_IN_R_1DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[0]_net_1\);
    
    \ARB_BYTE_RNI8SLR[5]\ : MX2
      port map(A => \ARB_BYTE[5]_net_1\, B => \ARB_BYTE[9]_net_1\, 
        S => BIT_OS_SEL_2(2), Y => N_22);
    
    \ARB_WRD_40M_FIXED[10]\ : DFN1C0
      port map(D => \Q[10]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[10]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SER320M_3_34_14 is

    port( ELK_TX_DAT                 : in    std_logic_vector(7 downto 0);
          MASTER_SALT_POR_B_i_0_i_2  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_5  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_10 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_0  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_12 : in    std_logic;
          ELK_OUT_R                  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_15 : in    std_logic;
          ELK_OUT_F                  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_7  : in    std_logic;
          CCC_160M_FXD               : in    std_logic;
          CLK_40M_GL                 : in    std_logic
        );

end SER320M_3_34_14;

architecture DEF_ARCH of SER320M_3_34_14 is 

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \N_SER_CMD_WORD_R[0]\, \START_RISE\, 
        \N_SER_CMD_WORD_F[0]\, \N_SER_CMD_WORD_R[3]\, 
        \SER_CMD_WORD_R[2]_net_1\, \N_SER_CMD_WORD_R[2]\, 
        \SER_CMD_WORD_R[1]_net_1\, \N_SER_CMD_WORD_R[1]\, 
        \SER_CMD_WORD_R[0]_net_1\, \N_SER_CMD_WORD_F[3]\, 
        \SER_CMD_WORD_F[2]_net_1\, \N_SER_CMD_WORD_F[2]\, 
        \SER_CMD_WORD_F[1]_net_1\, \N_SER_CMD_WORD_F[1]\, 
        \SER_CMD_WORD_F[0]_net_1\, N_START_RISE, 
        \CLK40M_GEN_DEL0\, \SER_OUT_FI\, \SER_OUT_RI\, 
        \SER_CMD_WORD_F[3]_net_1\, \SER_CMD_WORD_R[3]_net_1\, 
        \GND\, \VCC\ : std_logic;

begin 


    SER_OUT_FI : DFN1C0
      port map(D => \SER_CMD_WORD_F[3]_net_1\, CLK => 
        CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_10, Q => 
        \SER_OUT_FI\);
    
    \SER_CMD_WORD_F[3]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[3]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_5, Q => 
        \SER_CMD_WORD_F[3]_net_1\);
    
    \SER_CMD_WORD_R[1]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[1]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_2, Q => 
        \SER_CMD_WORD_R[1]_net_1\);
    
    \SER_CMD_WORD_R[2]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[2]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_2, Q => 
        \SER_CMD_WORD_R[2]_net_1\);
    
    \SER_CMD_WORD_R_RNO[3]\ : MX2
      port map(A => \SER_CMD_WORD_R[2]_net_1\, B => ELK_TX_DAT(7), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_R[3]\);
    
    \SER_CMD_WORD_R_RNO[0]\ : NOR2B
      port map(A => \START_RISE\, B => ELK_TX_DAT(1), Y => 
        \N_SER_CMD_WORD_R[0]\);
    
    \SER_CMD_WORD_F[0]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[0]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_5, Q => 
        \SER_CMD_WORD_F[0]_net_1\);
    
    \SER_CMD_WORD_R_RNO[1]\ : MX2
      port map(A => \SER_CMD_WORD_R[0]_net_1\, B => ELK_TX_DAT(3), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_R[1]\);
    
    \SER_CMD_WORD_F_RNO[2]\ : MX2
      port map(A => \SER_CMD_WORD_F[1]_net_1\, B => ELK_TX_DAT(4), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_F[2]\);
    
    \SER_CMD_WORD_F_RNO[3]\ : MX2
      port map(A => \SER_CMD_WORD_F[2]_net_1\, B => ELK_TX_DAT(6), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_F[3]\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    CLK40M_GEN_DEL0 : DFN1C0
      port map(D => CLK_40M_GL, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_7, Q => \CLK40M_GEN_DEL0\);
    
    SER_OUT_RI : DFN1C0
      port map(D => \SER_CMD_WORD_R[3]_net_1\, CLK => 
        CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_10, Q => 
        \SER_OUT_RI\);
    
    \SER_CMD_WORD_F[2]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[2]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_5, Q => 
        \SER_CMD_WORD_F[2]_net_1\);
    
    \SER_CMD_WORD_F_RNO[1]\ : MX2
      port map(A => \SER_CMD_WORD_F[0]_net_1\, B => ELK_TX_DAT(2), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_F[1]\);
    
    \SER_CMD_WORD_R[0]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[0]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_2, Q => 
        \SER_CMD_WORD_R[0]_net_1\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    START_RISE : DFN1C0
      port map(D => N_START_RISE, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_0, Q => \START_RISE\);
    
    \SER_CMD_WORD_R[3]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[3]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_2, Q => 
        \SER_CMD_WORD_R[3]_net_1\);
    
    \SER_CMD_WORD_F_RNO[0]\ : NOR2B
      port map(A => \START_RISE\, B => ELK_TX_DAT(0), Y => 
        \N_SER_CMD_WORD_F[0]\);
    
    SER_OUT_RDEL : DFN1C0
      port map(D => \SER_OUT_RI\, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_12, Q => ELK_OUT_R);
    
    \SER_CMD_WORD_F[1]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[1]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_5, Q => 
        \SER_CMD_WORD_F[1]_net_1\);
    
    START_RISE_RNO : NOR2B
      port map(A => \CLK40M_GEN_DEL0\, B => CLK_40M_GL, Y => 
        N_START_RISE);
    
    \SER_CMD_WORD_R_RNO[2]\ : MX2
      port map(A => \SER_CMD_WORD_R[1]_net_1\, B => ELK_TX_DAT(5), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_R[2]\);
    
    SER_OUT_FDEL : DFN1C0
      port map(D => \SER_OUT_FI\, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_15, Q => ELK_OUT_F);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity DDR_BIDIR_LVDS_DUAL_CLK_14 is

    port( DCB_SALT_SEL_c_i : in    std_logic;
          ELK14_DAT_P      : inout std_logic := 'Z';
          ELK14_DAT_N      : inout std_logic := 'Z';
          ELK_OUT_R        : in    std_logic;
          ELK_OUT_F        : in    std_logic;
          CCC_160M_FXD     : in    std_logic;
          CCC_160M_ADJ     : in    std_logic;
          ELK_IN_DDR_R     : out   std_logic;
          ELK_IN_DDR_F     : out   std_logic
        );

end DDR_BIDIR_LVDS_DUAL_CLK_14;

architecture DEF_ARCH of DDR_BIDIR_LVDS_DUAL_CLK_14 is 

  component DDR_REG
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          QR  : out   std_logic;
          QF  : out   std_logic
        );
  end component;

  component DDR_OUT
    port( DR  : in    std_logic := 'U';
          DF  : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component BIBUF_LVDS
    port( PADP : inout   std_logic;
          PADN : inout   std_logic;
          D    : in    std_logic := 'U';
          E    : in    std_logic := 'U';
          Y    : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal DDR_BIDIR_LVDS_DUAL_CLK_14_GND, BIBUF_LVDS_0_Y, 
        DDR_OUT_0_Q, \VCC\ : std_logic;

begin 


    DDR_REG_0 : DDR_REG
      port map(D => BIBUF_LVDS_0_Y, CLK => CCC_160M_ADJ, CLR => 
        DDR_BIDIR_LVDS_DUAL_CLK_14_GND, QR => ELK_IN_DDR_R, QF
         => ELK_IN_DDR_F);
    
    DDR_OUT_0 : DDR_OUT
      port map(DR => ELK_OUT_R, DF => ELK_OUT_F, CLK => 
        CCC_160M_FXD, CLR => DDR_BIDIR_LVDS_DUAL_CLK_14_GND, Q
         => DDR_OUT_0_Q);
    
    BIBUF_LVDS_0 : BIBUF_LVDS
      port map(PADP => ELK14_DAT_P, PADN => ELK14_DAT_N, D => 
        DDR_OUT_0_Q, E => DCB_SALT_SEL_c_i, Y => BIBUF_LVDS_0_Y);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    GND_i : GND
      port map(Y => DDR_BIDIR_LVDS_DUAL_CLK_14_GND);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SYNC_DAT_SEL_14 is

    port( ELK_TX_DAT                : out   std_logic_vector(7 downto 0);
          PATT_ELK_DAT_14           : in    std_logic_vector(7 downto 0);
          OP_MODE_c_2_0             : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_6 : in    std_logic;
          CLK_40M_GL                : in    std_logic
        );

end SYNC_DAT_SEL_14;

architecture DEF_ARCH of SYNC_DAT_SEL_14 is 

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \N_SERDAT[0]\, \N_SERDAT[1]\, \N_SERDAT[2]\, 
        \N_SERDAT[3]\, \N_SERDAT[4]\, \N_SERDAT[7]\, 
        \N_SERDAT[6]\, \N_SERDAT[5]\, \GND\, \VCC\ : std_logic;

begin 


    \SERDAT_RNO[4]\ : NOR2A
      port map(A => PATT_ELK_DAT_14(4), B => OP_MODE_c_2_0, Y => 
        \N_SERDAT[4]\);
    
    \SERDAT_RNO[0]\ : NOR2A
      port map(A => PATT_ELK_DAT_14(0), B => OP_MODE_c_2_0, Y => 
        \N_SERDAT[0]\);
    
    \SERDAT[6]\ : DFN1C0
      port map(D => \N_SERDAT[6]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_6, Q => ELK_TX_DAT(6));
    
    \SERDAT[4]\ : DFN1C0
      port map(D => \N_SERDAT[4]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_6, Q => ELK_TX_DAT(4));
    
    \SERDAT_RNO[7]\ : OR2
      port map(A => PATT_ELK_DAT_14(7), B => OP_MODE_c_2_0, Y => 
        \N_SERDAT[7]\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \SERDAT_RNO[3]\ : OR2
      port map(A => PATT_ELK_DAT_14(3), B => OP_MODE_c_2_0, Y => 
        \N_SERDAT[3]\);
    
    \SERDAT_RNO[2]\ : OR2
      port map(A => PATT_ELK_DAT_14(2), B => OP_MODE_c_2_0, Y => 
        \N_SERDAT[2]\);
    
    \SERDAT[5]\ : DFN1C0
      port map(D => \N_SERDAT[5]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_6, Q => ELK_TX_DAT(5));
    
    \SERDAT[7]\ : DFN1C0
      port map(D => \N_SERDAT[7]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_6, Q => ELK_TX_DAT(7));
    
    GND_i : GND
      port map(Y => \GND\);
    
    \SERDAT_RNO[5]\ : NOR2A
      port map(A => PATT_ELK_DAT_14(5), B => OP_MODE_c_2_0, Y => 
        \N_SERDAT[5]\);
    
    \SERDAT[0]\ : DFN1C0
      port map(D => \N_SERDAT[0]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_6, Q => ELK_TX_DAT(0));
    
    \SERDAT_RNO[6]\ : NOR2A
      port map(A => PATT_ELK_DAT_14(6), B => OP_MODE_c_2_0, Y => 
        \N_SERDAT[6]\);
    
    \SERDAT[1]\ : DFN1C0
      port map(D => \N_SERDAT[1]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_6, Q => ELK_TX_DAT(1));
    
    \SERDAT_RNO[1]\ : OR2
      port map(A => PATT_ELK_DAT_14(1), B => OP_MODE_c_2_0, Y => 
        \N_SERDAT[1]\);
    
    \SERDAT[3]\ : DFN1C0
      port map(D => \N_SERDAT[3]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_6, Q => ELK_TX_DAT(3));
    
    \SERDAT[2]\ : DFN1C0
      port map(D => \N_SERDAT[2]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_6, Q => ELK_TX_DAT(2));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity ELINK_SLAVE_15_9 is

    port( BIT_OS_SEL_2               : in    std_logic_vector(2 downto 1);
          BIT_OS_SEL_5_0             : in    std_logic;
          BIT_OS_SEL_3_0             : in    std_logic;
          BIT_OS_SEL_4               : in    std_logic_vector(1 downto 0);
          ELK_RX_SER_WORD_14         : out   std_logic_vector(7 downto 0);
          OP_MODE_c_2_0              : in    std_logic;
          PATT_ELK_DAT_14            : in    std_logic_vector(7 downto 0);
          MASTER_DCB_POR_B_i_0_i     : in    std_logic;
          ELK14_DAT_N                : inout std_logic := 'Z';
          ELK14_DAT_P                : inout std_logic := 'Z';
          DCB_SALT_SEL_c_i           : in    std_logic;
          CCC_160M_FXD               : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_7  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_15 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_12 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_0  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_10 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_5  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_2  : in    std_logic;
          CLK_40M_GL                 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_6  : in    std_logic;
          DEV_RST_B_c                : in    std_logic;
          CCC_160M_ADJ               : in    std_logic
        );

end ELINK_SLAVE_15_9;

architecture DEF_ARCH of ELINK_SLAVE_15_9 is 

  component SLAVE_DES320S_1_17_12
    port( ELK_RX_SER_WORD_14     : out   std_logic_vector(7 downto 0);
          BIT_OS_SEL_4           : in    std_logic_vector(1 downto 0) := (others => 'U');
          BIT_OS_SEL_3_0         : in    std_logic := 'U';
          BIT_OS_SEL_5_0         : in    std_logic := 'U';
          BIT_OS_SEL_2           : in    std_logic_vector(2 downto 1) := (others => 'U');
          CLK_40M_GL             : in    std_logic := 'U';
          CCC_160M_FXD           : in    std_logic := 'U';
          ELK_IN_R               : in    std_logic := 'U';
          ELK_IN_F               : in    std_logic := 'U';
          MASTER_DCB_POR_B_i_0_i : in    std_logic := 'U';
          CCC_160M_ADJ           : in    std_logic := 'U'
        );
  end component;

  component SER320M_3_34_14
    port( ELK_TX_DAT                 : in    std_logic_vector(7 downto 0) := (others => 'U');
          MASTER_SALT_POR_B_i_0_i_2  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_5  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_10 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_0  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_12 : in    std_logic := 'U';
          ELK_OUT_R                  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_15 : in    std_logic := 'U';
          ELK_OUT_F                  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_7  : in    std_logic := 'U';
          CCC_160M_FXD               : in    std_logic := 'U';
          CLK_40M_GL                 : in    std_logic := 'U'
        );
  end component;

  component DDR_BIDIR_LVDS_DUAL_CLK_14
    port( DCB_SALT_SEL_c_i : in    std_logic := 'U';
          ELK14_DAT_P      : inout   std_logic;
          ELK14_DAT_N      : inout   std_logic;
          ELK_OUT_R        : in    std_logic := 'U';
          ELK_OUT_F        : in    std_logic := 'U';
          CCC_160M_FXD     : in    std_logic := 'U';
          CCC_160M_ADJ     : in    std_logic := 'U';
          ELK_IN_DDR_R     : out   std_logic;
          ELK_IN_DDR_F     : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component SYNC_DAT_SEL_14
    port( ELK_TX_DAT                : out   std_logic_vector(7 downto 0);
          PATT_ELK_DAT_14           : in    std_logic_vector(7 downto 0) := (others => 'U');
          OP_MODE_c_2_0             : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_6 : in    std_logic := 'U';
          CLK_40M_GL                : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \ELK_IN_F\, ELK_IN_DDR_F, \ELK_IN_R\, ELK_IN_DDR_R, 
        \ELK_TX_DAT[0]\, \ELK_TX_DAT[1]\, \ELK_TX_DAT[2]\, 
        \ELK_TX_DAT[3]\, \ELK_TX_DAT[4]\, \ELK_TX_DAT[5]\, 
        \ELK_TX_DAT[6]\, \ELK_TX_DAT[7]\, ELK_OUT_R, ELK_OUT_F, 
        \GND\, \VCC\ : std_logic;

    for all : SLAVE_DES320S_1_17_12
	Use entity work.SLAVE_DES320S_1_17_12(DEF_ARCH);
    for all : SER320M_3_34_14
	Use entity work.SER320M_3_34_14(DEF_ARCH);
    for all : DDR_BIDIR_LVDS_DUAL_CLK_14
	Use entity work.DDR_BIDIR_LVDS_DUAL_CLK_14(DEF_ARCH);
    for all : SYNC_DAT_SEL_14
	Use entity work.SYNC_DAT_SEL_14(DEF_ARCH);
begin 


    U_SLAVE_1ELK : SLAVE_DES320S_1_17_12
      port map(ELK_RX_SER_WORD_14(7) => ELK_RX_SER_WORD_14(7), 
        ELK_RX_SER_WORD_14(6) => ELK_RX_SER_WORD_14(6), 
        ELK_RX_SER_WORD_14(5) => ELK_RX_SER_WORD_14(5), 
        ELK_RX_SER_WORD_14(4) => ELK_RX_SER_WORD_14(4), 
        ELK_RX_SER_WORD_14(3) => ELK_RX_SER_WORD_14(3), 
        ELK_RX_SER_WORD_14(2) => ELK_RX_SER_WORD_14(2), 
        ELK_RX_SER_WORD_14(1) => ELK_RX_SER_WORD_14(1), 
        ELK_RX_SER_WORD_14(0) => ELK_RX_SER_WORD_14(0), 
        BIT_OS_SEL_4(1) => BIT_OS_SEL_4(1), BIT_OS_SEL_4(0) => 
        BIT_OS_SEL_4(0), BIT_OS_SEL_3_0 => BIT_OS_SEL_3_0, 
        BIT_OS_SEL_5_0 => BIT_OS_SEL_5_0, BIT_OS_SEL_2(2) => 
        BIT_OS_SEL_2(2), BIT_OS_SEL_2(1) => BIT_OS_SEL_2(1), 
        CLK_40M_GL => CLK_40M_GL, CCC_160M_FXD => CCC_160M_FXD, 
        ELK_IN_R => \ELK_IN_R\, ELK_IN_F => \ELK_IN_F\, 
        MASTER_DCB_POR_B_i_0_i => MASTER_DCB_POR_B_i_0_i, 
        CCC_160M_ADJ => CCC_160M_ADJ);
    
    U_ELK1_CMD_TX : SER320M_3_34_14
      port map(ELK_TX_DAT(7) => \ELK_TX_DAT[7]\, ELK_TX_DAT(6)
         => \ELK_TX_DAT[6]\, ELK_TX_DAT(5) => \ELK_TX_DAT[5]\, 
        ELK_TX_DAT(4) => \ELK_TX_DAT[4]\, ELK_TX_DAT(3) => 
        \ELK_TX_DAT[3]\, ELK_TX_DAT(2) => \ELK_TX_DAT[2]\, 
        ELK_TX_DAT(1) => \ELK_TX_DAT[1]\, ELK_TX_DAT(0) => 
        \ELK_TX_DAT[0]\, MASTER_SALT_POR_B_i_0_i_2 => 
        MASTER_SALT_POR_B_i_0_i_2, MASTER_SALT_POR_B_i_0_i_5 => 
        MASTER_SALT_POR_B_i_0_i_5, MASTER_SALT_POR_B_i_0_i_10 => 
        MASTER_SALT_POR_B_i_0_i_10, MASTER_SALT_POR_B_i_0_i_0 => 
        MASTER_SALT_POR_B_i_0_i_0, MASTER_SALT_POR_B_i_0_i_12 => 
        MASTER_SALT_POR_B_i_0_i_12, ELK_OUT_R => ELK_OUT_R, 
        MASTER_SALT_POR_B_i_0_i_15 => MASTER_SALT_POR_B_i_0_i_15, 
        ELK_OUT_F => ELK_OUT_F, MASTER_SALT_POR_B_i_0_i_7 => 
        MASTER_SALT_POR_B_i_0_i_7, CCC_160M_FXD => CCC_160M_FXD, 
        CLK_40M_GL => CLK_40M_GL);
    
    U_DDR_ELK1 : DDR_BIDIR_LVDS_DUAL_CLK_14
      port map(DCB_SALT_SEL_c_i => DCB_SALT_SEL_c_i, ELK14_DAT_P
         => ELK14_DAT_P, ELK14_DAT_N => ELK14_DAT_N, ELK_OUT_R
         => ELK_OUT_R, ELK_OUT_F => ELK_OUT_F, CCC_160M_FXD => 
        CCC_160M_FXD, CCC_160M_ADJ => CCC_160M_ADJ, ELK_IN_DDR_R
         => ELK_IN_DDR_R, ELK_IN_DDR_F => ELK_IN_DDR_F);
    
    ELK_IN_F : DFN1C0
      port map(D => ELK_IN_DDR_F, CLK => CCC_160M_ADJ, CLR => 
        DEV_RST_B_c, Q => \ELK_IN_F\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    U_ELK1_SERDAT_SOURCE : SYNC_DAT_SEL_14
      port map(ELK_TX_DAT(7) => \ELK_TX_DAT[7]\, ELK_TX_DAT(6)
         => \ELK_TX_DAT[6]\, ELK_TX_DAT(5) => \ELK_TX_DAT[5]\, 
        ELK_TX_DAT(4) => \ELK_TX_DAT[4]\, ELK_TX_DAT(3) => 
        \ELK_TX_DAT[3]\, ELK_TX_DAT(2) => \ELK_TX_DAT[2]\, 
        ELK_TX_DAT(1) => \ELK_TX_DAT[1]\, ELK_TX_DAT(0) => 
        \ELK_TX_DAT[0]\, PATT_ELK_DAT_14(7) => PATT_ELK_DAT_14(7), 
        PATT_ELK_DAT_14(6) => PATT_ELK_DAT_14(6), 
        PATT_ELK_DAT_14(5) => PATT_ELK_DAT_14(5), 
        PATT_ELK_DAT_14(4) => PATT_ELK_DAT_14(4), 
        PATT_ELK_DAT_14(3) => PATT_ELK_DAT_14(3), 
        PATT_ELK_DAT_14(2) => PATT_ELK_DAT_14(2), 
        PATT_ELK_DAT_14(1) => PATT_ELK_DAT_14(1), 
        PATT_ELK_DAT_14(0) => PATT_ELK_DAT_14(0), OP_MODE_c_2_0
         => OP_MODE_c_2_0, MASTER_SALT_POR_B_i_0_i_6 => 
        MASTER_SALT_POR_B_i_0_i_6, CLK_40M_GL => CLK_40M_GL);
    
    ELK_IN_R : DFN1C0
      port map(D => ELK_IN_DDR_R, CLK => CCC_160M_ADJ, CLR => 
        DEV_RST_B_c, Q => \ELK_IN_R\);
    
    GND_i : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity tristate_buf_0 is

    port( P_USB_MASTER_EN_c : in    std_logic;
          USB_WR_BI         : in    std_logic;
          USB_WR_B          : out   std_logic
        );

end tristate_buf_0;

architecture DEF_ARCH of tristate_buf_0 is 

  component TRIBUFF_F_24U
    port( D   : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          PAD : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \GND\, \VCC\ : std_logic;

begin 


    \TRIBUFF_F_24U[0]\ : TRIBUFF_F_24U
      port map(D => USB_WR_BI, E => P_USB_MASTER_EN_c, PAD => 
        USB_WR_B);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    GND_i : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SLAVE_DES320S_1_17_0 is

    port( ELK_RX_SER_WORD_2      : out   std_logic_vector(7 downto 0);
          BIT_OS_SEL_1           : in    std_logic_vector(1 downto 0);
          BIT_OS_SEL_0_0         : in    std_logic;
          BIT_OS_SEL             : in    std_logic_vector(2 downto 1);
          BIT_OS_SEL_7_0         : in    std_logic;
          CLK_40M_GL             : in    std_logic;
          CCC_160M_FXD           : in    std_logic;
          ELK_IN_R               : in    std_logic;
          ELK_IN_F               : in    std_logic;
          MASTER_DCB_POR_B_i_0_i : in    std_logic;
          CCC_160M_ADJ           : in    std_logic
        );

end SLAVE_DES320S_1_17_0;

architecture DEF_ARCH of SLAVE_DES320S_1_17_0 is 

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal N_17, \ARB_BYTE[0]_net_1\, \ARB_BYTE[4]_net_1\, N_18, 
        \ARB_BYTE[1]_net_1\, \ARB_BYTE[5]_net_1\, N_19, 
        \ARB_BYTE[2]_net_1\, \ARB_BYTE[6]_net_1\, N_20, 
        \ARB_BYTE[3]_net_1\, \ARB_BYTE[7]_net_1\, N_21, 
        \ARB_BYTE[8]_net_1\, N_22, \ARB_BYTE[9]_net_1\, N_23, 
        \ARB_BYTE[10]_net_1\, N_24, \ARB_BYTE[11]_net_1\, N_31, 
        \ARB_BYTE[12]_net_1\, N_32, \ARB_BYTE[13]_net_1\, N_33, 
        N_34, N_35, N_36, N_37, N_38, N_39, N_40, N_56, 
        \ARB_BYTE[14]_net_1\, N_64, \N_RECD_SER_WORD[0]\, 
        \N_RECD_SER_WORD[1]\, \N_RECD_SER_WORD[2]\, 
        \N_RECD_SER_WORD[3]\, \N_RECD_SER_WORD[4]\, 
        \N_RECD_SER_WORD[5]\, \N_RECD_SER_WORD[6]\, 
        \N_RECD_SER_WORD[7]\, \ADJ_SER_IN_F_0DEL\, 
        \ADJ_SER_IN_R_0DEL\, \ADJ_SER_IN_F_1DEL\, 
        \ADJ_SER_IN_R_1DEL\, \Q[0]_net_1\, \ADJ_Q[0]_net_1\, 
        \Q[1]_net_1\, \ADJ_Q[1]_net_1\, \Q[2]_net_1\, 
        \ADJ_Q[2]_net_1\, \Q[3]_net_1\, \ADJ_Q[3]_net_1\, 
        \Q[4]_net_1\, \ADJ_Q[4]_net_1\, \Q[5]_net_1\, 
        \ADJ_Q[5]_net_1\, \Q[6]_net_1\, \ADJ_Q[6]_net_1\, 
        \Q[7]_net_1\, \ADJ_Q[7]_net_1\, \Q[8]_net_1\, 
        \ADJ_Q[8]_net_1\, \Q[9]_net_1\, \ADJ_Q[9]_net_1\, 
        \Q[10]_net_1\, \ADJ_Q[10]_net_1\, \Q[11]_net_1\, 
        \ADJ_Q[11]_net_1\, \Q[12]_net_1\, \ADJ_Q[12]_net_1\, 
        \Q[13]_net_1\, \ADJ_Q[13]_net_1\, \Q[14]_net_1\, 
        \ADJ_Q[14]_net_1\, \ARB_WRD_40M_FIXED[0]_net_1\, 
        \ARB_WRD_40M_FIXED[1]_net_1\, 
        \ARB_WRD_40M_FIXED[2]_net_1\, 
        \ARB_WRD_40M_FIXED[3]_net_1\, 
        \ARB_WRD_40M_FIXED[4]_net_1\, 
        \ARB_WRD_40M_FIXED[5]_net_1\, 
        \ARB_WRD_40M_FIXED[6]_net_1\, 
        \ARB_WRD_40M_FIXED[7]_net_1\, 
        \ARB_WRD_40M_FIXED[8]_net_1\, 
        \ARB_WRD_40M_FIXED[9]_net_1\, 
        \ARB_WRD_40M_FIXED[10]_net_1\, 
        \ARB_WRD_40M_FIXED[11]_net_1\, 
        \ARB_WRD_40M_FIXED[12]_net_1\, 
        \ARB_WRD_40M_FIXED[13]_net_1\, 
        \ARB_WRD_40M_FIXED[14]_net_1\, \GND\, \VCC\ : std_logic;

begin 


    \RECD_SER_WORD_RNO[5]\ : MX2
      port map(A => N_38, B => N_39, S => BIT_OS_SEL_1(0), Y => 
        \N_RECD_SER_WORD[5]\);
    
    \ARB_WRD_40M_FIXED[9]\ : DFN1C0
      port map(D => \Q[9]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[9]_net_1\);
    
    \ADJ_Q[4]\ : DFN1C0
      port map(D => \ADJ_Q[2]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[4]_net_1\);
    
    \ARB_BYTE[6]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[6]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[6]_net_1\);
    
    ADJ_SER_IN_F_1DEL : DFN1C0
      port map(D => \ADJ_SER_IN_F_0DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_F_1DEL\);
    
    \ARB_BYTE[0]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[0]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[0]_net_1\);
    
    \Q[11]\ : DFN1C0
      port map(D => \ADJ_Q[11]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[11]_net_1\);
    
    \ARB_BYTE_RNIH7KF1[10]\ : MX2
      port map(A => N_21, B => N_23, S => BIT_OS_SEL(1), Y => 
        N_37);
    
    \ADJ_Q[8]\ : DFN1C0
      port map(D => \ADJ_Q[6]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[8]_net_1\);
    
    \ADJ_Q[6]\ : DFN1C0
      port map(D => \ADJ_Q[4]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[6]_net_1\);
    
    \ADJ_Q[12]\ : DFN1C0
      port map(D => \ADJ_Q[10]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[12]_net_1\);
    
    \RECD_SER_WORD_RNO_1[0]\ : MX2
      port map(A => \ARB_BYTE[0]_net_1\, B => \ARB_BYTE[4]_net_1\, 
        S => BIT_OS_SEL_7_0, Y => N_17);
    
    \Q[1]\ : DFN1C0
      port map(D => \ADJ_Q[1]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[1]_net_1\);
    
    \ARB_BYTE[4]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[4]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[4]_net_1\);
    
    \ADJ_Q[2]\ : DFN1C0
      port map(D => \ADJ_Q[0]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[2]_net_1\);
    
    \RECD_SER_WORD_RNO_1[7]\ : MX2
      port map(A => \ARB_BYTE[10]_net_1\, B => 
        \ARB_BYTE[14]_net_1\, S => BIT_OS_SEL_0_0, Y => N_56);
    
    \RECD_SER_WORD[4]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[4]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_2(4));
    
    \Q[5]\ : DFN1C0
      port map(D => \ADJ_Q[5]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[5]_net_1\);
    
    \ADJ_Q[11]\ : DFN1C0
      port map(D => \ADJ_Q[9]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[11]_net_1\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \ADJ_Q[3]\ : DFN1C0
      port map(D => \ADJ_Q[1]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[3]_net_1\);
    
    \Q[10]\ : DFN1C0
      port map(D => \ADJ_Q[10]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[10]_net_1\);
    
    \ARB_WRD_40M_FIXED[6]\ : DFN1C0
      port map(D => \Q[6]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[6]_net_1\);
    
    \ARB_WRD_40M_FIXED[1]\ : DFN1C0
      port map(D => \Q[1]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[1]_net_1\);
    
    \RECD_SER_WORD[3]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[3]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_2(3));
    
    \RECD_SER_WORD[0]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[0]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_2(0));
    
    \RECD_SER_WORD_RNO[3]\ : MX2
      port map(A => N_36, B => N_37, S => BIT_OS_SEL_1(0), Y => 
        \N_RECD_SER_WORD[3]\);
    
    \Q[0]\ : DFN1C0
      port map(D => \ADJ_Q[0]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[0]_net_1\);
    
    \ARB_BYTE_RNIUROM1[1]\ : MX2
      port map(A => N_18, B => N_20, S => BIT_OS_SEL(1), Y => 
        N_34);
    
    \RECD_SER_WORD_RNO_0[7]\ : MX2
      port map(A => N_31, B => N_56, S => BIT_OS_SEL_1(1), Y => 
        N_64);
    
    \Q[7]\ : DFN1C0
      port map(D => \ADJ_Q[7]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[7]_net_1\);
    
    \ARB_BYTE[14]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[14]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[14]_net_1\);
    
    \ARB_WRD_40M_FIXED[2]\ : DFN1C0
      port map(D => \Q[2]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[2]_net_1\);
    
    \ARB_WRD_40M_FIXED[14]\ : DFN1C0
      port map(D => \Q[14]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[14]_net_1\);
    
    \RECD_SER_WORD_RNO[2]\ : MX2
      port map(A => N_35, B => N_36, S => BIT_OS_SEL_1(0), Y => 
        \N_RECD_SER_WORD[2]\);
    
    \ARB_BYTE[2]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[2]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[2]_net_1\);
    
    \ADJ_Q[7]\ : DFN1C0
      port map(D => \ADJ_Q[5]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[7]_net_1\);
    
    \ARB_BYTE[8]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[8]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[8]_net_1\);
    
    \RECD_SER_WORD[5]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[5]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_2(5));
    
    \ARB_BYTE[12]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[12]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[12]_net_1\);
    
    \ARB_BYTE_RNI7UDN[5]\ : MX2
      port map(A => \ARB_BYTE[5]_net_1\, B => \ARB_BYTE[9]_net_1\, 
        S => BIT_OS_SEL_7_0, Y => N_22);
    
    \RECD_SER_WORD[1]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[1]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_2(1));
    
    \ARB_BYTE_RNI64PM1[3]\ : MX2
      port map(A => N_20, B => N_22, S => BIT_OS_SEL(1), Y => 
        N_36);
    
    \ARB_BYTE_RNI5SDN[4]\ : MX2
      port map(A => \ARB_BYTE[4]_net_1\, B => \ARB_BYTE[8]_net_1\, 
        S => BIT_OS_SEL_7_0, Y => N_21);
    
    \Q[3]\ : DFN1C0
      port map(D => \ADJ_Q[3]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[3]_net_1\);
    
    ADJ_SER_IN_F_0DEL : DFN1C0
      port map(D => ELK_IN_F, CLK => CCC_160M_ADJ, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_F_0DEL\);
    
    \RECD_SER_WORD_RNO[7]\ : MX2
      port map(A => N_40, B => N_64, S => BIT_OS_SEL_1(0), Y => 
        \N_RECD_SER_WORD[7]\);
    
    \RECD_SER_WORD_RNO[1]\ : MX2
      port map(A => N_34, B => N_35, S => BIT_OS_SEL_1(0), Y => 
        \N_RECD_SER_WORD[1]\);
    
    \ARB_WRD_40M_FIXED[4]\ : DFN1C0
      port map(D => \Q[4]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[4]_net_1\);
    
    \ARB_BYTE_RNILBKF1[11]\ : MX2
      port map(A => N_22, B => N_24, S => BIT_OS_SEL(1), Y => 
        N_38);
    
    \RECD_SER_WORD_RNO[0]\ : MX2
      port map(A => N_33, B => N_34, S => BIT_OS_SEL_1(0), Y => 
        \N_RECD_SER_WORD[0]\);
    
    \Q[6]\ : DFN1C0
      port map(D => \ADJ_Q[6]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[6]_net_1\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \ARB_WRD_40M_FIXED[8]\ : DFN1C0
      port map(D => \Q[8]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[8]_net_1\);
    
    \ARB_BYTE_RNIGV8G[10]\ : MX2
      port map(A => \ARB_BYTE[6]_net_1\, B => 
        \ARB_BYTE[10]_net_1\, S => BIT_OS_SEL_7_0, Y => N_23);
    
    \ARB_BYTE[11]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[11]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[11]_net_1\);
    
    \Q[9]\ : DFN1C0
      port map(D => \ADJ_Q[9]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[9]_net_1\);
    
    \ARB_BYTE_RNIE7HA1[13]\ : MX2
      port map(A => N_24, B => N_32, S => BIT_OS_SEL(1), Y => 
        N_40);
    
    \Q[14]\ : DFN1C0
      port map(D => \ADJ_Q[14]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[14]_net_1\);
    
    ADJ_SER_IN_R_0DEL : DFN1C0
      port map(D => ELK_IN_R, CLK => CCC_160M_ADJ, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_R_0DEL\);
    
    \Q[13]\ : DFN1C0
      port map(D => \ADJ_Q[13]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[13]_net_1\);
    
    \ARB_BYTE[9]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[9]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[9]_net_1\);
    
    ADJ_SER_IN_R_1DEL : DFN1C0
      port map(D => \ADJ_SER_IN_R_0DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_R_1DEL\);
    
    \ARB_BYTE[10]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[10]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[10]_net_1\);
    
    \ADJ_Q[9]\ : DFN1C0
      port map(D => \ADJ_Q[7]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[9]_net_1\);
    
    \RECD_SER_WORD[7]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[7]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_2(7));
    
    \ARB_WRD_40M_FIXED[5]\ : DFN1C0
      port map(D => \Q[5]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[5]_net_1\);
    
    \ARB_WRD_40M_FIXED[12]\ : DFN1C0
      port map(D => \Q[12]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[12]_net_1\);
    
    \ARB_WRD_40M_FIXED[11]\ : DFN1C0
      port map(D => \Q[11]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[11]_net_1\);
    
    \ARB_BYTE_RNI0FF81[10]\ : MX2
      port map(A => N_23, B => N_31, S => BIT_OS_SEL(1), Y => 
        N_39);
    
    \ARB_WRD_40M_FIXED[0]\ : DFN1C0
      port map(D => \Q[0]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[0]_net_1\);
    
    \ADJ_Q[10]\ : DFN1C0
      port map(D => \ADJ_Q[8]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[10]_net_1\);
    
    \Q[2]\ : DFN1C0
      port map(D => \ADJ_Q[2]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[2]_net_1\);
    
    \ARB_BYTE_RNIVLDN[1]\ : MX2
      port map(A => \ARB_BYTE[1]_net_1\, B => \ARB_BYTE[5]_net_1\, 
        S => BIT_OS_SEL_7_0, Y => N_18);
    
    \ADJ_Q[1]\ : DFN1C0
      port map(D => \ADJ_SER_IN_F_1DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[1]_net_1\);
    
    \RECD_SER_WORD[6]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[6]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_2(6));
    
    \RECD_SER_WORD[2]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[2]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_2(2));
    
    \ADJ_Q[13]\ : DFN1C0
      port map(D => \ADJ_Q[11]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[13]_net_1\);
    
    \Q[8]\ : DFN1C0
      port map(D => \ADJ_Q[8]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[8]_net_1\);
    
    \ARB_BYTE_RNI3QDN[3]\ : MX2
      port map(A => \ARB_BYTE[3]_net_1\, B => \ARB_BYTE[7]_net_1\, 
        S => BIT_OS_SEL_7_0, Y => N_20);
    
    \ARB_BYTE[5]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[5]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[5]_net_1\);
    
    \ADJ_Q[14]\ : DFN1C0
      port map(D => \ADJ_Q[12]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[14]_net_1\);
    
    \RECD_SER_WORD_RNO[4]\ : MX2
      port map(A => N_37, B => N_38, S => BIT_OS_SEL_1(0), Y => 
        \N_RECD_SER_WORD[4]\);
    
    \Q[12]\ : DFN1C0
      port map(D => \ADJ_Q[12]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[12]_net_1\);
    
    \ARB_BYTE[13]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[13]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[13]_net_1\);
    
    \ARB_WRD_40M_FIXED[3]\ : DFN1C0
      port map(D => \Q[3]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[3]_net_1\);
    
    \ARB_BYTE[7]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[7]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[7]_net_1\);
    
    \RECD_SER_WORD_RNO_0[0]\ : MX2
      port map(A => N_17, B => N_19, S => BIT_OS_SEL(1), Y => 
        N_33);
    
    \Q[4]\ : DFN1C0
      port map(D => \ADJ_Q[4]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[4]_net_1\);
    
    \ARB_WRD_40M_FIXED[7]\ : DFN1C0
      port map(D => \Q[7]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[7]_net_1\);
    
    \ARB_BYTE_RNII19G[11]\ : MX2
      port map(A => \ARB_BYTE[7]_net_1\, B => 
        \ARB_BYTE[11]_net_1\, S => BIT_OS_SEL_7_0, Y => N_24);
    
    \ARB_BYTE_RNIK39G[12]\ : MX2
      port map(A => \ARB_BYTE[8]_net_1\, B => 
        \ARB_BYTE[12]_net_1\, S => BIT_OS_SEL_7_0, Y => N_31);
    
    \RECD_SER_WORD_RNO[6]\ : MX2
      port map(A => N_39, B => N_40, S => BIT_OS_SEL_1(0), Y => 
        \N_RECD_SER_WORD[6]\);
    
    \ARB_BYTE_RNI1ODN[2]\ : MX2
      port map(A => \ARB_BYTE[2]_net_1\, B => \ARB_BYTE[6]_net_1\, 
        S => BIT_OS_SEL_7_0, Y => N_19);
    
    \ARB_BYTE[3]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[3]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[3]_net_1\);
    
    \ARB_BYTE_RNI20PM1[2]\ : MX2
      port map(A => N_19, B => N_21, S => BIT_OS_SEL(1), Y => 
        N_35);
    
    \ADJ_Q[5]\ : DFN1C0
      port map(D => \ADJ_Q[3]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[5]_net_1\);
    
    \ARB_BYTE[1]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[1]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[1]_net_1\);
    
    \ARB_WRD_40M_FIXED[13]\ : DFN1C0
      port map(D => \Q[13]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[13]_net_1\);
    
    \ADJ_Q[0]\ : DFN1C0
      port map(D => \ADJ_SER_IN_R_1DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[0]_net_1\);
    
    \ARB_BYTE_RNI0QAI[13]\ : MX2
      port map(A => \ARB_BYTE[9]_net_1\, B => 
        \ARB_BYTE[13]_net_1\, S => BIT_OS_SEL(2), Y => N_32);
    
    \ARB_WRD_40M_FIXED[10]\ : DFN1C0
      port map(D => \Q[10]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[10]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SER320M_3_34_2 is

    port( ELK_TX_DAT                 : in    std_logic_vector(7 downto 0);
          MASTER_SALT_POR_B_i_0_i_5  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_13 : in    std_logic;
          ELK_OUT_R                  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_12 : in    std_logic;
          ELK_OUT_F                  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_8  : in    std_logic;
          CCC_160M_FXD               : in    std_logic;
          CLK_40M_GL                 : in    std_logic
        );

end SER320M_3_34_2;

architecture DEF_ARCH of SER320M_3_34_2 is 

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \N_SER_CMD_WORD_R[0]\, \START_RISE\, 
        \N_SER_CMD_WORD_F[0]\, \N_SER_CMD_WORD_R[3]\, 
        \SER_CMD_WORD_R[2]_net_1\, \N_SER_CMD_WORD_R[2]\, 
        \SER_CMD_WORD_R[1]_net_1\, \N_SER_CMD_WORD_R[1]\, 
        \SER_CMD_WORD_R[0]_net_1\, \N_SER_CMD_WORD_F[3]\, 
        \SER_CMD_WORD_F[2]_net_1\, \N_SER_CMD_WORD_F[2]\, 
        \SER_CMD_WORD_F[1]_net_1\, \N_SER_CMD_WORD_F[1]\, 
        \SER_CMD_WORD_F[0]_net_1\, N_START_RISE, 
        \CLK40M_GEN_DEL0\, \SER_OUT_FI\, \SER_OUT_RI\, 
        \SER_CMD_WORD_F[3]_net_1\, \SER_CMD_WORD_R[3]_net_1\, 
        \GND\, \VCC\ : std_logic;

begin 


    SER_OUT_FI : DFN1C0
      port map(D => \SER_CMD_WORD_F[3]_net_1\, CLK => 
        CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_5, Q => 
        \SER_OUT_FI\);
    
    \SER_CMD_WORD_F[3]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[3]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_12, Q => 
        \SER_CMD_WORD_F[3]_net_1\);
    
    \SER_CMD_WORD_R[1]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[1]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_8, Q => 
        \SER_CMD_WORD_R[1]_net_1\);
    
    \SER_CMD_WORD_R[2]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[2]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_8, Q => 
        \SER_CMD_WORD_R[2]_net_1\);
    
    \SER_CMD_WORD_R_RNO[3]\ : MX2
      port map(A => \SER_CMD_WORD_R[2]_net_1\, B => ELK_TX_DAT(7), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_R[3]\);
    
    \SER_CMD_WORD_R_RNO[0]\ : NOR2B
      port map(A => \START_RISE\, B => ELK_TX_DAT(1), Y => 
        \N_SER_CMD_WORD_R[0]\);
    
    \SER_CMD_WORD_F[0]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[0]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_12, Q => 
        \SER_CMD_WORD_F[0]_net_1\);
    
    \SER_CMD_WORD_R_RNO[1]\ : MX2
      port map(A => \SER_CMD_WORD_R[0]_net_1\, B => ELK_TX_DAT(3), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_R[1]\);
    
    \SER_CMD_WORD_F_RNO[2]\ : MX2
      port map(A => \SER_CMD_WORD_F[1]_net_1\, B => ELK_TX_DAT(4), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_F[2]\);
    
    \SER_CMD_WORD_F_RNO[3]\ : MX2
      port map(A => \SER_CMD_WORD_F[2]_net_1\, B => ELK_TX_DAT(6), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_F[3]\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    CLK40M_GEN_DEL0 : DFN1C0
      port map(D => CLK_40M_GL, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_8, Q => \CLK40M_GEN_DEL0\);
    
    SER_OUT_RI : DFN1C0
      port map(D => \SER_CMD_WORD_R[3]_net_1\, CLK => 
        CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_5, Q => 
        \SER_OUT_RI\);
    
    \SER_CMD_WORD_F[2]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[2]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_12, Q => 
        \SER_CMD_WORD_F[2]_net_1\);
    
    \SER_CMD_WORD_F_RNO[1]\ : MX2
      port map(A => \SER_CMD_WORD_F[0]_net_1\, B => ELK_TX_DAT(2), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_F[1]\);
    
    \SER_CMD_WORD_R[0]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[0]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_8, Q => 
        \SER_CMD_WORD_R[0]_net_1\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    START_RISE : DFN1C0
      port map(D => N_START_RISE, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_13, Q => \START_RISE\);
    
    \SER_CMD_WORD_R[3]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[3]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_8, Q => 
        \SER_CMD_WORD_R[3]_net_1\);
    
    \SER_CMD_WORD_F_RNO[0]\ : NOR2B
      port map(A => \START_RISE\, B => ELK_TX_DAT(0), Y => 
        \N_SER_CMD_WORD_F[0]\);
    
    SER_OUT_RDEL : DFN1C0
      port map(D => \SER_OUT_RI\, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_8, Q => ELK_OUT_R);
    
    \SER_CMD_WORD_F[1]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[1]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_12, Q => 
        \SER_CMD_WORD_F[1]_net_1\);
    
    START_RISE_RNO : NOR2B
      port map(A => \CLK40M_GEN_DEL0\, B => CLK_40M_GL, Y => 
        N_START_RISE);
    
    \SER_CMD_WORD_R_RNO[2]\ : MX2
      port map(A => \SER_CMD_WORD_R[1]_net_1\, B => ELK_TX_DAT(5), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_R[2]\);
    
    SER_OUT_FDEL : DFN1C0
      port map(D => \SER_OUT_FI\, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_12, Q => ELK_OUT_F);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity DDR_BIDIR_LVDS_DUAL_CLK_2 is

    port( DCB_SALT_SEL_c_i : in    std_logic;
          ELK2_DAT_P       : inout std_logic := 'Z';
          ELK2_DAT_N       : inout std_logic := 'Z';
          ELK_OUT_R        : in    std_logic;
          ELK_OUT_F        : in    std_logic;
          CCC_160M_FXD     : in    std_logic;
          CCC_160M_ADJ     : in    std_logic;
          ELK_IN_DDR_R     : out   std_logic;
          ELK_IN_DDR_F     : out   std_logic
        );

end DDR_BIDIR_LVDS_DUAL_CLK_2;

architecture DEF_ARCH of DDR_BIDIR_LVDS_DUAL_CLK_2 is 

  component DDR_REG
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          QR  : out   std_logic;
          QF  : out   std_logic
        );
  end component;

  component DDR_OUT
    port( DR  : in    std_logic := 'U';
          DF  : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component BIBUF_LVDS
    port( PADP : inout   std_logic;
          PADN : inout   std_logic;
          D    : in    std_logic := 'U';
          E    : in    std_logic := 'U';
          Y    : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal DDR_BIDIR_LVDS_DUAL_CLK_2_GND, BIBUF_LVDS_0_Y, 
        DDR_OUT_0_Q, \VCC\ : std_logic;

begin 


    DDR_REG_0 : DDR_REG
      port map(D => BIBUF_LVDS_0_Y, CLK => CCC_160M_ADJ, CLR => 
        DDR_BIDIR_LVDS_DUAL_CLK_2_GND, QR => ELK_IN_DDR_R, QF => 
        ELK_IN_DDR_F);
    
    DDR_OUT_0 : DDR_OUT
      port map(DR => ELK_OUT_R, DF => ELK_OUT_F, CLK => 
        CCC_160M_FXD, CLR => DDR_BIDIR_LVDS_DUAL_CLK_2_GND, Q => 
        DDR_OUT_0_Q);
    
    BIBUF_LVDS_0 : BIBUF_LVDS
      port map(PADP => ELK2_DAT_P, PADN => ELK2_DAT_N, D => 
        DDR_OUT_0_Q, E => DCB_SALT_SEL_c_i, Y => BIBUF_LVDS_0_Y);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    GND_i : GND
      port map(Y => DDR_BIDIR_LVDS_DUAL_CLK_2_GND);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SYNC_DAT_SEL_2 is

    port( ELK_TX_DAT                 : out   std_logic_vector(7 downto 0);
          PATT_ELK_DAT_2             : in    std_logic_vector(7 downto 0);
          OP_MODE_c_1_0              : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_13 : in    std_logic;
          CLK_40M_GL                 : in    std_logic
        );

end SYNC_DAT_SEL_2;

architecture DEF_ARCH of SYNC_DAT_SEL_2 is 

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \N_SERDAT[0]\, \N_SERDAT[1]\, \N_SERDAT[2]\, 
        \N_SERDAT[3]\, \N_SERDAT[4]\, \N_SERDAT[5]\, 
        \N_SERDAT[6]\, \N_SERDAT[7]\, \GND\, \VCC\ : std_logic;

begin 


    \SERDAT_RNO[4]\ : NOR2A
      port map(A => PATT_ELK_DAT_2(4), B => OP_MODE_c_1_0, Y => 
        \N_SERDAT[4]\);
    
    \SERDAT_RNO[0]\ : NOR2A
      port map(A => PATT_ELK_DAT_2(0), B => OP_MODE_c_1_0, Y => 
        \N_SERDAT[0]\);
    
    \SERDAT[6]\ : DFN1C0
      port map(D => \N_SERDAT[6]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_13, Q => ELK_TX_DAT(6));
    
    \SERDAT[4]\ : DFN1C0
      port map(D => \N_SERDAT[4]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_13, Q => ELK_TX_DAT(4));
    
    \SERDAT_RNO[7]\ : OR2
      port map(A => PATT_ELK_DAT_2(7), B => OP_MODE_c_1_0, Y => 
        \N_SERDAT[7]\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \SERDAT_RNO[3]\ : OR2
      port map(A => PATT_ELK_DAT_2(3), B => OP_MODE_c_1_0, Y => 
        \N_SERDAT[3]\);
    
    \SERDAT_RNO[2]\ : OR2
      port map(A => PATT_ELK_DAT_2(2), B => OP_MODE_c_1_0, Y => 
        \N_SERDAT[2]\);
    
    \SERDAT[5]\ : DFN1C0
      port map(D => \N_SERDAT[5]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_13, Q => ELK_TX_DAT(5));
    
    \SERDAT[7]\ : DFN1C0
      port map(D => \N_SERDAT[7]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_13, Q => ELK_TX_DAT(7));
    
    GND_i : GND
      port map(Y => \GND\);
    
    \SERDAT_RNO[5]\ : NOR2A
      port map(A => PATT_ELK_DAT_2(5), B => OP_MODE_c_1_0, Y => 
        \N_SERDAT[5]\);
    
    \SERDAT[0]\ : DFN1C0
      port map(D => \N_SERDAT[0]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_13, Q => ELK_TX_DAT(0));
    
    \SERDAT_RNO[6]\ : NOR2A
      port map(A => PATT_ELK_DAT_2(6), B => OP_MODE_c_1_0, Y => 
        \N_SERDAT[6]\);
    
    \SERDAT[1]\ : DFN1C0
      port map(D => \N_SERDAT[1]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_13, Q => ELK_TX_DAT(1));
    
    \SERDAT_RNO[1]\ : OR2
      port map(A => PATT_ELK_DAT_2(1), B => OP_MODE_c_1_0, Y => 
        \N_SERDAT[1]\);
    
    \SERDAT[3]\ : DFN1C0
      port map(D => \N_SERDAT[3]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_13, Q => ELK_TX_DAT(3));
    
    \SERDAT[2]\ : DFN1C0
      port map(D => \N_SERDAT[2]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_13, Q => ELK_TX_DAT(2));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity ELINK_SLAVE_15 is

    port( BIT_OS_SEL_7_0             : in    std_logic;
          BIT_OS_SEL                 : in    std_logic_vector(2 downto 1);
          BIT_OS_SEL_0_0             : in    std_logic;
          BIT_OS_SEL_1               : in    std_logic_vector(1 downto 0);
          ELK_RX_SER_WORD_2          : out   std_logic_vector(7 downto 0);
          OP_MODE_c_1_0              : in    std_logic;
          PATT_ELK_DAT_2             : in    std_logic_vector(7 downto 0);
          MASTER_DCB_POR_B_i_0_i     : in    std_logic;
          ELK2_DAT_N                 : inout std_logic := 'Z';
          ELK2_DAT_P                 : inout std_logic := 'Z';
          DCB_SALT_SEL_c_i           : in    std_logic;
          CCC_160M_FXD               : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_8  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_12 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_5  : in    std_logic;
          CLK_40M_GL                 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_13 : in    std_logic;
          DEV_RST_B_c_0              : in    std_logic;
          CCC_160M_ADJ               : in    std_logic
        );

end ELINK_SLAVE_15;

architecture DEF_ARCH of ELINK_SLAVE_15 is 

  component SLAVE_DES320S_1_17_0
    port( ELK_RX_SER_WORD_2      : out   std_logic_vector(7 downto 0);
          BIT_OS_SEL_1           : in    std_logic_vector(1 downto 0) := (others => 'U');
          BIT_OS_SEL_0_0         : in    std_logic := 'U';
          BIT_OS_SEL             : in    std_logic_vector(2 downto 1) := (others => 'U');
          BIT_OS_SEL_7_0         : in    std_logic := 'U';
          CLK_40M_GL             : in    std_logic := 'U';
          CCC_160M_FXD           : in    std_logic := 'U';
          ELK_IN_R               : in    std_logic := 'U';
          ELK_IN_F               : in    std_logic := 'U';
          MASTER_DCB_POR_B_i_0_i : in    std_logic := 'U';
          CCC_160M_ADJ           : in    std_logic := 'U'
        );
  end component;

  component SER320M_3_34_2
    port( ELK_TX_DAT                 : in    std_logic_vector(7 downto 0) := (others => 'U');
          MASTER_SALT_POR_B_i_0_i_5  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_13 : in    std_logic := 'U';
          ELK_OUT_R                  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_12 : in    std_logic := 'U';
          ELK_OUT_F                  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_8  : in    std_logic := 'U';
          CCC_160M_FXD               : in    std_logic := 'U';
          CLK_40M_GL                 : in    std_logic := 'U'
        );
  end component;

  component DDR_BIDIR_LVDS_DUAL_CLK_2
    port( DCB_SALT_SEL_c_i : in    std_logic := 'U';
          ELK2_DAT_P       : inout   std_logic;
          ELK2_DAT_N       : inout   std_logic;
          ELK_OUT_R        : in    std_logic := 'U';
          ELK_OUT_F        : in    std_logic := 'U';
          CCC_160M_FXD     : in    std_logic := 'U';
          CCC_160M_ADJ     : in    std_logic := 'U';
          ELK_IN_DDR_R     : out   std_logic;
          ELK_IN_DDR_F     : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component SYNC_DAT_SEL_2
    port( ELK_TX_DAT                 : out   std_logic_vector(7 downto 0);
          PATT_ELK_DAT_2             : in    std_logic_vector(7 downto 0) := (others => 'U');
          OP_MODE_c_1_0              : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_13 : in    std_logic := 'U';
          CLK_40M_GL                 : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \ELK_IN_F\, ELK_IN_DDR_F, \ELK_IN_R\, ELK_IN_DDR_R, 
        \ELK_TX_DAT[0]\, \ELK_TX_DAT[1]\, \ELK_TX_DAT[2]\, 
        \ELK_TX_DAT[3]\, \ELK_TX_DAT[4]\, \ELK_TX_DAT[5]\, 
        \ELK_TX_DAT[6]\, \ELK_TX_DAT[7]\, ELK_OUT_R, ELK_OUT_F, 
        \GND\, \VCC\ : std_logic;

    for all : SLAVE_DES320S_1_17_0
	Use entity work.SLAVE_DES320S_1_17_0(DEF_ARCH);
    for all : SER320M_3_34_2
	Use entity work.SER320M_3_34_2(DEF_ARCH);
    for all : DDR_BIDIR_LVDS_DUAL_CLK_2
	Use entity work.DDR_BIDIR_LVDS_DUAL_CLK_2(DEF_ARCH);
    for all : SYNC_DAT_SEL_2
	Use entity work.SYNC_DAT_SEL_2(DEF_ARCH);
begin 


    U_SLAVE_1ELK : SLAVE_DES320S_1_17_0
      port map(ELK_RX_SER_WORD_2(7) => ELK_RX_SER_WORD_2(7), 
        ELK_RX_SER_WORD_2(6) => ELK_RX_SER_WORD_2(6), 
        ELK_RX_SER_WORD_2(5) => ELK_RX_SER_WORD_2(5), 
        ELK_RX_SER_WORD_2(4) => ELK_RX_SER_WORD_2(4), 
        ELK_RX_SER_WORD_2(3) => ELK_RX_SER_WORD_2(3), 
        ELK_RX_SER_WORD_2(2) => ELK_RX_SER_WORD_2(2), 
        ELK_RX_SER_WORD_2(1) => ELK_RX_SER_WORD_2(1), 
        ELK_RX_SER_WORD_2(0) => ELK_RX_SER_WORD_2(0), 
        BIT_OS_SEL_1(1) => BIT_OS_SEL_1(1), BIT_OS_SEL_1(0) => 
        BIT_OS_SEL_1(0), BIT_OS_SEL_0_0 => BIT_OS_SEL_0_0, 
        BIT_OS_SEL(2) => BIT_OS_SEL(2), BIT_OS_SEL(1) => 
        BIT_OS_SEL(1), BIT_OS_SEL_7_0 => BIT_OS_SEL_7_0, 
        CLK_40M_GL => CLK_40M_GL, CCC_160M_FXD => CCC_160M_FXD, 
        ELK_IN_R => \ELK_IN_R\, ELK_IN_F => \ELK_IN_F\, 
        MASTER_DCB_POR_B_i_0_i => MASTER_DCB_POR_B_i_0_i, 
        CCC_160M_ADJ => CCC_160M_ADJ);
    
    U_ELK1_CMD_TX : SER320M_3_34_2
      port map(ELK_TX_DAT(7) => \ELK_TX_DAT[7]\, ELK_TX_DAT(6)
         => \ELK_TX_DAT[6]\, ELK_TX_DAT(5) => \ELK_TX_DAT[5]\, 
        ELK_TX_DAT(4) => \ELK_TX_DAT[4]\, ELK_TX_DAT(3) => 
        \ELK_TX_DAT[3]\, ELK_TX_DAT(2) => \ELK_TX_DAT[2]\, 
        ELK_TX_DAT(1) => \ELK_TX_DAT[1]\, ELK_TX_DAT(0) => 
        \ELK_TX_DAT[0]\, MASTER_SALT_POR_B_i_0_i_5 => 
        MASTER_SALT_POR_B_i_0_i_5, MASTER_SALT_POR_B_i_0_i_13 => 
        MASTER_SALT_POR_B_i_0_i_13, ELK_OUT_R => ELK_OUT_R, 
        MASTER_SALT_POR_B_i_0_i_12 => MASTER_SALT_POR_B_i_0_i_12, 
        ELK_OUT_F => ELK_OUT_F, MASTER_SALT_POR_B_i_0_i_8 => 
        MASTER_SALT_POR_B_i_0_i_8, CCC_160M_FXD => CCC_160M_FXD, 
        CLK_40M_GL => CLK_40M_GL);
    
    U_DDR_ELK1 : DDR_BIDIR_LVDS_DUAL_CLK_2
      port map(DCB_SALT_SEL_c_i => DCB_SALT_SEL_c_i, ELK2_DAT_P
         => ELK2_DAT_P, ELK2_DAT_N => ELK2_DAT_N, ELK_OUT_R => 
        ELK_OUT_R, ELK_OUT_F => ELK_OUT_F, CCC_160M_FXD => 
        CCC_160M_FXD, CCC_160M_ADJ => CCC_160M_ADJ, ELK_IN_DDR_R
         => ELK_IN_DDR_R, ELK_IN_DDR_F => ELK_IN_DDR_F);
    
    ELK_IN_F : DFN1C0
      port map(D => ELK_IN_DDR_F, CLK => CCC_160M_ADJ, CLR => 
        DEV_RST_B_c_0, Q => \ELK_IN_F\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    U_ELK1_SERDAT_SOURCE : SYNC_DAT_SEL_2
      port map(ELK_TX_DAT(7) => \ELK_TX_DAT[7]\, ELK_TX_DAT(6)
         => \ELK_TX_DAT[6]\, ELK_TX_DAT(5) => \ELK_TX_DAT[5]\, 
        ELK_TX_DAT(4) => \ELK_TX_DAT[4]\, ELK_TX_DAT(3) => 
        \ELK_TX_DAT[3]\, ELK_TX_DAT(2) => \ELK_TX_DAT[2]\, 
        ELK_TX_DAT(1) => \ELK_TX_DAT[1]\, ELK_TX_DAT(0) => 
        \ELK_TX_DAT[0]\, PATT_ELK_DAT_2(7) => PATT_ELK_DAT_2(7), 
        PATT_ELK_DAT_2(6) => PATT_ELK_DAT_2(6), PATT_ELK_DAT_2(5)
         => PATT_ELK_DAT_2(5), PATT_ELK_DAT_2(4) => 
        PATT_ELK_DAT_2(4), PATT_ELK_DAT_2(3) => PATT_ELK_DAT_2(3), 
        PATT_ELK_DAT_2(2) => PATT_ELK_DAT_2(2), PATT_ELK_DAT_2(1)
         => PATT_ELK_DAT_2(1), PATT_ELK_DAT_2(0) => 
        PATT_ELK_DAT_2(0), OP_MODE_c_1_0 => OP_MODE_c_1_0, 
        MASTER_SALT_POR_B_i_0_i_13 => MASTER_SALT_POR_B_i_0_i_13, 
        CLK_40M_GL => CLK_40M_GL);
    
    ELK_IN_R : DFN1C0
      port map(D => ELK_IN_DDR_R, CLK => CCC_160M_ADJ, CLR => 
        DEV_RST_B_c_0, Q => \ELK_IN_R\);
    
    GND_i : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SLAVE_DES320S_1_17_2 is

    port( ELK_RX_SER_WORD_4      : out   std_logic_vector(7 downto 0);
          BIT_OS_SEL_1_0         : in    std_logic;
          BIT_OS_SEL_0           : in    std_logic_vector(1 downto 0);
          BIT_OS_SEL_0_d0        : in    std_logic;
          BIT_OS_SEL_6           : in    std_logic_vector(2 downto 1);
          BIT_OS_SEL_7_0         : in    std_logic;
          CLK_40M_GL             : in    std_logic;
          CCC_160M_FXD           : in    std_logic;
          ELK_IN_R               : in    std_logic;
          ELK_IN_F               : in    std_logic;
          MASTER_DCB_POR_B_i_0_i : in    std_logic;
          CCC_160M_ADJ           : in    std_logic
        );

end SLAVE_DES320S_1_17_2;

architecture DEF_ARCH of SLAVE_DES320S_1_17_2 is 

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal N_17, \ARB_BYTE[0]_net_1\, \ARB_BYTE[4]_net_1\, N_18, 
        \ARB_BYTE[1]_net_1\, \ARB_BYTE[5]_net_1\, N_19, 
        \ARB_BYTE[2]_net_1\, \ARB_BYTE[6]_net_1\, N_20, 
        \ARB_BYTE[3]_net_1\, \ARB_BYTE[7]_net_1\, N_21, 
        \ARB_BYTE[8]_net_1\, N_22, \ARB_BYTE[9]_net_1\, N_23, 
        \ARB_BYTE[10]_net_1\, N_24, \ARB_BYTE[11]_net_1\, N_31, 
        \ARB_BYTE[12]_net_1\, N_32, \ARB_BYTE[13]_net_1\, N_33, 
        N_34, N_35, N_36, N_37, N_38, N_39, N_40, N_56, 
        \ARB_BYTE[14]_net_1\, N_64, \N_RECD_SER_WORD[0]\, 
        \N_RECD_SER_WORD[1]\, \N_RECD_SER_WORD[2]\, 
        \N_RECD_SER_WORD[3]\, \N_RECD_SER_WORD[4]\, 
        \N_RECD_SER_WORD[5]\, \N_RECD_SER_WORD[6]\, 
        \N_RECD_SER_WORD[7]\, \ADJ_SER_IN_F_0DEL\, 
        \ADJ_SER_IN_R_0DEL\, \ADJ_SER_IN_F_1DEL\, 
        \ADJ_SER_IN_R_1DEL\, \Q[0]_net_1\, \ADJ_Q[0]_net_1\, 
        \Q[1]_net_1\, \ADJ_Q[1]_net_1\, \Q[2]_net_1\, 
        \ADJ_Q[2]_net_1\, \Q[3]_net_1\, \ADJ_Q[3]_net_1\, 
        \Q[4]_net_1\, \ADJ_Q[4]_net_1\, \Q[5]_net_1\, 
        \ADJ_Q[5]_net_1\, \Q[6]_net_1\, \ADJ_Q[6]_net_1\, 
        \Q[7]_net_1\, \ADJ_Q[7]_net_1\, \Q[8]_net_1\, 
        \ADJ_Q[8]_net_1\, \Q[9]_net_1\, \ADJ_Q[9]_net_1\, 
        \Q[10]_net_1\, \ADJ_Q[10]_net_1\, \Q[11]_net_1\, 
        \ADJ_Q[11]_net_1\, \Q[12]_net_1\, \ADJ_Q[12]_net_1\, 
        \Q[13]_net_1\, \ADJ_Q[13]_net_1\, \Q[14]_net_1\, 
        \ADJ_Q[14]_net_1\, \ARB_WRD_40M_FIXED[0]_net_1\, 
        \ARB_WRD_40M_FIXED[1]_net_1\, 
        \ARB_WRD_40M_FIXED[2]_net_1\, 
        \ARB_WRD_40M_FIXED[3]_net_1\, 
        \ARB_WRD_40M_FIXED[4]_net_1\, 
        \ARB_WRD_40M_FIXED[5]_net_1\, 
        \ARB_WRD_40M_FIXED[6]_net_1\, 
        \ARB_WRD_40M_FIXED[7]_net_1\, 
        \ARB_WRD_40M_FIXED[8]_net_1\, 
        \ARB_WRD_40M_FIXED[9]_net_1\, 
        \ARB_WRD_40M_FIXED[10]_net_1\, 
        \ARB_WRD_40M_FIXED[11]_net_1\, 
        \ARB_WRD_40M_FIXED[12]_net_1\, 
        \ARB_WRD_40M_FIXED[13]_net_1\, 
        \ARB_WRD_40M_FIXED[14]_net_1\, \GND\, \VCC\ : std_logic;

begin 


    \RECD_SER_WORD_RNO[5]\ : MX2
      port map(A => N_38, B => N_39, S => BIT_OS_SEL_0(0), Y => 
        \N_RECD_SER_WORD[5]\);
    
    \ARB_WRD_40M_FIXED[9]\ : DFN1C0
      port map(D => \Q[9]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[9]_net_1\);
    
    \ADJ_Q[4]\ : DFN1C0
      port map(D => \ADJ_Q[2]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[4]_net_1\);
    
    \ARB_BYTE[6]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[6]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[6]_net_1\);
    
    ADJ_SER_IN_F_1DEL : DFN1C0
      port map(D => \ADJ_SER_IN_F_0DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_F_1DEL\);
    
    \ARB_BYTE[0]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[0]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[0]_net_1\);
    
    \Q[11]\ : DFN1C0
      port map(D => \ADJ_Q[11]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[11]_net_1\);
    
    \ADJ_Q[8]\ : DFN1C0
      port map(D => \ADJ_Q[6]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[8]_net_1\);
    
    \ADJ_Q[6]\ : DFN1C0
      port map(D => \ADJ_Q[4]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[6]_net_1\);
    
    \ADJ_Q[12]\ : DFN1C0
      port map(D => \ADJ_Q[10]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[12]_net_1\);
    
    \RECD_SER_WORD_RNO_1[0]\ : MX2
      port map(A => \ARB_BYTE[0]_net_1\, B => \ARB_BYTE[4]_net_1\, 
        S => BIT_OS_SEL_6(2), Y => N_17);
    
    \ARB_BYTE_RNI89ML[4]\ : MX2
      port map(A => \ARB_BYTE[4]_net_1\, B => \ARB_BYTE[8]_net_1\, 
        S => BIT_OS_SEL_6(2), Y => N_21);
    
    \Q[1]\ : DFN1C0
      port map(D => \ADJ_Q[1]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[1]_net_1\);
    
    \ARB_BYTE[4]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[4]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[4]_net_1\);
    
    \ADJ_Q[2]\ : DFN1C0
      port map(D => \ADJ_Q[0]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[2]_net_1\);
    
    \RECD_SER_WORD_RNO_1[7]\ : MX2
      port map(A => \ARB_BYTE[10]_net_1\, B => 
        \ARB_BYTE[14]_net_1\, S => BIT_OS_SEL_0_d0, Y => N_56);
    
    \RECD_SER_WORD[4]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[4]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_4(4));
    
    \Q[5]\ : DFN1C0
      port map(D => \ADJ_Q[5]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[5]_net_1\);
    
    \ADJ_Q[11]\ : DFN1C0
      port map(D => \ADJ_Q[9]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[11]_net_1\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \ADJ_Q[3]\ : DFN1C0
      port map(D => \ADJ_Q[1]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[3]_net_1\);
    
    \Q[10]\ : DFN1C0
      port map(D => \ADJ_Q[10]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[10]_net_1\);
    
    \ARB_WRD_40M_FIXED[6]\ : DFN1C0
      port map(D => \Q[6]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[6]_net_1\);
    
    \ARB_WRD_40M_FIXED[1]\ : DFN1C0
      port map(D => \Q[1]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[1]_net_1\);
    
    \RECD_SER_WORD[3]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[3]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_4(3));
    
    \RECD_SER_WORD[0]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[0]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_4(0));
    
    \RECD_SER_WORD_RNO[3]\ : MX2
      port map(A => N_36, B => N_37, S => BIT_OS_SEL_0(0), Y => 
        \N_RECD_SER_WORD[3]\);
    
    \Q[0]\ : DFN1C0
      port map(D => \ADJ_Q[0]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[0]_net_1\);
    
    \ARB_BYTE_RNI0TEE1[13]\ : MX2
      port map(A => N_24, B => N_32, S => BIT_OS_SEL_6(1), Y => 
        N_40);
    
    \ARB_BYTE_RNILG9K[11]\ : MX2
      port map(A => \ARB_BYTE[7]_net_1\, B => 
        \ARB_BYTE[11]_net_1\, S => BIT_OS_SEL_6(2), Y => N_24);
    
    \RECD_SER_WORD_RNO_0[7]\ : MX2
      port map(A => N_31, B => N_56, S => BIT_OS_SEL_0(1), Y => 
        N_64);
    
    \Q[7]\ : DFN1C0
      port map(D => \ADJ_Q[7]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[7]_net_1\);
    
    \ARB_BYTE[14]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[14]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[14]_net_1\);
    
    \ARB_WRD_40M_FIXED[2]\ : DFN1C0
      port map(D => \Q[2]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[2]_net_1\);
    
    \ARB_WRD_40M_FIXED[14]\ : DFN1C0
      port map(D => \Q[14]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[14]_net_1\);
    
    \RECD_SER_WORD_RNO[2]\ : MX2
      port map(A => N_35, B => N_36, S => BIT_OS_SEL_0(0), Y => 
        \N_RECD_SER_WORD[2]\);
    
    \ARB_BYTE_RNIRLBD1[10]\ : MX2
      port map(A => N_23, B => N_31, S => BIT_OS_SEL_6(1), Y => 
        N_39);
    
    \ARB_BYTE[2]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[2]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[2]_net_1\);
    
    \ADJ_Q[7]\ : DFN1C0
      port map(D => \ADJ_Q[5]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[7]_net_1\);
    
    \ARB_BYTE[8]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[8]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[8]_net_1\);
    
    \RECD_SER_WORD[5]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[5]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_4(5));
    
    \ARB_BYTE[12]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[12]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[12]_net_1\);
    
    \ARB_BYTE_RNINI9K[12]\ : MX2
      port map(A => \ARB_BYTE[8]_net_1\, B => 
        \ARB_BYTE[12]_net_1\, S => BIT_OS_SEL_6(2), Y => N_31);
    
    \RECD_SER_WORD[1]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[1]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_4(1));
    
    \ARB_BYTE_RNIJE9K[10]\ : MX2
      port map(A => \ARB_BYTE[6]_net_1\, B => 
        \ARB_BYTE[10]_net_1\, S => BIT_OS_SEL_6(2), Y => N_23);
    
    \Q[3]\ : DFN1C0
      port map(D => \ADJ_Q[3]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[3]_net_1\);
    
    \ARB_BYTE_RNI23ML[1]\ : MX2
      port map(A => \ARB_BYTE[1]_net_1\, B => \ARB_BYTE[5]_net_1\, 
        S => BIT_OS_SEL_6(2), Y => N_18);
    
    ADJ_SER_IN_F_0DEL : DFN1C0
      port map(D => ELK_IN_F, CLK => CCC_160M_ADJ, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_F_0DEL\);
    
    \RECD_SER_WORD_RNO[7]\ : MX2
      port map(A => N_40, B => N_64, S => BIT_OS_SEL_1_0, Y => 
        \N_RECD_SER_WORD[7]\);
    
    \RECD_SER_WORD_RNO[1]\ : MX2
      port map(A => N_34, B => N_35, S => BIT_OS_SEL_0(0), Y => 
        \N_RECD_SER_WORD[1]\);
    
    \ARB_WRD_40M_FIXED[4]\ : DFN1C0
      port map(D => \Q[4]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[4]_net_1\);
    
    \RECD_SER_WORD_RNO[0]\ : MX2
      port map(A => N_33, B => N_34, S => BIT_OS_SEL_0(0), Y => 
        \N_RECD_SER_WORD[0]\);
    
    \Q[6]\ : DFN1C0
      port map(D => \ADJ_Q[6]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[6]_net_1\);
    
    \ARB_BYTE_RNIGGOE1[11]\ : MX2
      port map(A => N_22, B => N_24, S => BIT_OS_SEL_6(1), Y => 
        N_38);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \ARB_WRD_40M_FIXED[8]\ : DFN1C0
      port map(D => \Q[8]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[8]_net_1\);
    
    \ARB_BYTE[11]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[11]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[11]_net_1\);
    
    \Q[9]\ : DFN1C0
      port map(D => \ADJ_Q[9]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[9]_net_1\);
    
    \Q[14]\ : DFN1C0
      port map(D => \ADJ_Q[14]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[14]_net_1\);
    
    ADJ_SER_IN_R_0DEL : DFN1C0
      port map(D => ELK_IN_R, CLK => CCC_160M_ADJ, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_R_0DEL\);
    
    \Q[13]\ : DFN1C0
      port map(D => \ADJ_Q[13]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[13]_net_1\);
    
    \ARB_BYTE[9]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[9]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[9]_net_1\);
    
    ADJ_SER_IN_R_1DEL : DFN1C0
      port map(D => \ADJ_SER_IN_R_0DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_R_1DEL\);
    
    \ARB_BYTE[10]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[10]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[10]_net_1\);
    
    \ADJ_Q[9]\ : DFN1C0
      port map(D => \ADJ_Q[7]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[9]_net_1\);
    
    \RECD_SER_WORD[7]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[7]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_4(7));
    
    \ARB_WRD_40M_FIXED[5]\ : DFN1C0
      port map(D => \Q[5]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[5]_net_1\);
    
    \ARB_WRD_40M_FIXED[12]\ : DFN1C0
      port map(D => \Q[12]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[12]_net_1\);
    
    \ARB_BYTE_RNIPU4G1[1]\ : MX2
      port map(A => N_18, B => N_20, S => BIT_OS_SEL_6(1), Y => 
        N_34);
    
    \ARB_WRD_40M_FIXED[11]\ : DFN1C0
      port map(D => \Q[11]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[11]_net_1\);
    
    \ARB_WRD_40M_FIXED[0]\ : DFN1C0
      port map(D => \Q[0]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[0]_net_1\);
    
    \ADJ_Q[10]\ : DFN1C0
      port map(D => \ADJ_Q[8]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[10]_net_1\);
    
    \Q[2]\ : DFN1C0
      port map(D => \ADJ_Q[2]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[2]_net_1\);
    
    \ADJ_Q[1]\ : DFN1C0
      port map(D => \ADJ_SER_IN_F_1DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[1]_net_1\);
    
    \RECD_SER_WORD[6]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[6]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_4(6));
    
    \RECD_SER_WORD[2]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[2]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_4(2));
    
    \ARB_BYTE_RNI67ML[3]\ : MX2
      port map(A => \ARB_BYTE[3]_net_1\, B => \ARB_BYTE[7]_net_1\, 
        S => BIT_OS_SEL_6(2), Y => N_20);
    
    \ADJ_Q[13]\ : DFN1C0
      port map(D => \ADJ_Q[11]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[13]_net_1\);
    
    \ARB_BYTE_RNIT25G1[2]\ : MX2
      port map(A => N_19, B => N_21, S => BIT_OS_SEL_6(1), Y => 
        N_35);
    
    \Q[8]\ : DFN1C0
      port map(D => \ADJ_Q[8]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[8]_net_1\);
    
    \ARB_BYTE[5]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[5]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[5]_net_1\);
    
    \ADJ_Q[14]\ : DFN1C0
      port map(D => \ADJ_Q[12]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[14]_net_1\);
    
    \ARB_BYTE_RNI45ML[2]\ : MX2
      port map(A => \ARB_BYTE[2]_net_1\, B => \ARB_BYTE[6]_net_1\, 
        S => BIT_OS_SEL_6(2), Y => N_19);
    
    \RECD_SER_WORD_RNO[4]\ : MX2
      port map(A => N_37, B => N_38, S => BIT_OS_SEL_0(0), Y => 
        \N_RECD_SER_WORD[4]\);
    
    \Q[12]\ : DFN1C0
      port map(D => \ADJ_Q[12]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[12]_net_1\);
    
    \ARB_BYTE_RNIABML[5]\ : MX2
      port map(A => \ARB_BYTE[5]_net_1\, B => \ARB_BYTE[9]_net_1\, 
        S => BIT_OS_SEL_6(2), Y => N_22);
    
    \ARB_BYTE[13]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[13]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[13]_net_1\);
    
    \ARB_WRD_40M_FIXED[3]\ : DFN1C0
      port map(D => \Q[3]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[3]_net_1\);
    
    \ARB_BYTE[7]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[7]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[7]_net_1\);
    
    \RECD_SER_WORD_RNO_0[0]\ : MX2
      port map(A => N_17, B => N_19, S => BIT_OS_SEL_6(1), Y => 
        N_33);
    
    \Q[4]\ : DFN1C0
      port map(D => \ADJ_Q[4]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[4]_net_1\);
    
    \ARB_WRD_40M_FIXED[7]\ : DFN1C0
      port map(D => \Q[7]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[7]_net_1\);
    
    \RECD_SER_WORD_RNO[6]\ : MX2
      port map(A => N_39, B => N_40, S => BIT_OS_SEL_0(0), Y => 
        \N_RECD_SER_WORD[6]\);
    
    \ARB_BYTE_RNICCOE1[10]\ : MX2
      port map(A => N_21, B => N_23, S => BIT_OS_SEL_6(1), Y => 
        N_37);
    
    \ARB_BYTE[3]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[3]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[3]_net_1\);
    
    \ADJ_Q[5]\ : DFN1C0
      port map(D => \ADJ_Q[3]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[5]_net_1\);
    
    \ARB_BYTE[1]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[1]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[1]_net_1\);
    
    \ARB_BYTE_RNI175G1[3]\ : MX2
      port map(A => N_20, B => N_22, S => BIT_OS_SEL_6(1), Y => 
        N_36);
    
    \ARB_WRD_40M_FIXED[13]\ : DFN1C0
      port map(D => \Q[13]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[13]_net_1\);
    
    \ADJ_Q[0]\ : DFN1C0
      port map(D => \ADJ_SER_IN_R_1DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[0]_net_1\);
    
    \ARB_BYTE_RNIQNCL[13]\ : MX2
      port map(A => \ARB_BYTE[9]_net_1\, B => 
        \ARB_BYTE[13]_net_1\, S => BIT_OS_SEL_7_0, Y => N_32);
    
    \ARB_WRD_40M_FIXED[10]\ : DFN1C0
      port map(D => \Q[10]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[10]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SER320M_3_34_4 is

    port( ELK_TX_DAT                 : in    std_logic_vector(7 downto 0);
          MASTER_SALT_POR_B_i_0_i_17 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_1  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_13 : in    std_logic;
          ELK_OUT_R_i_0              : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_16 : in    std_logic;
          ELK_OUT_F_i_0              : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_9  : in    std_logic;
          CLK_40M_GL                 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_4  : in    std_logic;
          CCC_160M_FXD               : in    std_logic
        );

end SER320M_3_34_4;

architecture DEF_ARCH of SER320M_3_34_4 is 

  component DFI1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          QN  : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component DFN1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

    signal SER_OUT_RI_i, \SER_CMD_WORD_R[3]_net_1\, SER_OUT_FI_i, 
        \SER_CMD_WORD_F[3]_net_1\, \N_SER_CMD_WORD_R[0]\, 
        \START_RISE\, \N_SER_CMD_WORD_F[0]\, 
        \N_SER_CMD_WORD_R[3]\, \SER_CMD_WORD_R[2]_net_1\, 
        \N_SER_CMD_WORD_R[2]\, \SER_CMD_WORD_R[1]_net_1\, 
        \N_SER_CMD_WORD_R[1]\, \SER_CMD_WORD_R[0]_net_1\, 
        \N_SER_CMD_WORD_F[3]\, \SER_CMD_WORD_F[2]_net_1\, 
        \N_SER_CMD_WORD_F[2]\, \SER_CMD_WORD_F[1]_net_1\, 
        \N_SER_CMD_WORD_F[1]\, \SER_CMD_WORD_F[0]_net_1\, 
        N_START_RISE, \CLK40M_GEN_DEL0\, \GND\, \VCC\
         : std_logic;

begin 


    SER_OUT_FI : DFI1C0
      port map(D => \SER_CMD_WORD_F[3]_net_1\, CLK => 
        CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_4, QN => 
        SER_OUT_FI_i);
    
    \SER_CMD_WORD_F[3]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[3]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_1, Q => 
        \SER_CMD_WORD_F[3]_net_1\);
    
    \SER_CMD_WORD_R[1]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[1]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_17, Q => 
        \SER_CMD_WORD_R[1]_net_1\);
    
    \SER_CMD_WORD_R[2]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[2]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_17, Q => 
        \SER_CMD_WORD_R[2]_net_1\);
    
    \SER_CMD_WORD_R_RNO[3]\ : MX2
      port map(A => \SER_CMD_WORD_R[2]_net_1\, B => ELK_TX_DAT(7), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_R[3]\);
    
    \SER_CMD_WORD_R_RNO[0]\ : NOR2B
      port map(A => \START_RISE\, B => ELK_TX_DAT(1), Y => 
        \N_SER_CMD_WORD_R[0]\);
    
    \SER_CMD_WORD_F[0]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[0]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_1, Q => 
        \SER_CMD_WORD_F[0]_net_1\);
    
    \SER_CMD_WORD_R_RNO[1]\ : MX2
      port map(A => \SER_CMD_WORD_R[0]_net_1\, B => ELK_TX_DAT(3), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_R[1]\);
    
    \SER_CMD_WORD_F_RNO[2]\ : MX2
      port map(A => \SER_CMD_WORD_F[1]_net_1\, B => ELK_TX_DAT(4), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_F[2]\);
    
    \SER_CMD_WORD_F_RNO[3]\ : MX2
      port map(A => \SER_CMD_WORD_F[2]_net_1\, B => ELK_TX_DAT(6), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_F[3]\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    CLK40M_GEN_DEL0 : DFN1C0
      port map(D => CLK_40M_GL, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_9, Q => \CLK40M_GEN_DEL0\);
    
    SER_OUT_RI : DFI1C0
      port map(D => \SER_CMD_WORD_R[3]_net_1\, CLK => 
        CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_4, QN => 
        SER_OUT_RI_i);
    
    \SER_CMD_WORD_F[2]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[2]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_1, Q => 
        \SER_CMD_WORD_F[2]_net_1\);
    
    \SER_CMD_WORD_F_RNO[1]\ : MX2
      port map(A => \SER_CMD_WORD_F[0]_net_1\, B => ELK_TX_DAT(2), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_F[1]\);
    
    \SER_CMD_WORD_R[0]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[0]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_16, Q => 
        \SER_CMD_WORD_R[0]_net_1\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    START_RISE : DFN1C0
      port map(D => N_START_RISE, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_13, Q => \START_RISE\);
    
    \SER_CMD_WORD_R[3]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[3]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_17, Q => 
        \SER_CMD_WORD_R[3]_net_1\);
    
    \SER_CMD_WORD_F_RNO[0]\ : NOR2B
      port map(A => \START_RISE\, B => ELK_TX_DAT(0), Y => 
        \N_SER_CMD_WORD_F[0]\);
    
    SER_OUT_RDEL : DFN1P0
      port map(D => SER_OUT_RI_i, CLK => CCC_160M_FXD, PRE => 
        MASTER_SALT_POR_B_i_0_i_13, Q => ELK_OUT_R_i_0);
    
    \SER_CMD_WORD_F[1]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[1]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_1, Q => 
        \SER_CMD_WORD_F[1]_net_1\);
    
    START_RISE_RNO : NOR2B
      port map(A => \CLK40M_GEN_DEL0\, B => CLK_40M_GL, Y => 
        N_START_RISE);
    
    \SER_CMD_WORD_R_RNO[2]\ : MX2
      port map(A => \SER_CMD_WORD_R[1]_net_1\, B => ELK_TX_DAT(5), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_R[2]\);
    
    SER_OUT_FDEL : DFN1P0
      port map(D => SER_OUT_FI_i, CLK => CCC_160M_FXD, PRE => 
        MASTER_SALT_POR_B_i_0_i_16, Q => ELK_OUT_F_i_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity DDR_BIDIR_LVDS_DUAL_CLK_4 is

    port( DCB_SALT_SEL_c_i : in    std_logic;
          ELK4_DAT_P       : inout std_logic := 'Z';
          ELK4_DAT_N       : inout std_logic := 'Z';
          ELK_OUT_R_i_0    : in    std_logic;
          ELK_OUT_F_i_0    : in    std_logic;
          CCC_160M_FXD     : in    std_logic;
          CCC_160M_ADJ     : in    std_logic;
          ELK_IN_DDR_F_i   : out   std_logic;
          ELK_IN_DDR_R_i   : out   std_logic
        );

end DDR_BIDIR_LVDS_DUAL_CLK_4;

architecture DEF_ARCH of DDR_BIDIR_LVDS_DUAL_CLK_4 is 

  component INV
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DDR_REG
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          QR  : out   std_logic;
          QF  : out   std_logic
        );
  end component;

  component DDR_OUT
    port( DR  : in    std_logic := 'U';
          DF  : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component BIBUF_LVDS
    port( PADP : inout   std_logic;
          PADN : inout   std_logic;
          D    : in    std_logic := 'U';
          E    : in    std_logic := 'U';
          Y    : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal ELK_IN_DDR_R, ELK_IN_DDR_F, 
        DDR_BIDIR_LVDS_DUAL_CLK_4_GND, BIBUF_LVDS_0_Y, 
        DDR_OUT_0_Q, \VCC\ : std_logic;

begin 


    DDR_REG_0_RNIA1NA : INV
      port map(A => ELK_IN_DDR_F, Y => ELK_IN_DDR_F_i);
    
    DDR_REG_0 : DDR_REG
      port map(D => BIBUF_LVDS_0_Y, CLK => CCC_160M_ADJ, CLR => 
        DDR_BIDIR_LVDS_DUAL_CLK_4_GND, QR => ELK_IN_DDR_R, QF => 
        ELK_IN_DDR_F);
    
    DDR_OUT_0 : DDR_OUT
      port map(DR => ELK_OUT_R_i_0, DF => ELK_OUT_F_i_0, CLK => 
        CCC_160M_FXD, CLR => DDR_BIDIR_LVDS_DUAL_CLK_4_GND, Q => 
        DDR_OUT_0_Q);
    
    BIBUF_LVDS_0 : BIBUF_LVDS
      port map(PADP => ELK4_DAT_P, PADN => ELK4_DAT_N, D => 
        DDR_OUT_0_Q, E => DCB_SALT_SEL_c_i, Y => BIBUF_LVDS_0_Y);
    
    DDR_REG_0_RNIA1NA_0 : INV
      port map(A => ELK_IN_DDR_R, Y => ELK_IN_DDR_R_i);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    GND_i : GND
      port map(Y => DDR_BIDIR_LVDS_DUAL_CLK_4_GND);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SYNC_DAT_SEL_4 is

    port( ELK_TX_DAT                 : out   std_logic_vector(7 downto 0);
          PATT_ELK_DAT_4             : in    std_logic_vector(7 downto 0);
          OP_MODE_c_1_0              : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_16 : in    std_logic;
          CLK_40M_GL                 : in    std_logic
        );

end SYNC_DAT_SEL_4;

architecture DEF_ARCH of SYNC_DAT_SEL_4 is 

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \N_SERDAT[0]\, \N_SERDAT[1]\, \N_SERDAT[2]\, 
        \N_SERDAT[3]\, \N_SERDAT[4]\, \N_SERDAT[5]\, 
        \N_SERDAT[6]\, \N_SERDAT[7]\, \GND\, \VCC\ : std_logic;

begin 


    \SERDAT_RNO[4]\ : NOR2A
      port map(A => PATT_ELK_DAT_4(4), B => OP_MODE_c_1_0, Y => 
        \N_SERDAT[4]\);
    
    \SERDAT_RNO[0]\ : NOR2A
      port map(A => PATT_ELK_DAT_4(0), B => OP_MODE_c_1_0, Y => 
        \N_SERDAT[0]\);
    
    \SERDAT[6]\ : DFN1C0
      port map(D => \N_SERDAT[6]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_16, Q => ELK_TX_DAT(6));
    
    \SERDAT[4]\ : DFN1C0
      port map(D => \N_SERDAT[4]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_16, Q => ELK_TX_DAT(4));
    
    \SERDAT_RNO[7]\ : OR2
      port map(A => PATT_ELK_DAT_4(7), B => OP_MODE_c_1_0, Y => 
        \N_SERDAT[7]\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \SERDAT_RNO[3]\ : OR2
      port map(A => PATT_ELK_DAT_4(3), B => OP_MODE_c_1_0, Y => 
        \N_SERDAT[3]\);
    
    \SERDAT_RNO[2]\ : OR2
      port map(A => PATT_ELK_DAT_4(2), B => OP_MODE_c_1_0, Y => 
        \N_SERDAT[2]\);
    
    \SERDAT[5]\ : DFN1C0
      port map(D => \N_SERDAT[5]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_16, Q => ELK_TX_DAT(5));
    
    \SERDAT[7]\ : DFN1C0
      port map(D => \N_SERDAT[7]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_16, Q => ELK_TX_DAT(7));
    
    GND_i : GND
      port map(Y => \GND\);
    
    \SERDAT_RNO[5]\ : NOR2A
      port map(A => PATT_ELK_DAT_4(5), B => OP_MODE_c_1_0, Y => 
        \N_SERDAT[5]\);
    
    \SERDAT[0]\ : DFN1C0
      port map(D => \N_SERDAT[0]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_16, Q => ELK_TX_DAT(0));
    
    \SERDAT_RNO[6]\ : NOR2A
      port map(A => PATT_ELK_DAT_4(6), B => OP_MODE_c_1_0, Y => 
        \N_SERDAT[6]\);
    
    \SERDAT[1]\ : DFN1C0
      port map(D => \N_SERDAT[1]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_16, Q => ELK_TX_DAT(1));
    
    \SERDAT_RNO[1]\ : OR2
      port map(A => PATT_ELK_DAT_4(1), B => OP_MODE_c_1_0, Y => 
        \N_SERDAT[1]\);
    
    \SERDAT[3]\ : DFN1C0
      port map(D => \N_SERDAT[3]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_16, Q => ELK_TX_DAT(3));
    
    \SERDAT[2]\ : DFN1C0
      port map(D => \N_SERDAT[2]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_16, Q => ELK_TX_DAT(2));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity ELINK_SLAVE_INV_2_1 is

    port( BIT_OS_SEL_7_0             : in    std_logic;
          BIT_OS_SEL_6               : in    std_logic_vector(2 downto 1);
          BIT_OS_SEL_0_d0            : in    std_logic;
          BIT_OS_SEL_0               : in    std_logic_vector(1 downto 0);
          BIT_OS_SEL_1_0             : in    std_logic;
          ELK_RX_SER_WORD_4          : out   std_logic_vector(7 downto 0);
          OP_MODE_c_1_0              : in    std_logic;
          PATT_ELK_DAT_4             : in    std_logic_vector(7 downto 0);
          MASTER_DCB_POR_B_i_0_i     : in    std_logic;
          ELK4_DAT_N                 : inout std_logic := 'Z';
          ELK4_DAT_P                 : inout std_logic := 'Z';
          DCB_SALT_SEL_c_i           : in    std_logic;
          CCC_160M_FXD               : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_4  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_9  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_13 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_1  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_17 : in    std_logic;
          CLK_40M_GL                 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_16 : in    std_logic;
          DEV_RST_B_c                : in    std_logic;
          CCC_160M_ADJ               : in    std_logic
        );

end ELINK_SLAVE_INV_2_1;

architecture DEF_ARCH of ELINK_SLAVE_INV_2_1 is 

  component SLAVE_DES320S_1_17_2
    port( ELK_RX_SER_WORD_4      : out   std_logic_vector(7 downto 0);
          BIT_OS_SEL_1_0         : in    std_logic := 'U';
          BIT_OS_SEL_0           : in    std_logic_vector(1 downto 0) := (others => 'U');
          BIT_OS_SEL_0_d0        : in    std_logic := 'U';
          BIT_OS_SEL_6           : in    std_logic_vector(2 downto 1) := (others => 'U');
          BIT_OS_SEL_7_0         : in    std_logic := 'U';
          CLK_40M_GL             : in    std_logic := 'U';
          CCC_160M_FXD           : in    std_logic := 'U';
          ELK_IN_R               : in    std_logic := 'U';
          ELK_IN_F               : in    std_logic := 'U';
          MASTER_DCB_POR_B_i_0_i : in    std_logic := 'U';
          CCC_160M_ADJ           : in    std_logic := 'U'
        );
  end component;

  component SER320M_3_34_4
    port( ELK_TX_DAT                 : in    std_logic_vector(7 downto 0) := (others => 'U');
          MASTER_SALT_POR_B_i_0_i_17 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_1  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_13 : in    std_logic := 'U';
          ELK_OUT_R_i_0              : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_16 : in    std_logic := 'U';
          ELK_OUT_F_i_0              : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_9  : in    std_logic := 'U';
          CLK_40M_GL                 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_4  : in    std_logic := 'U';
          CCC_160M_FXD               : in    std_logic := 'U'
        );
  end component;

  component DDR_BIDIR_LVDS_DUAL_CLK_4
    port( DCB_SALT_SEL_c_i : in    std_logic := 'U';
          ELK4_DAT_P       : inout   std_logic;
          ELK4_DAT_N       : inout   std_logic;
          ELK_OUT_R_i_0    : in    std_logic := 'U';
          ELK_OUT_F_i_0    : in    std_logic := 'U';
          CCC_160M_FXD     : in    std_logic := 'U';
          CCC_160M_ADJ     : in    std_logic := 'U';
          ELK_IN_DDR_F_i   : out   std_logic;
          ELK_IN_DDR_R_i   : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component SYNC_DAT_SEL_4
    port( ELK_TX_DAT                 : out   std_logic_vector(7 downto 0);
          PATT_ELK_DAT_4             : in    std_logic_vector(7 downto 0) := (others => 'U');
          OP_MODE_c_1_0              : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_16 : in    std_logic := 'U';
          CLK_40M_GL                 : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \ELK_IN_F\, ELK_IN_DDR_F_i, \ELK_IN_R\, 
        ELK_IN_DDR_R_i, \ELK_TX_DAT[0]\, \ELK_TX_DAT[1]\, 
        \ELK_TX_DAT[2]\, \ELK_TX_DAT[3]\, \ELK_TX_DAT[4]\, 
        \ELK_TX_DAT[5]\, \ELK_TX_DAT[6]\, \ELK_TX_DAT[7]\, 
        ELK_OUT_R_i_0, ELK_OUT_F_i_0, \GND\, \VCC\ : std_logic;

    for all : SLAVE_DES320S_1_17_2
	Use entity work.SLAVE_DES320S_1_17_2(DEF_ARCH);
    for all : SER320M_3_34_4
	Use entity work.SER320M_3_34_4(DEF_ARCH);
    for all : DDR_BIDIR_LVDS_DUAL_CLK_4
	Use entity work.DDR_BIDIR_LVDS_DUAL_CLK_4(DEF_ARCH);
    for all : SYNC_DAT_SEL_4
	Use entity work.SYNC_DAT_SEL_4(DEF_ARCH);
begin 


    U_SLAVE_1ELK : SLAVE_DES320S_1_17_2
      port map(ELK_RX_SER_WORD_4(7) => ELK_RX_SER_WORD_4(7), 
        ELK_RX_SER_WORD_4(6) => ELK_RX_SER_WORD_4(6), 
        ELK_RX_SER_WORD_4(5) => ELK_RX_SER_WORD_4(5), 
        ELK_RX_SER_WORD_4(4) => ELK_RX_SER_WORD_4(4), 
        ELK_RX_SER_WORD_4(3) => ELK_RX_SER_WORD_4(3), 
        ELK_RX_SER_WORD_4(2) => ELK_RX_SER_WORD_4(2), 
        ELK_RX_SER_WORD_4(1) => ELK_RX_SER_WORD_4(1), 
        ELK_RX_SER_WORD_4(0) => ELK_RX_SER_WORD_4(0), 
        BIT_OS_SEL_1_0 => BIT_OS_SEL_1_0, BIT_OS_SEL_0(1) => 
        BIT_OS_SEL_0(1), BIT_OS_SEL_0(0) => BIT_OS_SEL_0(0), 
        BIT_OS_SEL_0_d0 => BIT_OS_SEL_0_d0, BIT_OS_SEL_6(2) => 
        BIT_OS_SEL_6(2), BIT_OS_SEL_6(1) => BIT_OS_SEL_6(1), 
        BIT_OS_SEL_7_0 => BIT_OS_SEL_7_0, CLK_40M_GL => 
        CLK_40M_GL, CCC_160M_FXD => CCC_160M_FXD, ELK_IN_R => 
        \ELK_IN_R\, ELK_IN_F => \ELK_IN_F\, 
        MASTER_DCB_POR_B_i_0_i => MASTER_DCB_POR_B_i_0_i, 
        CCC_160M_ADJ => CCC_160M_ADJ);
    
    U_ELK1_CMD_TX : SER320M_3_34_4
      port map(ELK_TX_DAT(7) => \ELK_TX_DAT[7]\, ELK_TX_DAT(6)
         => \ELK_TX_DAT[6]\, ELK_TX_DAT(5) => \ELK_TX_DAT[5]\, 
        ELK_TX_DAT(4) => \ELK_TX_DAT[4]\, ELK_TX_DAT(3) => 
        \ELK_TX_DAT[3]\, ELK_TX_DAT(2) => \ELK_TX_DAT[2]\, 
        ELK_TX_DAT(1) => \ELK_TX_DAT[1]\, ELK_TX_DAT(0) => 
        \ELK_TX_DAT[0]\, MASTER_SALT_POR_B_i_0_i_17 => 
        MASTER_SALT_POR_B_i_0_i_17, MASTER_SALT_POR_B_i_0_i_1 => 
        MASTER_SALT_POR_B_i_0_i_1, MASTER_SALT_POR_B_i_0_i_13 => 
        MASTER_SALT_POR_B_i_0_i_13, ELK_OUT_R_i_0 => 
        ELK_OUT_R_i_0, MASTER_SALT_POR_B_i_0_i_16 => 
        MASTER_SALT_POR_B_i_0_i_16, ELK_OUT_F_i_0 => 
        ELK_OUT_F_i_0, MASTER_SALT_POR_B_i_0_i_9 => 
        MASTER_SALT_POR_B_i_0_i_9, CLK_40M_GL => CLK_40M_GL, 
        MASTER_SALT_POR_B_i_0_i_4 => MASTER_SALT_POR_B_i_0_i_4, 
        CCC_160M_FXD => CCC_160M_FXD);
    
    U_DDR_ELK1 : DDR_BIDIR_LVDS_DUAL_CLK_4
      port map(DCB_SALT_SEL_c_i => DCB_SALT_SEL_c_i, ELK4_DAT_P
         => ELK4_DAT_P, ELK4_DAT_N => ELK4_DAT_N, ELK_OUT_R_i_0
         => ELK_OUT_R_i_0, ELK_OUT_F_i_0 => ELK_OUT_F_i_0, 
        CCC_160M_FXD => CCC_160M_FXD, CCC_160M_ADJ => 
        CCC_160M_ADJ, ELK_IN_DDR_F_i => ELK_IN_DDR_F_i, 
        ELK_IN_DDR_R_i => ELK_IN_DDR_R_i);
    
    ELK_IN_F : DFN1C0
      port map(D => ELK_IN_DDR_F_i, CLK => CCC_160M_ADJ, CLR => 
        DEV_RST_B_c, Q => \ELK_IN_F\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    U_ELK1_SERDAT_SOURCE : SYNC_DAT_SEL_4
      port map(ELK_TX_DAT(7) => \ELK_TX_DAT[7]\, ELK_TX_DAT(6)
         => \ELK_TX_DAT[6]\, ELK_TX_DAT(5) => \ELK_TX_DAT[5]\, 
        ELK_TX_DAT(4) => \ELK_TX_DAT[4]\, ELK_TX_DAT(3) => 
        \ELK_TX_DAT[3]\, ELK_TX_DAT(2) => \ELK_TX_DAT[2]\, 
        ELK_TX_DAT(1) => \ELK_TX_DAT[1]\, ELK_TX_DAT(0) => 
        \ELK_TX_DAT[0]\, PATT_ELK_DAT_4(7) => PATT_ELK_DAT_4(7), 
        PATT_ELK_DAT_4(6) => PATT_ELK_DAT_4(6), PATT_ELK_DAT_4(5)
         => PATT_ELK_DAT_4(5), PATT_ELK_DAT_4(4) => 
        PATT_ELK_DAT_4(4), PATT_ELK_DAT_4(3) => PATT_ELK_DAT_4(3), 
        PATT_ELK_DAT_4(2) => PATT_ELK_DAT_4(2), PATT_ELK_DAT_4(1)
         => PATT_ELK_DAT_4(1), PATT_ELK_DAT_4(0) => 
        PATT_ELK_DAT_4(0), OP_MODE_c_1_0 => OP_MODE_c_1_0, 
        MASTER_SALT_POR_B_i_0_i_16 => MASTER_SALT_POR_B_i_0_i_16, 
        CLK_40M_GL => CLK_40M_GL);
    
    ELK_IN_R : DFN1C0
      port map(D => ELK_IN_DDR_R_i, CLK => CCC_160M_ADJ, CLR => 
        DEV_RST_B_c, Q => \ELK_IN_R\);
    
    GND_i : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity DDR_BIDIR_LVDS_DUAL_CLK is

    port( DCB_SALT_SEL_c : in    std_logic;
          TFC_DAT_0P     : inout std_logic := 'Z';
          TFC_DAT_0N     : inout std_logic := 'Z';
          TFC_OUT_R      : in    std_logic;
          TFC_OUT_F      : in    std_logic;
          CCC_160M_FXD   : in    std_logic;
          CCC_160M_ADJ   : in    std_logic;
          TFC_IN_DDR_R   : out   std_logic;
          TFC_IN_DDR_F   : out   std_logic
        );

end DDR_BIDIR_LVDS_DUAL_CLK;

architecture DEF_ARCH of DDR_BIDIR_LVDS_DUAL_CLK is 

  component DDR_REG
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          QR  : out   std_logic;
          QF  : out   std_logic
        );
  end component;

  component DDR_OUT
    port( DR  : in    std_logic := 'U';
          DF  : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component BIBUF_LVDS
    port( PADP : inout   std_logic;
          PADN : inout   std_logic;
          D    : in    std_logic := 'U';
          E    : in    std_logic := 'U';
          Y    : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal DDR_BIDIR_LVDS_DUAL_CLK_GND, BIBUF_LVDS_0_Y, 
        DDR_OUT_0_Q, \VCC\ : std_logic;

begin 


    DDR_REG_0 : DDR_REG
      port map(D => BIBUF_LVDS_0_Y, CLK => CCC_160M_ADJ, CLR => 
        DDR_BIDIR_LVDS_DUAL_CLK_GND, QR => TFC_IN_DDR_R, QF => 
        TFC_IN_DDR_F);
    
    DDR_OUT_0 : DDR_OUT
      port map(DR => TFC_OUT_R, DF => TFC_OUT_F, CLK => 
        CCC_160M_FXD, CLR => DDR_BIDIR_LVDS_DUAL_CLK_GND, Q => 
        DDR_OUT_0_Q);
    
    BIBUF_LVDS_0 : BIBUF_LVDS
      port map(PADP => TFC_DAT_0P, PADN => TFC_DAT_0N, D => 
        DDR_OUT_0_Q, E => DCB_SALT_SEL_c, Y => BIBUF_LVDS_0_Y);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    GND_i : GND
      port map(Y => DDR_BIDIR_LVDS_DUAL_CLK_GND);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity tristate_buf is

    port( P_USB_MASTER_EN_c : in    std_logic;
          USB_RD_BI         : in    std_logic;
          USB_RD_B          : out   std_logic
        );

end tristate_buf;

architecture DEF_ARCH of tristate_buf is 

  component TRIBUFF_F_24U
    port( D   : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          PAD : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \GND\, \VCC\ : std_logic;

begin 


    \TRIBUFF_F_24U[0]\ : TRIBUFF_F_24U
      port map(D => USB_RD_BI, E => P_USB_MASTER_EN_c, PAD => 
        USB_RD_B);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    GND_i : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity REF_CLK_DIV_GEN is

    port( DEV_RST_B_c_1   : in    std_logic;
          Y               : in    std_logic;
          CLK40M_10NS_REF : out   std_logic
        );

end REF_CLK_DIV_GEN;

architecture DEF_ARCH of REF_CLK_DIV_GEN is 

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component XA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal un14_gen_40m_refcnt, \GEN_40M_REFCNT[1]_net_1\, 
        \GEN_40M_REFCNT[2]_net_1\, SUM1, 
        \GEN_40M_REFCNT[0]_net_1\, \N_GEN_40M_REFCNT[2]\, 
        \N_GEN_40M_REFCNT[0]\, \GND\, \VCC\ : std_logic;

begin 


    GEN_40M_REF : DFN1C0
      port map(D => un14_gen_40m_refcnt, CLK => Y, CLR => 
        DEV_RST_B_c_1, Q => CLK40M_10NS_REF);
    
    un2_n_gen_40m_refcnt_1_SUM1 : XOR2
      port map(A => \GEN_40M_REFCNT[0]_net_1\, B => 
        \GEN_40M_REFCNT[1]_net_1\, Y => SUM1);
    
    GEN_40M_REF_RNO : NOR2
      port map(A => \GEN_40M_REFCNT[1]_net_1\, B => 
        \GEN_40M_REFCNT[2]_net_1\, Y => un14_gen_40m_refcnt);
    
    \GEN_40M_REFCNT[0]\ : DFN1C0
      port map(D => \N_GEN_40M_REFCNT[0]\, CLK => Y, CLR => 
        DEV_RST_B_c_1, Q => \GEN_40M_REFCNT[0]_net_1\);
    
    \GEN_40M_REFCNT[2]\ : DFN1C0
      port map(D => \N_GEN_40M_REFCNT[2]\, CLK => Y, CLR => 
        DEV_RST_B_c_1, Q => \GEN_40M_REFCNT[2]_net_1\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \GEN_40M_REFCNT[1]\ : DFN1C0
      port map(D => SUM1, CLK => Y, CLR => DEV_RST_B_c_1, Q => 
        \GEN_40M_REFCNT[1]_net_1\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \GEN_40M_REFCNT_RNO[2]\ : XA1
      port map(A => \GEN_40M_REFCNT[0]_net_1\, B => 
        \GEN_40M_REFCNT[2]_net_1\, C => \GEN_40M_REFCNT[1]_net_1\, 
        Y => \N_GEN_40M_REFCNT[2]\);
    
    \GEN_40M_REFCNT_RNO[0]\ : OA1C
      port map(A => \GEN_40M_REFCNT[2]_net_1\, B => 
        \GEN_40M_REFCNT[1]_net_1\, C => \GEN_40M_REFCNT[0]_net_1\, 
        Y => \N_GEN_40M_REFCNT[0]\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SLAVE_DES320S_1_17_4 is

    port( ELK_RX_SER_WORD_6      : out   std_logic_vector(7 downto 0);
          BIT_OS_SEL_0           : in    std_logic;
          BIT_OS_SEL_6_0         : in    std_logic;
          BIT_OS_SEL_7_0         : in    std_logic;
          BIT_OS_SEL_5           : in    std_logic_vector(2 downto 1);
          CLK_40M_GL             : in    std_logic;
          CCC_160M_FXD           : in    std_logic;
          ELK_IN_R               : in    std_logic;
          ELK_IN_F               : in    std_logic;
          MASTER_DCB_POR_B_i_0_i : in    std_logic;
          CCC_160M_ADJ           : in    std_logic
        );

end SLAVE_DES320S_1_17_4;

architecture DEF_ARCH of SLAVE_DES320S_1_17_4 is 

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal N_17, \ARB_BYTE[0]_net_1\, \ARB_BYTE[4]_net_1\, N_18, 
        \ARB_BYTE[1]_net_1\, \ARB_BYTE[5]_net_1\, N_19, 
        \ARB_BYTE[2]_net_1\, \ARB_BYTE[6]_net_1\, N_20, 
        \ARB_BYTE[3]_net_1\, \ARB_BYTE[7]_net_1\, N_21, 
        \ARB_BYTE[8]_net_1\, N_22, \ARB_BYTE[9]_net_1\, N_23, 
        \ARB_BYTE[10]_net_1\, N_24, \ARB_BYTE[11]_net_1\, N_31, 
        \ARB_BYTE[12]_net_1\, N_32, \ARB_BYTE[13]_net_1\, N_33, 
        N_34, N_35, N_36, N_37, N_38, N_39, N_40, N_56, 
        \ARB_BYTE[14]_net_1\, N_64, \N_RECD_SER_WORD[0]\, 
        \N_RECD_SER_WORD[1]\, \N_RECD_SER_WORD[2]\, 
        \N_RECD_SER_WORD[3]\, \N_RECD_SER_WORD[4]\, 
        \N_RECD_SER_WORD[5]\, \N_RECD_SER_WORD[6]\, 
        \N_RECD_SER_WORD[7]\, \ADJ_SER_IN_F_0DEL\, 
        \ADJ_SER_IN_R_0DEL\, \ADJ_SER_IN_F_1DEL\, 
        \ADJ_SER_IN_R_1DEL\, \Q[0]_net_1\, \ADJ_Q[0]_net_1\, 
        \Q[1]_net_1\, \ADJ_Q[1]_net_1\, \Q[2]_net_1\, 
        \ADJ_Q[2]_net_1\, \Q[3]_net_1\, \ADJ_Q[3]_net_1\, 
        \Q[4]_net_1\, \ADJ_Q[4]_net_1\, \Q[5]_net_1\, 
        \ADJ_Q[5]_net_1\, \Q[6]_net_1\, \ADJ_Q[6]_net_1\, 
        \Q[7]_net_1\, \ADJ_Q[7]_net_1\, \Q[8]_net_1\, 
        \ADJ_Q[8]_net_1\, \Q[9]_net_1\, \ADJ_Q[9]_net_1\, 
        \Q[10]_net_1\, \ADJ_Q[10]_net_1\, \Q[11]_net_1\, 
        \ADJ_Q[11]_net_1\, \Q[12]_net_1\, \ADJ_Q[12]_net_1\, 
        \Q[13]_net_1\, \ADJ_Q[13]_net_1\, \Q[14]_net_1\, 
        \ADJ_Q[14]_net_1\, \ARB_WRD_40M_FIXED[0]_net_1\, 
        \ARB_WRD_40M_FIXED[1]_net_1\, 
        \ARB_WRD_40M_FIXED[2]_net_1\, 
        \ARB_WRD_40M_FIXED[3]_net_1\, 
        \ARB_WRD_40M_FIXED[4]_net_1\, 
        \ARB_WRD_40M_FIXED[5]_net_1\, 
        \ARB_WRD_40M_FIXED[6]_net_1\, 
        \ARB_WRD_40M_FIXED[7]_net_1\, 
        \ARB_WRD_40M_FIXED[8]_net_1\, 
        \ARB_WRD_40M_FIXED[9]_net_1\, 
        \ARB_WRD_40M_FIXED[10]_net_1\, 
        \ARB_WRD_40M_FIXED[11]_net_1\, 
        \ARB_WRD_40M_FIXED[12]_net_1\, 
        \ARB_WRD_40M_FIXED[13]_net_1\, 
        \ARB_WRD_40M_FIXED[14]_net_1\, \GND\, \VCC\ : std_logic;

begin 


    \RECD_SER_WORD_RNO[5]\ : MX2
      port map(A => N_38, B => N_39, S => BIT_OS_SEL_0, Y => 
        \N_RECD_SER_WORD[5]\);
    
    \ARB_WRD_40M_FIXED[9]\ : DFN1C0
      port map(D => \Q[9]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[9]_net_1\);
    
    \ADJ_Q[4]\ : DFN1C0
      port map(D => \ADJ_Q[2]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[4]_net_1\);
    
    \ARB_BYTE[6]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[6]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[6]_net_1\);
    
    ADJ_SER_IN_F_1DEL : DFN1C0
      port map(D => \ADJ_SER_IN_F_0DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_F_1DEL\);
    
    \ARB_BYTE[0]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[0]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[0]_net_1\);
    
    \Q[11]\ : DFN1C0
      port map(D => \ADJ_Q[11]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[11]_net_1\);
    
    \ADJ_Q[8]\ : DFN1C0
      port map(D => \ADJ_Q[6]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[8]_net_1\);
    
    \ARB_BYTE_RNI0H9K1[6]\ : MX2
      port map(A => N_23, B => N_31, S => BIT_OS_SEL_5(1), Y => 
        N_39);
    
    \ADJ_Q[6]\ : DFN1C0
      port map(D => \ADJ_Q[4]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[6]_net_1\);
    
    \ADJ_Q[12]\ : DFN1C0
      port map(D => \ADJ_Q[10]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[12]_net_1\);
    
    \RECD_SER_WORD_RNO_1[0]\ : MX2
      port map(A => \ARB_BYTE[0]_net_1\, B => \ARB_BYTE[4]_net_1\, 
        S => BIT_OS_SEL_5(2), Y => N_17);
    
    \Q[1]\ : DFN1C0
      port map(D => \ADJ_Q[1]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[1]_net_1\);
    
    \ARB_BYTE_RNIL9UF1[5]\ : MX2
      port map(A => N_22, B => N_24, S => BIT_OS_SEL_5(1), Y => 
        N_38);
    
    \ARB_BYTE[4]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[4]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[4]_net_1\);
    
    \ADJ_Q[2]\ : DFN1C0
      port map(D => \ADJ_Q[0]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[2]_net_1\);
    
    \RECD_SER_WORD_RNO_1[7]\ : MX2
      port map(A => \ARB_BYTE[10]_net_1\, B => 
        \ARB_BYTE[14]_net_1\, S => BIT_OS_SEL_7_0, Y => N_56);
    
    \RECD_SER_WORD[4]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[4]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_6(4));
    
    \Q[5]\ : DFN1C0
      port map(D => \ADJ_Q[5]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[5]_net_1\);
    
    \ADJ_Q[11]\ : DFN1C0
      port map(D => \ADJ_Q[9]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[11]_net_1\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \ADJ_Q[3]\ : DFN1C0
      port map(D => \ADJ_Q[1]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[3]_net_1\);
    
    \Q[10]\ : DFN1C0
      port map(D => \ADJ_Q[10]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[10]_net_1\);
    
    \ARB_WRD_40M_FIXED[6]\ : DFN1C0
      port map(D => \Q[6]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[6]_net_1\);
    
    \ARB_WRD_40M_FIXED[1]\ : DFN1C0
      port map(D => \Q[1]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[1]_net_1\);
    
    \RECD_SER_WORD[3]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[3]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_6(3));
    
    \ARB_BYTE_RNIBMUJ[4]\ : MX2
      port map(A => \ARB_BYTE[4]_net_1\, B => \ARB_BYTE[8]_net_1\, 
        S => BIT_OS_SEL_5(2), Y => N_21);
    
    \RECD_SER_WORD[0]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[0]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_6(0));
    
    \RECD_SER_WORD_RNO[3]\ : MX2
      port map(A => N_36, B => N_37, S => BIT_OS_SEL_0, Y => 
        \N_RECD_SER_WORD[3]\);
    
    \Q[0]\ : DFN1C0
      port map(D => \ADJ_Q[0]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[0]_net_1\);
    
    \RECD_SER_WORD_RNO_0[7]\ : MX2
      port map(A => N_31, B => N_56, S => BIT_OS_SEL_6_0, Y => 
        N_64);
    
    \Q[7]\ : DFN1C0
      port map(D => \ADJ_Q[7]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[7]_net_1\);
    
    \ARB_BYTE[14]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[14]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[14]_net_1\);
    
    \ARB_WRD_40M_FIXED[2]\ : DFN1C0
      port map(D => \Q[2]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[2]_net_1\);
    
    \ARB_WRD_40M_FIXED[14]\ : DFN1C0
      port map(D => \Q[14]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[14]_net_1\);
    
    \RECD_SER_WORD_RNO[2]\ : MX2
      port map(A => N_35, B => N_36, S => BIT_OS_SEL_0, Y => 
        \N_RECD_SER_WORD[2]\);
    
    \ARB_BYTE_RNI4L9K1[13]\ : MX2
      port map(A => N_24, B => N_32, S => BIT_OS_SEL_5(1), Y => 
        N_40);
    
    \ARB_BYTE[2]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[2]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[2]_net_1\);
    
    \ARB_BYTE_RNI2QIB1[2]\ : MX2
      port map(A => N_19, B => N_21, S => BIT_OS_SEL_5(1), Y => 
        N_35);
    
    \ADJ_Q[7]\ : DFN1C0
      port map(D => \ADJ_Q[5]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[7]_net_1\);
    
    \ARB_BYTE_RNIS3AO[13]\ : MX2
      port map(A => \ARB_BYTE[9]_net_1\, B => 
        \ARB_BYTE[13]_net_1\, S => BIT_OS_SEL_5(2), Y => N_32);
    
    \ARB_BYTE[8]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[8]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[8]_net_1\);
    
    \RECD_SER_WORD[5]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[5]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_6(5));
    
    \ARB_BYTE[12]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[12]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[12]_net_1\);
    
    \RECD_SER_WORD[1]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[1]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_6(1));
    
    \ARB_BYTE_RNIQ1AO[12]\ : MX2
      port map(A => \ARB_BYTE[8]_net_1\, B => 
        \ARB_BYTE[12]_net_1\, S => BIT_OS_SEL_5(2), Y => N_31);
    
    \ARB_BYTE_RNI5GUJ[1]\ : MX2
      port map(A => \ARB_BYTE[1]_net_1\, B => \ARB_BYTE[5]_net_1\, 
        S => BIT_OS_SEL_5(2), Y => N_18);
    
    \Q[3]\ : DFN1C0
      port map(D => \ADJ_Q[3]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[3]_net_1\);
    
    ADJ_SER_IN_F_0DEL : DFN1C0
      port map(D => ELK_IN_F, CLK => CCC_160M_ADJ, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_F_0DEL\);
    
    \RECD_SER_WORD_RNO[7]\ : MX2
      port map(A => N_40, B => N_64, S => BIT_OS_SEL_0, Y => 
        \N_RECD_SER_WORD[7]\);
    
    \RECD_SER_WORD_RNO[1]\ : MX2
      port map(A => N_34, B => N_35, S => BIT_OS_SEL_0, Y => 
        \N_RECD_SER_WORD[1]\);
    
    \ARB_WRD_40M_FIXED[4]\ : DFN1C0
      port map(D => \Q[4]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[4]_net_1\);
    
    \RECD_SER_WORD_RNO[0]\ : MX2
      port map(A => N_33, B => N_34, S => BIT_OS_SEL_0, Y => 
        \N_RECD_SER_WORD[0]\);
    
    \Q[6]\ : DFN1C0
      port map(D => \ADJ_Q[6]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[6]_net_1\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \ARB_WRD_40M_FIXED[8]\ : DFN1C0
      port map(D => \Q[8]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[8]_net_1\);
    
    \ARB_BYTE[11]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[11]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[11]_net_1\);
    
    \Q[9]\ : DFN1C0
      port map(D => \ADJ_Q[9]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[9]_net_1\);
    
    \ARB_BYTE_RNIOV9O[11]\ : MX2
      port map(A => \ARB_BYTE[7]_net_1\, B => 
        \ARB_BYTE[11]_net_1\, S => BIT_OS_SEL_5(2), Y => N_24);
    
    \Q[14]\ : DFN1C0
      port map(D => \ADJ_Q[14]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[14]_net_1\);
    
    ADJ_SER_IN_R_0DEL : DFN1C0
      port map(D => ELK_IN_R, CLK => CCC_160M_ADJ, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_R_0DEL\);
    
    \Q[13]\ : DFN1C0
      port map(D => \ADJ_Q[13]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[13]_net_1\);
    
    \ARB_BYTE[9]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[9]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[9]_net_1\);
    
    ADJ_SER_IN_R_1DEL : DFN1C0
      port map(D => \ADJ_SER_IN_R_0DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_R_1DEL\);
    
    \ARB_BYTE_RNI7IUJ[2]\ : MX2
      port map(A => \ARB_BYTE[2]_net_1\, B => \ARB_BYTE[6]_net_1\, 
        S => BIT_OS_SEL_5(2), Y => N_19);
    
    \ARB_BYTE[10]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[10]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[10]_net_1\);
    
    \ADJ_Q[9]\ : DFN1C0
      port map(D => \ADJ_Q[7]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[9]_net_1\);
    
    \RECD_SER_WORD[7]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[7]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_6(7));
    
    \ARB_WRD_40M_FIXED[5]\ : DFN1C0
      port map(D => \Q[5]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[5]_net_1\);
    
    \ARB_WRD_40M_FIXED[12]\ : DFN1C0
      port map(D => \Q[12]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[12]_net_1\);
    
    \ARB_WRD_40M_FIXED[11]\ : DFN1C0
      port map(D => \Q[11]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[11]_net_1\);
    
    \ARB_WRD_40M_FIXED[0]\ : DFN1C0
      port map(D => \Q[0]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[0]_net_1\);
    
    \ADJ_Q[10]\ : DFN1C0
      port map(D => \ADJ_Q[8]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[10]_net_1\);
    
    \Q[2]\ : DFN1C0
      port map(D => \ADJ_Q[2]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[2]_net_1\);
    
    \ADJ_Q[1]\ : DFN1C0
      port map(D => \ADJ_SER_IN_F_1DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[1]_net_1\);
    
    \RECD_SER_WORD[6]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[6]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_6(6));
    
    \ARB_BYTE_RNI6UIB1[3]\ : MX2
      port map(A => N_20, B => N_22, S => BIT_OS_SEL_5(1), Y => 
        N_36);
    
    \RECD_SER_WORD[2]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[2]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_6(2));
    
    \ARB_BYTE_RNIULIB1[1]\ : MX2
      port map(A => N_18, B => N_20, S => BIT_OS_SEL_5(1), Y => 
        N_34);
    
    \ADJ_Q[13]\ : DFN1C0
      port map(D => \ADJ_Q[11]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[13]_net_1\);
    
    \ARB_BYTE_RNIDOUJ[5]\ : MX2
      port map(A => \ARB_BYTE[5]_net_1\, B => \ARB_BYTE[9]_net_1\, 
        S => BIT_OS_SEL_5(2), Y => N_22);
    
    \Q[8]\ : DFN1C0
      port map(D => \ADJ_Q[8]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[8]_net_1\);
    
    \ARB_BYTE[5]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[5]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[5]_net_1\);
    
    \ARB_BYTE_RNIMT9O[6]\ : MX2
      port map(A => \ARB_BYTE[6]_net_1\, B => 
        \ARB_BYTE[10]_net_1\, S => BIT_OS_SEL_5(2), Y => N_23);
    
    \ADJ_Q[14]\ : DFN1C0
      port map(D => \ADJ_Q[12]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[14]_net_1\);
    
    \RECD_SER_WORD_RNO[4]\ : MX2
      port map(A => N_37, B => N_38, S => BIT_OS_SEL_0, Y => 
        \N_RECD_SER_WORD[4]\);
    
    \Q[12]\ : DFN1C0
      port map(D => \ADJ_Q[12]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[12]_net_1\);
    
    \ARB_BYTE_RNI9KUJ[3]\ : MX2
      port map(A => \ARB_BYTE[3]_net_1\, B => \ARB_BYTE[7]_net_1\, 
        S => BIT_OS_SEL_5(2), Y => N_20);
    
    \ARB_BYTE[13]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[13]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[13]_net_1\);
    
    \ARB_WRD_40M_FIXED[3]\ : DFN1C0
      port map(D => \Q[3]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[3]_net_1\);
    
    \ARB_BYTE[7]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[7]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[7]_net_1\);
    
    \RECD_SER_WORD_RNO_0[0]\ : MX2
      port map(A => N_17, B => N_19, S => BIT_OS_SEL_5(1), Y => 
        N_33);
    
    \Q[4]\ : DFN1C0
      port map(D => \ADJ_Q[4]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[4]_net_1\);
    
    \ARB_WRD_40M_FIXED[7]\ : DFN1C0
      port map(D => \Q[7]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[7]_net_1\);
    
    \RECD_SER_WORD_RNO[6]\ : MX2
      port map(A => N_39, B => N_40, S => BIT_OS_SEL_0, Y => 
        \N_RECD_SER_WORD[6]\);
    
    \ARB_BYTE_RNIH5UF1[4]\ : MX2
      port map(A => N_21, B => N_23, S => BIT_OS_SEL_5(1), Y => 
        N_37);
    
    \ARB_BYTE[3]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[3]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[3]_net_1\);
    
    \ADJ_Q[5]\ : DFN1C0
      port map(D => \ADJ_Q[3]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[5]_net_1\);
    
    \ARB_BYTE[1]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[1]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[1]_net_1\);
    
    \ARB_WRD_40M_FIXED[13]\ : DFN1C0
      port map(D => \Q[13]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[13]_net_1\);
    
    \ADJ_Q[0]\ : DFN1C0
      port map(D => \ADJ_SER_IN_R_1DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[0]_net_1\);
    
    \ARB_WRD_40M_FIXED[10]\ : DFN1C0
      port map(D => \Q[10]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[10]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SER320M_3_34_6 is

    port( ELK_TX_DAT                 : in    std_logic_vector(7 downto 0);
          MASTER_SALT_POR_B_i_0_i_6  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_9  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_3  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_12 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_16 : in    std_logic;
          ELK_OUT_R                  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_1  : in    std_logic;
          ELK_OUT_F                  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_10 : in    std_logic;
          CCC_160M_FXD               : in    std_logic;
          CLK_40M_GL                 : in    std_logic
        );

end SER320M_3_34_6;

architecture DEF_ARCH of SER320M_3_34_6 is 

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \N_SER_CMD_WORD_R[0]\, \START_RISE\, 
        \N_SER_CMD_WORD_F[0]\, \N_SER_CMD_WORD_R[3]\, 
        \SER_CMD_WORD_R[2]_net_1\, \N_SER_CMD_WORD_R[2]\, 
        \SER_CMD_WORD_R[1]_net_1\, \N_SER_CMD_WORD_R[1]\, 
        \SER_CMD_WORD_R[0]_net_1\, \N_SER_CMD_WORD_F[3]\, 
        \SER_CMD_WORD_F[2]_net_1\, \N_SER_CMD_WORD_F[2]\, 
        \SER_CMD_WORD_F[1]_net_1\, \N_SER_CMD_WORD_F[1]\, 
        \SER_CMD_WORD_F[0]_net_1\, N_START_RISE, 
        \CLK40M_GEN_DEL0\, \SER_OUT_FI\, \SER_OUT_RI\, 
        \SER_CMD_WORD_F[3]_net_1\, \SER_CMD_WORD_R[3]_net_1\, 
        \GND\, \VCC\ : std_logic;

begin 


    SER_OUT_FI : DFN1C0
      port map(D => \SER_CMD_WORD_F[3]_net_1\, CLK => 
        CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_3, Q => 
        \SER_OUT_FI\);
    
    \SER_CMD_WORD_F[3]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[3]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_9, Q => 
        \SER_CMD_WORD_F[3]_net_1\);
    
    \SER_CMD_WORD_R[1]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[1]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_6, Q => 
        \SER_CMD_WORD_R[1]_net_1\);
    
    \SER_CMD_WORD_R[2]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[2]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_6, Q => 
        \SER_CMD_WORD_R[2]_net_1\);
    
    \SER_CMD_WORD_R_RNO[3]\ : MX2
      port map(A => \SER_CMD_WORD_R[2]_net_1\, B => ELK_TX_DAT(7), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_R[3]\);
    
    \SER_CMD_WORD_R_RNO[0]\ : NOR2B
      port map(A => \START_RISE\, B => ELK_TX_DAT(1), Y => 
        \N_SER_CMD_WORD_R[0]\);
    
    \SER_CMD_WORD_F[0]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[0]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_9, Q => 
        \SER_CMD_WORD_F[0]_net_1\);
    
    \SER_CMD_WORD_R_RNO[1]\ : MX2
      port map(A => \SER_CMD_WORD_R[0]_net_1\, B => ELK_TX_DAT(3), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_R[1]\);
    
    \SER_CMD_WORD_F_RNO[2]\ : MX2
      port map(A => \SER_CMD_WORD_F[1]_net_1\, B => ELK_TX_DAT(4), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_F[2]\);
    
    \SER_CMD_WORD_F_RNO[3]\ : MX2
      port map(A => \SER_CMD_WORD_F[2]_net_1\, B => ELK_TX_DAT(6), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_F[3]\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    CLK40M_GEN_DEL0 : DFN1C0
      port map(D => CLK_40M_GL, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_10, Q => \CLK40M_GEN_DEL0\);
    
    SER_OUT_RI : DFN1C0
      port map(D => \SER_CMD_WORD_R[3]_net_1\, CLK => 
        CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_3, Q => 
        \SER_OUT_RI\);
    
    \SER_CMD_WORD_F[2]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[2]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_9, Q => 
        \SER_CMD_WORD_F[2]_net_1\);
    
    \SER_CMD_WORD_F_RNO[1]\ : MX2
      port map(A => \SER_CMD_WORD_F[0]_net_1\, B => ELK_TX_DAT(2), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_F[1]\);
    
    \SER_CMD_WORD_R[0]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[0]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_6, Q => 
        \SER_CMD_WORD_R[0]_net_1\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    START_RISE : DFN1C0
      port map(D => N_START_RISE, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_12, Q => \START_RISE\);
    
    \SER_CMD_WORD_R[3]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[3]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_6, Q => 
        \SER_CMD_WORD_R[3]_net_1\);
    
    \SER_CMD_WORD_F_RNO[0]\ : NOR2B
      port map(A => \START_RISE\, B => ELK_TX_DAT(0), Y => 
        \N_SER_CMD_WORD_F[0]\);
    
    SER_OUT_RDEL : DFN1C0
      port map(D => \SER_OUT_RI\, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_16, Q => ELK_OUT_R);
    
    \SER_CMD_WORD_F[1]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[1]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_9, Q => 
        \SER_CMD_WORD_F[1]_net_1\);
    
    START_RISE_RNO : NOR2B
      port map(A => \CLK40M_GEN_DEL0\, B => CLK_40M_GL, Y => 
        N_START_RISE);
    
    \SER_CMD_WORD_R_RNO[2]\ : MX2
      port map(A => \SER_CMD_WORD_R[1]_net_1\, B => ELK_TX_DAT(5), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_R[2]\);
    
    SER_OUT_FDEL : DFN1C0
      port map(D => \SER_OUT_FI\, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_1, Q => ELK_OUT_F);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity DDR_BIDIR_LVDS_DUAL_CLK_6 is

    port( DCB_SALT_SEL_c_i : in    std_logic;
          ELK6_DAT_P       : inout std_logic := 'Z';
          ELK6_DAT_N       : inout std_logic := 'Z';
          ELK_OUT_R        : in    std_logic;
          ELK_OUT_F        : in    std_logic;
          CCC_160M_FXD     : in    std_logic;
          CCC_160M_ADJ     : in    std_logic;
          ELK_IN_DDR_R     : out   std_logic;
          ELK_IN_DDR_F     : out   std_logic
        );

end DDR_BIDIR_LVDS_DUAL_CLK_6;

architecture DEF_ARCH of DDR_BIDIR_LVDS_DUAL_CLK_6 is 

  component DDR_REG
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          QR  : out   std_logic;
          QF  : out   std_logic
        );
  end component;

  component DDR_OUT
    port( DR  : in    std_logic := 'U';
          DF  : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component BIBUF_LVDS
    port( PADP : inout   std_logic;
          PADN : inout   std_logic;
          D    : in    std_logic := 'U';
          E    : in    std_logic := 'U';
          Y    : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal DDR_BIDIR_LVDS_DUAL_CLK_6_GND, BIBUF_LVDS_0_Y, 
        DDR_OUT_0_Q, \VCC\ : std_logic;

begin 


    DDR_REG_0 : DDR_REG
      port map(D => BIBUF_LVDS_0_Y, CLK => CCC_160M_ADJ, CLR => 
        DDR_BIDIR_LVDS_DUAL_CLK_6_GND, QR => ELK_IN_DDR_R, QF => 
        ELK_IN_DDR_F);
    
    DDR_OUT_0 : DDR_OUT
      port map(DR => ELK_OUT_R, DF => ELK_OUT_F, CLK => 
        CCC_160M_FXD, CLR => DDR_BIDIR_LVDS_DUAL_CLK_6_GND, Q => 
        DDR_OUT_0_Q);
    
    BIBUF_LVDS_0 : BIBUF_LVDS
      port map(PADP => ELK6_DAT_P, PADN => ELK6_DAT_N, D => 
        DDR_OUT_0_Q, E => DCB_SALT_SEL_c_i, Y => BIBUF_LVDS_0_Y);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    GND_i : GND
      port map(Y => DDR_BIDIR_LVDS_DUAL_CLK_6_GND);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SYNC_DAT_SEL_6 is

    port( ELK_TX_DAT                : out   std_logic_vector(7 downto 0);
          PATT_ELK_DAT_6            : in    std_logic_vector(7 downto 0);
          OP_MODE_c_1_0             : in    std_logic;
          OP_MODE_c_0_0             : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_2 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_1 : in    std_logic;
          CLK_40M_GL                : in    std_logic
        );

end SYNC_DAT_SEL_6;

architecture DEF_ARCH of SYNC_DAT_SEL_6 is 

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \N_SERDAT[0]\, \N_SERDAT[1]\, \N_SERDAT[2]\, 
        \N_SERDAT[3]\, \N_SERDAT[4]\, \N_SERDAT[5]\, 
        \N_SERDAT[6]\, \N_SERDAT[7]\, \GND\, \VCC\ : std_logic;

begin 


    \SERDAT_RNO[4]\ : NOR2A
      port map(A => PATT_ELK_DAT_6(4), B => OP_MODE_c_0_0, Y => 
        \N_SERDAT[4]\);
    
    \SERDAT_RNO[0]\ : NOR2A
      port map(A => PATT_ELK_DAT_6(0), B => OP_MODE_c_0_0, Y => 
        \N_SERDAT[0]\);
    
    \SERDAT[6]\ : DFN1C0
      port map(D => \N_SERDAT[6]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_2, Q => ELK_TX_DAT(6));
    
    \SERDAT[4]\ : DFN1C0
      port map(D => \N_SERDAT[4]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_1, Q => ELK_TX_DAT(4));
    
    \SERDAT_RNO[7]\ : OR2
      port map(A => PATT_ELK_DAT_6(7), B => OP_MODE_c_1_0, Y => 
        \N_SERDAT[7]\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \SERDAT_RNO[3]\ : OR2
      port map(A => PATT_ELK_DAT_6(3), B => OP_MODE_c_0_0, Y => 
        \N_SERDAT[3]\);
    
    \SERDAT_RNO[2]\ : OR2
      port map(A => PATT_ELK_DAT_6(2), B => OP_MODE_c_0_0, Y => 
        \N_SERDAT[2]\);
    
    \SERDAT[5]\ : DFN1C0
      port map(D => \N_SERDAT[5]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_1, Q => ELK_TX_DAT(5));
    
    \SERDAT[7]\ : DFN1C0
      port map(D => \N_SERDAT[7]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_2, Q => ELK_TX_DAT(7));
    
    GND_i : GND
      port map(Y => \GND\);
    
    \SERDAT_RNO[5]\ : NOR2A
      port map(A => PATT_ELK_DAT_6(5), B => OP_MODE_c_0_0, Y => 
        \N_SERDAT[5]\);
    
    \SERDAT[0]\ : DFN1C0
      port map(D => \N_SERDAT[0]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_1, Q => ELK_TX_DAT(0));
    
    \SERDAT_RNO[6]\ : NOR2A
      port map(A => PATT_ELK_DAT_6(6), B => OP_MODE_c_1_0, Y => 
        \N_SERDAT[6]\);
    
    \SERDAT[1]\ : DFN1C0
      port map(D => \N_SERDAT[1]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_1, Q => ELK_TX_DAT(1));
    
    \SERDAT_RNO[1]\ : OR2
      port map(A => PATT_ELK_DAT_6(1), B => OP_MODE_c_0_0, Y => 
        \N_SERDAT[1]\);
    
    \SERDAT[3]\ : DFN1C0
      port map(D => \N_SERDAT[3]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_1, Q => ELK_TX_DAT(3));
    
    \SERDAT[2]\ : DFN1C0
      port map(D => \N_SERDAT[2]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_1, Q => ELK_TX_DAT(2));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity ELINK_SLAVE_15_1 is

    port( BIT_OS_SEL_5               : in    std_logic_vector(2 downto 1);
          BIT_OS_SEL_7_0             : in    std_logic;
          BIT_OS_SEL_6_0             : in    std_logic;
          BIT_OS_SEL_0               : in    std_logic;
          ELK_RX_SER_WORD_6          : out   std_logic_vector(7 downto 0);
          OP_MODE_c_0_0              : in    std_logic;
          OP_MODE_c_1_0              : in    std_logic;
          PATT_ELK_DAT_6             : in    std_logic_vector(7 downto 0);
          MASTER_DCB_POR_B_i_0_i     : in    std_logic;
          ELK6_DAT_N                 : inout std_logic := 'Z';
          ELK6_DAT_P                 : inout std_logic := 'Z';
          DCB_SALT_SEL_c_i           : in    std_logic;
          CCC_160M_FXD               : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_10 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_16 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_12 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_3  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_9  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_6  : in    std_logic;
          CLK_40M_GL                 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_1  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_2  : in    std_logic;
          DEV_RST_B_c_1              : in    std_logic;
          CCC_160M_ADJ               : in    std_logic
        );

end ELINK_SLAVE_15_1;

architecture DEF_ARCH of ELINK_SLAVE_15_1 is 

  component SLAVE_DES320S_1_17_4
    port( ELK_RX_SER_WORD_6      : out   std_logic_vector(7 downto 0);
          BIT_OS_SEL_0           : in    std_logic := 'U';
          BIT_OS_SEL_6_0         : in    std_logic := 'U';
          BIT_OS_SEL_7_0         : in    std_logic := 'U';
          BIT_OS_SEL_5           : in    std_logic_vector(2 downto 1) := (others => 'U');
          CLK_40M_GL             : in    std_logic := 'U';
          CCC_160M_FXD           : in    std_logic := 'U';
          ELK_IN_R               : in    std_logic := 'U';
          ELK_IN_F               : in    std_logic := 'U';
          MASTER_DCB_POR_B_i_0_i : in    std_logic := 'U';
          CCC_160M_ADJ           : in    std_logic := 'U'
        );
  end component;

  component SER320M_3_34_6
    port( ELK_TX_DAT                 : in    std_logic_vector(7 downto 0) := (others => 'U');
          MASTER_SALT_POR_B_i_0_i_6  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_9  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_3  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_12 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_16 : in    std_logic := 'U';
          ELK_OUT_R                  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_1  : in    std_logic := 'U';
          ELK_OUT_F                  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_10 : in    std_logic := 'U';
          CCC_160M_FXD               : in    std_logic := 'U';
          CLK_40M_GL                 : in    std_logic := 'U'
        );
  end component;

  component DDR_BIDIR_LVDS_DUAL_CLK_6
    port( DCB_SALT_SEL_c_i : in    std_logic := 'U';
          ELK6_DAT_P       : inout   std_logic;
          ELK6_DAT_N       : inout   std_logic;
          ELK_OUT_R        : in    std_logic := 'U';
          ELK_OUT_F        : in    std_logic := 'U';
          CCC_160M_FXD     : in    std_logic := 'U';
          CCC_160M_ADJ     : in    std_logic := 'U';
          ELK_IN_DDR_R     : out   std_logic;
          ELK_IN_DDR_F     : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component SYNC_DAT_SEL_6
    port( ELK_TX_DAT                : out   std_logic_vector(7 downto 0);
          PATT_ELK_DAT_6            : in    std_logic_vector(7 downto 0) := (others => 'U');
          OP_MODE_c_1_0             : in    std_logic := 'U';
          OP_MODE_c_0_0             : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_2 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_1 : in    std_logic := 'U';
          CLK_40M_GL                : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \ELK_IN_F\, ELK_IN_DDR_F, \ELK_IN_R\, ELK_IN_DDR_R, 
        \ELK_TX_DAT[0]\, \ELK_TX_DAT[1]\, \ELK_TX_DAT[2]\, 
        \ELK_TX_DAT[3]\, \ELK_TX_DAT[4]\, \ELK_TX_DAT[5]\, 
        \ELK_TX_DAT[6]\, \ELK_TX_DAT[7]\, ELK_OUT_R, ELK_OUT_F, 
        \GND\, \VCC\ : std_logic;

    for all : SLAVE_DES320S_1_17_4
	Use entity work.SLAVE_DES320S_1_17_4(DEF_ARCH);
    for all : SER320M_3_34_6
	Use entity work.SER320M_3_34_6(DEF_ARCH);
    for all : DDR_BIDIR_LVDS_DUAL_CLK_6
	Use entity work.DDR_BIDIR_LVDS_DUAL_CLK_6(DEF_ARCH);
    for all : SYNC_DAT_SEL_6
	Use entity work.SYNC_DAT_SEL_6(DEF_ARCH);
begin 


    U_SLAVE_1ELK : SLAVE_DES320S_1_17_4
      port map(ELK_RX_SER_WORD_6(7) => ELK_RX_SER_WORD_6(7), 
        ELK_RX_SER_WORD_6(6) => ELK_RX_SER_WORD_6(6), 
        ELK_RX_SER_WORD_6(5) => ELK_RX_SER_WORD_6(5), 
        ELK_RX_SER_WORD_6(4) => ELK_RX_SER_WORD_6(4), 
        ELK_RX_SER_WORD_6(3) => ELK_RX_SER_WORD_6(3), 
        ELK_RX_SER_WORD_6(2) => ELK_RX_SER_WORD_6(2), 
        ELK_RX_SER_WORD_6(1) => ELK_RX_SER_WORD_6(1), 
        ELK_RX_SER_WORD_6(0) => ELK_RX_SER_WORD_6(0), 
        BIT_OS_SEL_0 => BIT_OS_SEL_0, BIT_OS_SEL_6_0 => 
        BIT_OS_SEL_6_0, BIT_OS_SEL_7_0 => BIT_OS_SEL_7_0, 
        BIT_OS_SEL_5(2) => BIT_OS_SEL_5(2), BIT_OS_SEL_5(1) => 
        BIT_OS_SEL_5(1), CLK_40M_GL => CLK_40M_GL, CCC_160M_FXD
         => CCC_160M_FXD, ELK_IN_R => \ELK_IN_R\, ELK_IN_F => 
        \ELK_IN_F\, MASTER_DCB_POR_B_i_0_i => 
        MASTER_DCB_POR_B_i_0_i, CCC_160M_ADJ => CCC_160M_ADJ);
    
    U_ELK1_CMD_TX : SER320M_3_34_6
      port map(ELK_TX_DAT(7) => \ELK_TX_DAT[7]\, ELK_TX_DAT(6)
         => \ELK_TX_DAT[6]\, ELK_TX_DAT(5) => \ELK_TX_DAT[5]\, 
        ELK_TX_DAT(4) => \ELK_TX_DAT[4]\, ELK_TX_DAT(3) => 
        \ELK_TX_DAT[3]\, ELK_TX_DAT(2) => \ELK_TX_DAT[2]\, 
        ELK_TX_DAT(1) => \ELK_TX_DAT[1]\, ELK_TX_DAT(0) => 
        \ELK_TX_DAT[0]\, MASTER_SALT_POR_B_i_0_i_6 => 
        MASTER_SALT_POR_B_i_0_i_6, MASTER_SALT_POR_B_i_0_i_9 => 
        MASTER_SALT_POR_B_i_0_i_9, MASTER_SALT_POR_B_i_0_i_3 => 
        MASTER_SALT_POR_B_i_0_i_3, MASTER_SALT_POR_B_i_0_i_12 => 
        MASTER_SALT_POR_B_i_0_i_12, MASTER_SALT_POR_B_i_0_i_16
         => MASTER_SALT_POR_B_i_0_i_16, ELK_OUT_R => ELK_OUT_R, 
        MASTER_SALT_POR_B_i_0_i_1 => MASTER_SALT_POR_B_i_0_i_1, 
        ELK_OUT_F => ELK_OUT_F, MASTER_SALT_POR_B_i_0_i_10 => 
        MASTER_SALT_POR_B_i_0_i_10, CCC_160M_FXD => CCC_160M_FXD, 
        CLK_40M_GL => CLK_40M_GL);
    
    U_DDR_ELK1 : DDR_BIDIR_LVDS_DUAL_CLK_6
      port map(DCB_SALT_SEL_c_i => DCB_SALT_SEL_c_i, ELK6_DAT_P
         => ELK6_DAT_P, ELK6_DAT_N => ELK6_DAT_N, ELK_OUT_R => 
        ELK_OUT_R, ELK_OUT_F => ELK_OUT_F, CCC_160M_FXD => 
        CCC_160M_FXD, CCC_160M_ADJ => CCC_160M_ADJ, ELK_IN_DDR_R
         => ELK_IN_DDR_R, ELK_IN_DDR_F => ELK_IN_DDR_F);
    
    ELK_IN_F : DFN1C0
      port map(D => ELK_IN_DDR_F, CLK => CCC_160M_ADJ, CLR => 
        DEV_RST_B_c_1, Q => \ELK_IN_F\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    U_ELK1_SERDAT_SOURCE : SYNC_DAT_SEL_6
      port map(ELK_TX_DAT(7) => \ELK_TX_DAT[7]\, ELK_TX_DAT(6)
         => \ELK_TX_DAT[6]\, ELK_TX_DAT(5) => \ELK_TX_DAT[5]\, 
        ELK_TX_DAT(4) => \ELK_TX_DAT[4]\, ELK_TX_DAT(3) => 
        \ELK_TX_DAT[3]\, ELK_TX_DAT(2) => \ELK_TX_DAT[2]\, 
        ELK_TX_DAT(1) => \ELK_TX_DAT[1]\, ELK_TX_DAT(0) => 
        \ELK_TX_DAT[0]\, PATT_ELK_DAT_6(7) => PATT_ELK_DAT_6(7), 
        PATT_ELK_DAT_6(6) => PATT_ELK_DAT_6(6), PATT_ELK_DAT_6(5)
         => PATT_ELK_DAT_6(5), PATT_ELK_DAT_6(4) => 
        PATT_ELK_DAT_6(4), PATT_ELK_DAT_6(3) => PATT_ELK_DAT_6(3), 
        PATT_ELK_DAT_6(2) => PATT_ELK_DAT_6(2), PATT_ELK_DAT_6(1)
         => PATT_ELK_DAT_6(1), PATT_ELK_DAT_6(0) => 
        PATT_ELK_DAT_6(0), OP_MODE_c_1_0 => OP_MODE_c_1_0, 
        OP_MODE_c_0_0 => OP_MODE_c_0_0, MASTER_SALT_POR_B_i_0_i_2
         => MASTER_SALT_POR_B_i_0_i_2, MASTER_SALT_POR_B_i_0_i_1
         => MASTER_SALT_POR_B_i_0_i_1, CLK_40M_GL => CLK_40M_GL);
    
    ELK_IN_R : DFN1C0
      port map(D => ELK_IN_DDR_R, CLK => CCC_160M_ADJ, CLR => 
        DEV_RST_B_c_1, Q => \ELK_IN_R\);
    
    GND_i : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity CCC_DYN_TRIPLE_160M is

    port( AUX_SUPDATE      : in    std_logic;
          AUX_SSHIFT       : in    std_logic;
          AUX_SDIN         : in    std_logic;
          AUX_MODE         : in    std_logic;
          CCC_RX_CLK_LOCK  : out   std_logic;
          CCC_160M_2ADJ_1  : out   std_logic;
          CCC_160M_1ADJ_1  : out   std_logic;
          CCC_160M_ADJ_1   : out   std_logic;
          CLK_40M_BUF_RECD : in    std_logic;
          CLK_40M_GL       : in    std_logic
        );

end CCC_DYN_TRIPLE_160M;

architecture DEF_ARCH of CCC_DYN_TRIPLE_160M is 

  component DYNCCC
    generic (VCOFREQUENCY:real := 0.0);

    port( CLKA      : in    std_logic := 'U';
          EXTFB     : in    std_logic := 'U';
          POWERDOWN : in    std_logic := 'U';
          GLA       : out   std_logic;
          LOCK      : out   std_logic;
          CLKB      : in    std_logic := 'U';
          GLB       : out   std_logic;
          YB        : out   std_logic;
          CLKC      : in    std_logic := 'U';
          GLC       : out   std_logic;
          YC        : out   std_logic;
          SDIN      : in    std_logic := 'U';
          SCLK      : in    std_logic := 'U';
          SSHIFT    : in    std_logic := 'U';
          SUPDATE   : in    std_logic := 'U';
          MODE      : in    std_logic := 'U';
          SDOUT     : out   std_logic;
          OADIV0    : in    std_logic := 'U';
          OADIV1    : in    std_logic := 'U';
          OADIV2    : in    std_logic := 'U';
          OADIV3    : in    std_logic := 'U';
          OADIV4    : in    std_logic := 'U';
          OAMUX0    : in    std_logic := 'U';
          OAMUX1    : in    std_logic := 'U';
          OAMUX2    : in    std_logic := 'U';
          DLYGLA0   : in    std_logic := 'U';
          DLYGLA1   : in    std_logic := 'U';
          DLYGLA2   : in    std_logic := 'U';
          DLYGLA3   : in    std_logic := 'U';
          DLYGLA4   : in    std_logic := 'U';
          OBDIV0    : in    std_logic := 'U';
          OBDIV1    : in    std_logic := 'U';
          OBDIV2    : in    std_logic := 'U';
          OBDIV3    : in    std_logic := 'U';
          OBDIV4    : in    std_logic := 'U';
          OBMUX0    : in    std_logic := 'U';
          OBMUX1    : in    std_logic := 'U';
          OBMUX2    : in    std_logic := 'U';
          DLYYB0    : in    std_logic := 'U';
          DLYYB1    : in    std_logic := 'U';
          DLYYB2    : in    std_logic := 'U';
          DLYYB3    : in    std_logic := 'U';
          DLYYB4    : in    std_logic := 'U';
          DLYGLB0   : in    std_logic := 'U';
          DLYGLB1   : in    std_logic := 'U';
          DLYGLB2   : in    std_logic := 'U';
          DLYGLB3   : in    std_logic := 'U';
          DLYGLB4   : in    std_logic := 'U';
          OCDIV0    : in    std_logic := 'U';
          OCDIV1    : in    std_logic := 'U';
          OCDIV2    : in    std_logic := 'U';
          OCDIV3    : in    std_logic := 'U';
          OCDIV4    : in    std_logic := 'U';
          OCMUX0    : in    std_logic := 'U';
          OCMUX1    : in    std_logic := 'U';
          OCMUX2    : in    std_logic := 'U';
          DLYYC0    : in    std_logic := 'U';
          DLYYC1    : in    std_logic := 'U';
          DLYYC2    : in    std_logic := 'U';
          DLYYC3    : in    std_logic := 'U';
          DLYYC4    : in    std_logic := 'U';
          DLYGLC0   : in    std_logic := 'U';
          DLYGLC1   : in    std_logic := 'U';
          DLYGLC2   : in    std_logic := 'U';
          DLYGLC3   : in    std_logic := 'U';
          DLYGLC4   : in    std_logic := 'U';
          FINDIV0   : in    std_logic := 'U';
          FINDIV1   : in    std_logic := 'U';
          FINDIV2   : in    std_logic := 'U';
          FINDIV3   : in    std_logic := 'U';
          FINDIV4   : in    std_logic := 'U';
          FINDIV5   : in    std_logic := 'U';
          FINDIV6   : in    std_logic := 'U';
          FBDIV0    : in    std_logic := 'U';
          FBDIV1    : in    std_logic := 'U';
          FBDIV2    : in    std_logic := 'U';
          FBDIV3    : in    std_logic := 'U';
          FBDIV4    : in    std_logic := 'U';
          FBDIV5    : in    std_logic := 'U';
          FBDIV6    : in    std_logic := 'U';
          FBDLY0    : in    std_logic := 'U';
          FBDLY1    : in    std_logic := 'U';
          FBDLY2    : in    std_logic := 'U';
          FBDLY3    : in    std_logic := 'U';
          FBDLY4    : in    std_logic := 'U';
          FBSEL0    : in    std_logic := 'U';
          FBSEL1    : in    std_logic := 'U';
          XDLYSEL   : in    std_logic := 'U';
          VCOSEL0   : in    std_logic := 'U';
          VCOSEL1   : in    std_logic := 'U';
          VCOSEL2   : in    std_logic := 'U'
        );
  end component;

  component PLLINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component INV
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal CLK_40M_GL_c_i, CLKAP, SDOUT, Core_YB, Core_YC, 
        CCC_DYN_TRIPLE_160M_GND, CCC_DYN_TRIPLE_160M_VCC
         : std_logic;

begin 


    Core : DYNCCC
      generic map(VCOFREQUENCY => 160.0)

      port map(CLKA => CLKAP, EXTFB => CCC_DYN_TRIPLE_160M_GND, 
        POWERDOWN => CCC_DYN_TRIPLE_160M_VCC, GLA => 
        CCC_160M_ADJ_1, LOCK => CCC_RX_CLK_LOCK, CLKB => 
        CCC_DYN_TRIPLE_160M_GND, GLB => CCC_160M_1ADJ_1, YB => 
        Core_YB, CLKC => CCC_DYN_TRIPLE_160M_GND, GLC => 
        CCC_160M_2ADJ_1, YC => Core_YC, SDIN => AUX_SDIN, SCLK
         => CLK_40M_GL_c_i, SSHIFT => AUX_SSHIFT, SUPDATE => 
        AUX_SUPDATE, MODE => AUX_MODE, SDOUT => SDOUT, OADIV0 => 
        CCC_DYN_TRIPLE_160M_GND, OADIV1 => 
        CCC_DYN_TRIPLE_160M_GND, OADIV2 => 
        CCC_DYN_TRIPLE_160M_GND, OADIV3 => 
        CCC_DYN_TRIPLE_160M_GND, OADIV4 => 
        CCC_DYN_TRIPLE_160M_GND, OAMUX0 => 
        CCC_DYN_TRIPLE_160M_GND, OAMUX1 => 
        CCC_DYN_TRIPLE_160M_GND, OAMUX2 => 
        CCC_DYN_TRIPLE_160M_VCC, DLYGLA0 => 
        CCC_DYN_TRIPLE_160M_GND, DLYGLA1 => 
        CCC_DYN_TRIPLE_160M_GND, DLYGLA2 => 
        CCC_DYN_TRIPLE_160M_GND, DLYGLA3 => 
        CCC_DYN_TRIPLE_160M_GND, DLYGLA4 => 
        CCC_DYN_TRIPLE_160M_GND, OBDIV0 => 
        CCC_DYN_TRIPLE_160M_GND, OBDIV1 => 
        CCC_DYN_TRIPLE_160M_GND, OBDIV2 => 
        CCC_DYN_TRIPLE_160M_GND, OBDIV3 => 
        CCC_DYN_TRIPLE_160M_GND, OBDIV4 => 
        CCC_DYN_TRIPLE_160M_GND, OBMUX0 => 
        CCC_DYN_TRIPLE_160M_GND, OBMUX1 => 
        CCC_DYN_TRIPLE_160M_GND, OBMUX2 => 
        CCC_DYN_TRIPLE_160M_VCC, DLYYB0 => 
        CCC_DYN_TRIPLE_160M_GND, DLYYB1 => 
        CCC_DYN_TRIPLE_160M_GND, DLYYB2 => 
        CCC_DYN_TRIPLE_160M_GND, DLYYB3 => 
        CCC_DYN_TRIPLE_160M_GND, DLYYB4 => 
        CCC_DYN_TRIPLE_160M_GND, DLYGLB0 => 
        CCC_DYN_TRIPLE_160M_GND, DLYGLB1 => 
        CCC_DYN_TRIPLE_160M_GND, DLYGLB2 => 
        CCC_DYN_TRIPLE_160M_GND, DLYGLB3 => 
        CCC_DYN_TRIPLE_160M_GND, DLYGLB4 => 
        CCC_DYN_TRIPLE_160M_GND, OCDIV0 => 
        CCC_DYN_TRIPLE_160M_GND, OCDIV1 => 
        CCC_DYN_TRIPLE_160M_GND, OCDIV2 => 
        CCC_DYN_TRIPLE_160M_GND, OCDIV3 => 
        CCC_DYN_TRIPLE_160M_GND, OCDIV4 => 
        CCC_DYN_TRIPLE_160M_GND, OCMUX0 => 
        CCC_DYN_TRIPLE_160M_GND, OCMUX1 => 
        CCC_DYN_TRIPLE_160M_GND, OCMUX2 => 
        CCC_DYN_TRIPLE_160M_VCC, DLYYC0 => 
        CCC_DYN_TRIPLE_160M_GND, DLYYC1 => 
        CCC_DYN_TRIPLE_160M_GND, DLYYC2 => 
        CCC_DYN_TRIPLE_160M_GND, DLYYC3 => 
        CCC_DYN_TRIPLE_160M_GND, DLYYC4 => 
        CCC_DYN_TRIPLE_160M_GND, DLYGLC0 => 
        CCC_DYN_TRIPLE_160M_GND, DLYGLC1 => 
        CCC_DYN_TRIPLE_160M_GND, DLYGLC2 => 
        CCC_DYN_TRIPLE_160M_GND, DLYGLC3 => 
        CCC_DYN_TRIPLE_160M_GND, DLYGLC4 => 
        CCC_DYN_TRIPLE_160M_GND, FINDIV0 => 
        CCC_DYN_TRIPLE_160M_VCC, FINDIV1 => 
        CCC_DYN_TRIPLE_160M_VCC, FINDIV2 => 
        CCC_DYN_TRIPLE_160M_VCC, FINDIV3 => 
        CCC_DYN_TRIPLE_160M_GND, FINDIV4 => 
        CCC_DYN_TRIPLE_160M_GND, FINDIV5 => 
        CCC_DYN_TRIPLE_160M_GND, FINDIV6 => 
        CCC_DYN_TRIPLE_160M_GND, FBDIV0 => 
        CCC_DYN_TRIPLE_160M_VCC, FBDIV1 => 
        CCC_DYN_TRIPLE_160M_VCC, FBDIV2 => 
        CCC_DYN_TRIPLE_160M_VCC, FBDIV3 => 
        CCC_DYN_TRIPLE_160M_VCC, FBDIV4 => 
        CCC_DYN_TRIPLE_160M_VCC, FBDIV5 => 
        CCC_DYN_TRIPLE_160M_GND, FBDIV6 => 
        CCC_DYN_TRIPLE_160M_GND, FBDLY0 => 
        CCC_DYN_TRIPLE_160M_VCC, FBDLY1 => 
        CCC_DYN_TRIPLE_160M_VCC, FBDLY2 => 
        CCC_DYN_TRIPLE_160M_VCC, FBDLY3 => 
        CCC_DYN_TRIPLE_160M_GND, FBDLY4 => 
        CCC_DYN_TRIPLE_160M_VCC, FBSEL0 => 
        CCC_DYN_TRIPLE_160M_GND, FBSEL1 => 
        CCC_DYN_TRIPLE_160M_VCC, XDLYSEL => 
        CCC_DYN_TRIPLE_160M_GND, VCOSEL0 => 
        CCC_DYN_TRIPLE_160M_GND, VCOSEL1 => 
        CCC_DYN_TRIPLE_160M_GND, VCOSEL2 => 
        CCC_DYN_TRIPLE_160M_VCC);
    
    pllint1 : PLLINT
      port map(A => CLK_40M_BUF_RECD, Y => CLKAP);
    
    VCC_i : VCC
      port map(Y => CCC_DYN_TRIPLE_160M_VCC);
    
    Core_RNO : INV
      port map(A => CLK_40M_GL, Y => CLK_40M_GL_c_i);
    
    GND_i : GND
      port map(Y => CCC_DYN_TRIPLE_160M_GND);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity GP_CCC_SCONFIG is

    port( PHASE_ADJ_160_L       : in    std_logic_vector(4 downto 0);
          P_MASTER_POR_B_c_34   : in    std_logic;
          P_MASTER_POR_B_c_19   : in    std_logic;
          P_MASTER_POR_B_c_18   : in    std_logic;
          P_MASTER_POR_B_c_33   : in    std_logic;
          P_MASTER_POR_B_c_31   : in    std_logic;
          P_MASTER_POR_B_c_22   : in    std_logic;
          AUX_SSHIFT            : out   std_logic;
          P_MASTER_POR_B_c_13   : in    std_logic;
          AUX_SUPDATE           : out   std_logic;
          P_MASTER_POR_B_c_25   : in    std_logic;
          P_MASTER_POR_B_c_6    : in    std_logic;
          AUX_SDIN              : out   std_logic;
          P_MASTER_POR_B_c_14   : in    std_logic;
          CCC2_CONFIG_TRIG_i_0  : in    std_logic;
          AUX_MODE              : out   std_logic;
          P_MASTER_POR_B_c_22_0 : in    std_logic;
          CLK_40M_GL            : in    std_logic
        );

end GP_CCC_SCONFIG;

architecture DEF_ARCH of GP_CCC_SCONFIG is 

  component MX2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E0C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component DFN1E1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component AX1E
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component AO1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component AOI1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \SHIFT_SM_0[4]_net_1\, \SHIFT_SM_ns[2]\, m6_0, 
        \BITCNT[7]_net_1\, \BITCNT[6]_net_1\, m15_1, 
        \BITCNT[5]_net_1\, m36_1, \SHIFT_SM[0]_net_1\, m23_e_0, 
        \SHIFT_SM_i_0[1]\, \SHIFT_SM[3]_net_1\, N_74_mux, 
        \BITCNT[4]_net_1\, \BITCNT[3]_net_1\, 
        \SHIFT_SM_RNIGM97[3]_net_1\, \SHIFT_SM[5]_net_1\, 
        N_106_mux, \BITCNT[1]_net_1\, \ALL81BITS[34]_net_1\, 
        \BITCNT[0]_net_1\, N_108_mux, \ALL81BITS[31]_net_1\, N_39, 
        N_75_mux, \BITCNT[2]_net_1\, N_86_mux, N_805, 
        N_SUPDATE_0_sqmuxa, \CCC1_MODE_RNO\, \AUX_MODE\, 
        N_CCC1_MODE_0_sqmuxa, N_5_0, N_2, N_36_0, N_8_0, N_89_mux, 
        \SHIFT_SM[6]_net_1\, N_18_0, \ALL81BITS[71]_net_1\, 
        N_19_0, \ALL81BITS[44]_net_1\, \SHIFT_SM[4]_net_1\, 
        N_26_0, N_27_0, \ALL81BITS[11]_net_1\, N_28_0, 
        \ALL81BITS[10]_net_1\, N_29_0, \ALL81BITS[9]_net_1\, 
        N_31_0, \ALL81BITS[7]_net_1\, N_825, \ALL81BITS[2]_net_1\, 
        N_46, i8_mux, N_826, N_827, \ALL81BITS[50]_net_1\, N_55, 
        i17_mux, N_829, N_59, N_60, N_63, N_61, N_62, N_830, 
        i5_mux, i7_mux, N_831, i23_mux, N_832, N_833, 
        \ALL81BITS[42]_net_1\, N_834, i2_mux, N_837, i11_mux, 
        i4_mux, N_838, N_839, N_840, i14_mux, N_841, 
        \ALL81BITS[0]_net_1\, \ALL81BITS[1]_net_1\, 
        \ALL81BITS[48]_net_1\, \ALL81BITS[49]_net_1\, 
        \ALL81BITS[8]_net_1\, \ALL81BITS[72]_net_1\, 
        \ALL81BITS[73]_net_1\, \ALL81BITS[40]_net_1\, 
        \ALL81BITS[41]_net_1\, \ALL81BITS[76]_net_1\, 
        \ALL81BITS[77]_net_1\, \ALL81BITS[78]_net_1\, 
        \ALL81BITS[79]_net_1\, \ALL81BITS[46]_net_1\, 
        \ALL81BITS[47]_net_1\, N_SDIN, N_SDIN_2, \SHIFT_SM_ns[4]\, 
        N_77_mux, \SHIFT_SM[2]_net_1\, N_17_0, N_20_0, N_21_0, 
        N_40, N_44, N_80_mux, BITCNT_n7, N_47, BITCNT_n6, 
        BITCNT_n5, N_52, BITCNT_n4, BITCNT_n3, BITCNT_n2, N_58, 
        \SHIFT_SM_RNO[5]_net_1\, \SHIFT_SM_RNO[0]_net_1\, N_636, 
        N_93_mux, BITCNT_n1, N_11_0, \ALL81BITS_RNO[41]_net_1\, 
        N_25_0, \SHIFT_SM_RNO[1]_net_1\, N_50, N_828, N_57, 
        \ALL81BITS[37]_net_1\, \ALL81BITS[39]_net_1\, N_64, N_65, 
        N_66, N_835, N_836, N_842, N_843, N_34_0, N_33_0, N_32_0, 
        N_30_0, N_24_0, N_23_0, N_22_0, \ALL81BITS_RNO[42]_net_1\, 
        \ALL81BITS_RNO[73]_net_1\, N_16_0, N_15_0, N_14_0, N_13_0, 
        \ALL81BITS_RNO[72]_net_1\, \GND\, \VCC\ : std_logic;

begin 

    AUX_MODE <= \AUX_MODE\;

    SDIN_RNO_19 : MX2A
      port map(A => N_830, B => N_831, S => \BITCNT[6]_net_1\, Y
         => N_832);
    
    \BITCNT[0]\ : DFN1E0C0
      port map(D => N_11_0, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_14, E => N_93_mux, Q => 
        \BITCNT[0]_net_1\);
    
    \ALL81BITS_RNO[44]\ : OR2
      port map(A => \ALL81BITS[44]_net_1\, B => 
        \SHIFT_SM[4]_net_1\, Y => N_19_0);
    
    SDIN_RNO_14 : NOR2A
      port map(A => N_46, B => \BITCNT[6]_net_1\, Y => N_826);
    
    \BITCNT_RNO[4]\ : NOR2
      port map(A => N_52, B => N_21_0, Y => BITCNT_n4);
    
    \ALL81BITS_RNO[76]\ : OR2
      port map(A => \ALL81BITS[76]_net_1\, B => 
        \SHIFT_SM[4]_net_1\, Y => N_16_0);
    
    \BITCNT_RNI3USJ[3]\ : NOR2B
      port map(A => \BITCNT[3]_net_1\, B => \BITCNT[4]_net_1\, Y
         => N_805);
    
    \BITCNT[7]\ : DFN1E0C0
      port map(D => BITCNT_n7, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_14, E => N_93_mux, Q => 
        \BITCNT[7]_net_1\);
    
    \SHIFT_SM[6]\ : DFN1P0
      port map(D => N_89_mux, CLK => CLK_40M_GL, PRE => 
        P_MASTER_POR_B_c_22_0, Q => \SHIFT_SM[6]_net_1\);
    
    \ALL81BITS_RNO[9]\ : OR2
      port map(A => \ALL81BITS[9]_net_1\, B => 
        \SHIFT_SM[4]_net_1\, Y => N_29_0);
    
    \SHIFT_SM_RNO_0[5]\ : NOR2A
      port map(A => \SHIFT_SM[5]_net_1\, B => N_86_mux, Y => N_58);
    
    \BITCNT_RNID5RT_1[2]\ : NOR2
      port map(A => \BITCNT[2]_net_1\, B => N_39, Y => N_36_0);
    
    \SHIFT_SM_RNIO1E43[0]\ : NOR3C
      port map(A => N_5_0, B => m6_0, C => \SHIFT_SM[0]_net_1\, Y
         => N_8_0);
    
    \SHIFT_SM_RNIIMQ1[1]\ : NOR2A
      port map(A => \SHIFT_SM_i_0[1]\, B => \SHIFT_SM[3]_net_1\, 
        Y => m23_e_0);
    
    \ALL81BITS_RNO[72]\ : OR2
      port map(A => \SHIFT_SM_0[4]_net_1\, B => 
        \ALL81BITS[72]_net_1\, Y => \ALL81BITS_RNO[72]_net_1\);
    
    \BITCNT[5]\ : DFN1E0C0
      port map(D => BITCNT_n5, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_14, E => N_93_mux, Q => 
        \BITCNT[5]_net_1\);
    
    \BITCNT_RNIMERT[3]\ : NOR3
      port map(A => \BITCNT[4]_net_1\, B => \BITCNT[3]_net_1\, C
         => \BITCNT[5]_net_1\, Y => N_74_mux);
    
    SDIN_RNO_33 : NOR2A
      port map(A => \ALL81BITS[42]_net_1\, B => \BITCNT[0]_net_1\, 
        Y => N_833);
    
    SDIN_RNO_23 : MX2A
      port map(A => i8_mux, B => N_825, S => \BITCNT[1]_net_1\, Y
         => N_46);
    
    SDIN_RNO_40 : MX2C
      port map(A => \ALL81BITS[10]_net_1\, B => 
        \ALL81BITS[11]_net_1\, S => \BITCNT[0]_net_1\, Y => 
        i7_mux);
    
    SDIN_RNO_18 : MX2C
      port map(A => N_61, B => N_62, S => \BITCNT[1]_net_1\, Y
         => N_63);
    
    \ALL81BITS[79]\ : DFN1C0
      port map(D => N_13_0, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_34, Q => \ALL81BITS[79]_net_1\);
    
    SUPDATE : DFN1E1C0
      port map(D => N_SUPDATE_0_sqmuxa, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_13, E => \SHIFT_SM_RNIGM97[3]_net_1\, 
        Q => AUX_SUPDATE);
    
    \BITCNT_RNO_0[4]\ : AX1E
      port map(A => N_40, B => \BITCNT[3]_net_1\, C => 
        \BITCNT[4]_net_1\, Y => N_52);
    
    \SHIFT_SM_RNIG8VK5[5]\ : MX2A
      port map(A => N_8_0, B => N_86_mux, S => 
        \SHIFT_SM[5]_net_1\, Y => N_17_0);
    
    \BITCNT_RNO_0[7]\ : NOR3C
      port map(A => \BITCNT[5]_net_1\, B => N_80_mux, C => 
        \BITCNT[6]_net_1\, Y => N_44);
    
    \SHIFT_SM_0_RNIVOT57[4]\ : OA1A
      port map(A => m23_e_0, B => \SHIFT_SM_0[4]_net_1\, C => 
        N_21_0, Y => N_93_mux);
    
    SDIN_RNO_9 : NOR2B
      port map(A => N_55, B => \BITCNT[5]_net_1\, Y => N_828);
    
    SDIN_RNO_35 : NOR2A
      port map(A => \ALL81BITS[44]_net_1\, B => \BITCNT[0]_net_1\, 
        Y => N_839);
    
    \BITCNT_RNI94TJ[7]\ : NOR2
      port map(A => \BITCNT[7]_net_1\, B => \BITCNT[6]_net_1\, Y
         => m6_0);
    
    SDIN_RNO_3 : MX2
      port map(A => N_836, B => N_842, S => \BITCNT[2]_net_1\, Y
         => N_843);
    
    SDIN_RNO_25 : NOR2A
      port map(A => \ALL81BITS[50]_net_1\, B => \BITCNT[0]_net_1\, 
        Y => N_827);
    
    \ALL81BITS_RNO[0]\ : OR2
      port map(A => \ALL81BITS[0]_net_1\, B => 
        \SHIFT_SM[4]_net_1\, Y => N_34_0);
    
    SDIN_RNO_2 : MX2
      port map(A => N_57, B => N_65, S => \BITCNT[2]_net_1\, Y
         => N_66);
    
    CCC1_MODE_RNO : OR2
      port map(A => \AUX_MODE\, B => N_CCC1_MODE_0_sqmuxa, Y => 
        \CCC1_MODE_RNO\);
    
    \BITCNT_RNO[3]\ : XA1B
      port map(A => \BITCNT[3]_net_1\, B => N_40, C => N_21_0, Y
         => BITCNT_n3);
    
    \SHIFT_SM[4]\ : DFN1C0
      port map(D => \SHIFT_SM_ns[2]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_22, Q => \SHIFT_SM[4]_net_1\);
    
    \ALL81BITS[34]\ : DFN1C0
      port map(D => N_25_0, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_33, Q => \ALL81BITS[34]_net_1\);
    
    \SHIFT_SM_RNO[5]\ : MX2B
      port map(A => N_58, B => CCC2_CONFIG_TRIG_i_0, S => 
        \SHIFT_SM[6]_net_1\, Y => \SHIFT_SM_RNO[5]_net_1\);
    
    SDIN_RNO_41 : MX2C
      port map(A => \ALL81BITS[72]_net_1\, B => 
        \ALL81BITS[73]_net_1\, S => \BITCNT[0]_net_1\, Y => 
        i23_mux);
    
    SDIN_RNO_42 : MX2C
      port map(A => \ALL81BITS[76]_net_1\, B => 
        \ALL81BITS[77]_net_1\, S => \BITCNT[0]_net_1\, Y => 
        i11_mux);
    
    \ALL81BITS_RNO[31]\ : OR2
      port map(A => \ALL81BITS[31]_net_1\, B => 
        \SHIFT_SM[4]_net_1\, Y => N_26_0);
    
    SDIN_RNO_39 : MX2C
      port map(A => \ALL81BITS[8]_net_1\, B => 
        \ALL81BITS[9]_net_1\, S => \BITCNT[0]_net_1\, Y => i5_mux);
    
    \SHIFT_SM_0[4]\ : DFN1C0
      port map(D => \SHIFT_SM_ns[2]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_22_0, Q => \SHIFT_SM_0[4]_net_1\);
    
    SDIN_RNO_29 : NOR2B
      port map(A => \ALL81BITS[39]_net_1\, B => \BITCNT[0]_net_1\, 
        Y => N_62);
    
    \ALL81BITS_RNO[79]\ : OR2
      port map(A => \ALL81BITS[79]_net_1\, B => 
        \SHIFT_SM_0[4]_net_1\, Y => N_13_0);
    
    \ALL81BITS[78]\ : DFN1C0
      port map(D => N_14_0, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_34, Q => \ALL81BITS[78]_net_1\);
    
    SDIN_RNO_34 : MX2
      port map(A => i11_mux, B => i4_mux, S => \BITCNT[1]_net_1\, 
        Y => N_837);
    
    \BITCNT_RNO_0[6]\ : AX1C
      port map(A => \BITCNT[5]_net_1\, B => N_80_mux, C => 
        \BITCNT[6]_net_1\, Y => N_47);
    
    SDIN_RNO_24 : MX2C
      port map(A => \ALL81BITS[48]_net_1\, B => 
        \ALL81BITS[49]_net_1\, S => \BITCNT[0]_net_1\, Y => 
        i17_mux);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \ALL81BITS_RNO[78]\ : OR2
      port map(A => \ALL81BITS[78]_net_1\, B => 
        \SHIFT_SM_0[4]_net_1\, Y => N_14_0);
    
    SDIN_RNO_17 : MX2C
      port map(A => N_829, B => N_59, S => \BITCNT[6]_net_1\, Y
         => N_60);
    
    \SHIFT_SM_RNO[6]\ : AO1
      port map(A => \SHIFT_SM[6]_net_1\, B => 
        CCC2_CONFIG_TRIG_i_0, C => N_CCC1_MODE_0_sqmuxa, Y => 
        N_89_mux);
    
    \ALL81BITS_RNO[77]\ : OR2
      port map(A => \ALL81BITS[77]_net_1\, B => 
        \SHIFT_SM_0[4]_net_1\, Y => N_15_0);
    
    \BITCNT_RNO[0]\ : NOR2
      port map(A => \BITCNT[0]_net_1\, B => N_21_0, Y => N_11_0);
    
    \ALL81BITS[72]\ : DFN1C0
      port map(D => \ALL81BITS_RNO[72]_net_1\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_33, Q => \ALL81BITS[72]_net_1\);
    
    SDIN_RNO_16 : MX2A
      port map(A => i17_mux, B => N_827, S => \BITCNT[1]_net_1\, 
        Y => N_55);
    
    \BITCNT_RNI50TJ[4]\ : NOR2
      port map(A => \BITCNT[4]_net_1\, B => \BITCNT[5]_net_1\, Y
         => N_2);
    
    \BITCNT[1]\ : DFN1E0C0
      port map(D => BITCNT_n1, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_14, E => N_93_mux, Q => 
        \BITCNT[1]_net_1\);
    
    \SHIFT_SM_RNIJ6KU6[2]\ : MX2
      port map(A => N_17_0, B => N_20_0, S => \SHIFT_SM[2]_net_1\, 
        Y => N_21_0);
    
    SDIN_RNO_38 : NOR2A
      port map(A => \ALL81BITS[2]_net_1\, B => \BITCNT[0]_net_1\, 
        Y => N_825);
    
    \ALL81BITS_RNO[42]\ : OR2
      port map(A => \ALL81BITS[42]_net_1\, B => 
        \SHIFT_SM[4]_net_1\, Y => \ALL81BITS_RNO[42]_net_1\);
    
    \SHIFT_SM_RNO[1]\ : OR2A
      port map(A => \SHIFT_SM[2]_net_1\, B => N_77_mux, Y => 
        \SHIFT_SM_RNO[1]_net_1\);
    
    SDIN_RNO_28 : NOR2B
      port map(A => \ALL81BITS[37]_net_1\, B => \BITCNT[0]_net_1\, 
        Y => N_61);
    
    \BITCNT_RNO[6]\ : NOR2A
      port map(A => N_47, B => N_21_0, Y => BITCNT_n6);
    
    \ALL81BITS[77]\ : DFN1C0
      port map(D => N_15_0, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_33, Q => \ALL81BITS[77]_net_1\);
    
    \SHIFT_SM_RNO[2]\ : AO1
      port map(A => N_77_mux, B => \SHIFT_SM[2]_net_1\, C => 
        \SHIFT_SM[3]_net_1\, Y => \SHIFT_SM_ns[4]\);
    
    SDIN_RNO_10 : MX2
      port map(A => N_60, B => N_63, S => \BITCNT[5]_net_1\, Y
         => N_64);
    
    SDIN_RNO : NOR2A
      port map(A => N_SDIN_2, B => \SHIFT_SM[6]_net_1\, Y => 
        N_SDIN);
    
    \ALL81BITS[71]\ : DFN1C0
      port map(D => N_18_0, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_33, Q => \ALL81BITS[71]_net_1\);
    
    \BITCNT_RNO[5]\ : XA1B
      port map(A => \BITCNT[5]_net_1\, B => N_80_mux, C => N_21_0, 
        Y => BITCNT_n5);
    
    \ALL81BITS[2]\ : DFN1C0
      port map(D => N_32_0, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_31, Q => \ALL81BITS[2]_net_1\);
    
    \BITCNT[4]\ : DFN1E0C0
      port map(D => BITCNT_n4, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_14, E => N_93_mux, Q => 
        \BITCNT[4]_net_1\);
    
    SDIN_RNO_8 : MX2
      port map(A => N_826, B => N_106_mux, S => \BITCNT[5]_net_1\, 
        Y => N_50);
    
    \ALL81BITS[44]\ : DFN1C0
      port map(D => N_19_0, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_33, Q => \ALL81BITS[44]_net_1\);
    
    \ALL81BITS[39]\ : DFN1C0
      port map(D => N_23_0, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_33, Q => \ALL81BITS[39]_net_1\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \ALL81BITS[73]\ : DFN1C0
      port map(D => \ALL81BITS_RNO[73]_net_1\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_33, Q => \ALL81BITS[73]_net_1\);
    
    \ALL81BITS_RNO[8]\ : OR2
      port map(A => \ALL81BITS[8]_net_1\, B => 
        \SHIFT_SM[4]_net_1\, Y => N_30_0);
    
    \BITCNT_RNID5RT_0[2]\ : NOR2B
      port map(A => N_39, B => \BITCNT[2]_net_1\, Y => N_40);
    
    SDIN_RNO_11 : MX2
      port map(A => N_832, B => N_834, S => \BITCNT[5]_net_1\, Y
         => N_835);
    
    SDIN_RNO_12 : MX2A
      port map(A => N_838, B => N_840, S => \BITCNT[5]_net_1\, Y
         => N_841);
    
    SDIN_RNO_0 : NOR2
      port map(A => \SHIFT_SM[6]_net_1\, B => \SHIFT_SM[2]_net_1\, 
        Y => N_636);
    
    \BITCNT_RNICOJF2[5]\ : NOR3C
      port map(A => m15_1, B => N_805, C => N_75_mux, Y => 
        N_86_mux);
    
    \ALL81BITS[76]\ : DFN1C0
      port map(D => N_16_0, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_33, Q => \ALL81BITS[76]_net_1\);
    
    \ALL81BITS[7]\ : DFN1C0
      port map(D => N_31_0, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_31, Q => \ALL81BITS[7]_net_1\);
    
    SDIN_RNO_37 : MX2C
      port map(A => \ALL81BITS[0]_net_1\, B => 
        \ALL81BITS[1]_net_1\, S => \BITCNT[0]_net_1\, Y => i8_mux);
    
    SDIN_RNO_27 : NOR2B
      port map(A => \ALL81BITS[71]_net_1\, B => N_39, Y => N_59);
    
    \ALL81BITS_RNO[34]\ : OR2
      port map(A => \ALL81BITS[34]_net_1\, B => 
        \SHIFT_SM_0[4]_net_1\, Y => N_25_0);
    
    \SHIFT_SM_RNIO1E43_0[0]\ : AOI1B
      port map(A => m6_0, B => N_5_0, C => \SHIFT_SM[0]_net_1\, Y
         => N_CCC1_MODE_0_sqmuxa);
    
    SDIN_RNO_36 : MX2C
      port map(A => \ALL81BITS[46]_net_1\, B => 
        \ALL81BITS[47]_net_1\, S => \BITCNT[0]_net_1\, Y => 
        i14_mux);
    
    SDIN_RNO_26 : NOR2B
      port map(A => \ALL81BITS[7]_net_1\, B => N_39, Y => N_829);
    
    \BITCNT[2]\ : DFN1E0C0
      port map(D => BITCNT_n2, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_14, E => N_93_mux, Q => 
        \BITCNT[2]_net_1\);
    
    \ALL81BITS_RNO[7]\ : OR2
      port map(A => \ALL81BITS[7]_net_1\, B => 
        \SHIFT_SM[4]_net_1\, Y => N_31_0);
    
    \ALL81BITS_RNO[71]\ : OR2
      port map(A => \ALL81BITS[71]_net_1\, B => 
        \SHIFT_SM_0[4]_net_1\, Y => N_18_0);
    
    \BITCNT_RNI8KJF2[2]\ : MX2
      port map(A => N_74_mux, B => N_2, S => N_36_0, Y => N_5_0);
    
    SDIN_RNO_30 : MX2
      port map(A => i5_mux, B => i7_mux, S => \BITCNT[1]_net_1\, 
        Y => N_830);
    
    SDIN_RNO_20 : MX2A
      port map(A => i2_mux, B => N_833, S => \BITCNT[1]_net_1\, Y
         => N_834);
    
    \ALL81BITS[49]\ : DFN1E1C0
      port map(D => PHASE_ADJ_160_L(3), CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_19, E => \SHIFT_SM_0[4]_net_1\, Q
         => \ALL81BITS[49]_net_1\);
    
    \ALL81BITS_RNO[11]\ : OR2
      port map(A => \ALL81BITS[11]_net_1\, B => 
        \SHIFT_SM[4]_net_1\, Y => N_27_0);
    
    \SHIFT_SM_RNO[0]\ : OR2A
      port map(A => \SHIFT_SM_i_0[1]\, B => N_8_0, Y => 
        \SHIFT_SM_RNO[0]_net_1\);
    
    \SHIFT_SM[3]\ : DFN1C0
      port map(D => \SHIFT_SM_0[4]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_22, Q => \SHIFT_SM[3]_net_1\);
    
    \ALL81BITS[0]\ : DFN1C0
      port map(D => N_34_0, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_31, Q => \ALL81BITS[0]_net_1\);
    
    \ALL81BITS[37]\ : DFN1C0
      port map(D => N_24_0, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_33, Q => \ALL81BITS[37]_net_1\);
    
    \BITCNT_RNID5RT[2]\ : NOR3A
      port map(A => \BITCNT[1]_net_1\, B => \BITCNT[2]_net_1\, C
         => \BITCNT[0]_net_1\, Y => N_75_mux);
    
    \ALL81BITS[31]\ : DFN1C0
      port map(D => N_26_0, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_33, Q => \ALL81BITS[31]_net_1\);
    
    \BITCNT_RNITNSJ[1]\ : NOR2B
      port map(A => \BITCNT[1]_net_1\, B => \BITCNT[0]_net_1\, Y
         => N_39);
    
    \ALL81BITS[8]\ : DFN1C0
      port map(D => N_30_0, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_31, Q => \ALL81BITS[8]_net_1\);
    
    SDIN_RNO_31 : NOR2
      port map(A => i23_mux, B => \BITCNT[1]_net_1\, Y => N_831);
    
    SDIN_RNO_32 : MX2C
      port map(A => \ALL81BITS[40]_net_1\, B => 
        \ALL81BITS[41]_net_1\, S => \BITCNT[0]_net_1\, Y => 
        i2_mux);
    
    SDIN_RNO_21 : NOR2A
      port map(A => \BITCNT[6]_net_1\, B => N_837, Y => N_838);
    
    SDIN_RNO_22 : MX2A
      port map(A => N_839, B => i14_mux, S => \BITCNT[1]_net_1\, 
        Y => N_840);
    
    \ALL81BITS[1]\ : DFN1C0
      port map(D => N_33_0, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_31, Q => \ALL81BITS[1]_net_1\);
    
    \SHIFT_SM_RNIO6HG2[5]\ : NOR2B
      port map(A => N_86_mux, B => \SHIFT_SM[5]_net_1\, Y => 
        \SHIFT_SM_ns[2]\);
    
    \BITCNT_RNIG3OH1[3]\ : NOR2B
      port map(A => N_805, B => N_40, Y => N_80_mux);
    
    SSHIFT : DFN1E1C0
      port map(D => \SHIFT_SM[2]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_13, E => \SHIFT_SM_RNIGM97[3]_net_1\, 
        Q => AUX_SSHIFT);
    
    SDIN_RNO_43 : MX2C
      port map(A => \ALL81BITS[78]_net_1\, B => 
        \ALL81BITS[79]_net_1\, S => \BITCNT[0]_net_1\, Y => 
        i4_mux);
    
    \ALL81BITS[48]\ : DFN1E1C0
      port map(D => PHASE_ADJ_160_L(2), CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_19, E => \SHIFT_SM_0[4]_net_1\, Q
         => \ALL81BITS[48]_net_1\);
    
    \SHIFT_SM_RNIQIN81[5]\ : NOR2
      port map(A => N_77_mux, B => \SHIFT_SM[5]_net_1\, Y => 
        N_20_0);
    
    \BITCNT_RNIE4Q71[7]\ : OA1C
      port map(A => \BITCNT[6]_net_1\, B => N_2, C => 
        \BITCNT[7]_net_1\, Y => N_77_mux);
    
    \SHIFT_SM[5]\ : DFN1C0
      port map(D => \SHIFT_SM_RNO[5]_net_1\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_22_0, Q => \SHIFT_SM[5]_net_1\);
    
    \BITCNT_RNO[2]\ : XA1B
      port map(A => \BITCNT[2]_net_1\, B => N_39, C => N_21_0, Y
         => BITCNT_n2);
    
    \BITCNT_RNO[1]\ : XA1B
      port map(A => \BITCNT[0]_net_1\, B => \BITCNT[1]_net_1\, C
         => N_21_0, Y => BITCNT_n1);
    
    \ALL81BITS[9]\ : DFN1C0
      port map(D => N_29_0, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_31, Q => \ALL81BITS[9]_net_1\);
    
    \ALL81BITS[42]\ : DFN1C0
      port map(D => \ALL81BITS_RNO[42]_net_1\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_33, Q => \ALL81BITS[42]_net_1\);
    
    \ALL81BITS_RNO[10]\ : OR2
      port map(A => \ALL81BITS[10]_net_1\, B => 
        \SHIFT_SM[4]_net_1\, Y => N_28_0);
    
    SDIN_RNO_6 : NOR2A
      port map(A => N_835, B => \BITCNT[4]_net_1\, Y => N_836);
    
    SDIN_RNO_4 : MX2
      port map(A => N_50, B => N_828, S => \BITCNT[4]_net_1\, Y
         => N_57);
    
    SDIN_RNO_5 : NOR2
      port map(A => N_64, B => \BITCNT[4]_net_1\, Y => N_65);
    
    \ALL81BITS_RNO[41]\ : OR2
      port map(A => \ALL81BITS[41]_net_1\, B => 
        \SHIFT_SM[4]_net_1\, Y => \ALL81BITS_RNO[41]_net_1\);
    
    \ALL81BITS[47]\ : DFN1E1C0
      port map(D => PHASE_ADJ_160_L(1), CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_18, E => \SHIFT_SM_0[4]_net_1\, Q
         => \ALL81BITS[47]_net_1\);
    
    CCC1_MODE : DFN1C0
      port map(D => \CCC1_MODE_RNO\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_25, Q => \AUX_MODE\);
    
    \ALL81BITS_RNO[2]\ : OR2
      port map(A => \ALL81BITS[2]_net_1\, B => 
        \SHIFT_SM[4]_net_1\, Y => N_32_0);
    
    \SHIFT_SM[1]\ : DFN1P0
      port map(D => \SHIFT_SM_RNO[1]_net_1\, CLK => CLK_40M_GL, 
        PRE => P_MASTER_POR_B_c_22, Q => \SHIFT_SM_i_0[1]\);
    
    \SHIFT_SM_RNIGM97[3]\ : NOR3
      port map(A => \SHIFT_SM[5]_net_1\, B => \SHIFT_SM[3]_net_1\, 
        C => \SHIFT_SM_0[4]_net_1\, Y => 
        \SHIFT_SM_RNIGM97[3]_net_1\);
    
    \ALL81BITS[50]\ : DFN1E1C0
      port map(D => PHASE_ADJ_160_L(4), CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_19, E => \SHIFT_SM_0[4]_net_1\, Q
         => \ALL81BITS[50]_net_1\);
    
    \ALL81BITS[41]\ : DFN1C0
      port map(D => \ALL81BITS_RNO[41]_net_1\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_33, Q => \ALL81BITS[41]_net_1\);
    
    \ALL81BITS[11]\ : DFN1C0
      port map(D => N_27_0, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_33, Q => \ALL81BITS[11]_net_1\);
    
    \ALL81BITS[40]\ : DFN1C0
      port map(D => N_22_0, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_33, Q => \ALL81BITS[40]_net_1\);
    
    \ALL81BITS[10]\ : DFN1C0
      port map(D => N_28_0, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_33, Q => \ALL81BITS[10]_net_1\);
    
    \SHIFT_SM[0]\ : DFN1C0
      port map(D => \SHIFT_SM_RNO[0]_net_1\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_22, Q => \SHIFT_SM[0]_net_1\);
    
    \ALL81BITS_RNO[1]\ : OR2
      port map(A => \ALL81BITS[1]_net_1\, B => 
        \SHIFT_SM[4]_net_1\, Y => N_33_0);
    
    SDIN_RNO_7 : MX2A
      port map(A => N_841, B => N_108_mux, S => \BITCNT[4]_net_1\, 
        Y => N_842);
    
    \BITCNT_RNO[7]\ : XA1B
      port map(A => \BITCNT[7]_net_1\, B => N_44, C => N_21_0, Y
         => BITCNT_n7);
    
    SUPDATE_RNO_0 : NOR3A
      port map(A => \SHIFT_SM[0]_net_1\, B => \BITCNT[7]_net_1\, 
        C => \BITCNT[6]_net_1\, Y => m36_1);
    
    \BITCNT_RNISKRT[5]\ : NOR2A
      port map(A => m6_0, B => \BITCNT[5]_net_1\, Y => m15_1);
    
    \BITCNT[3]\ : DFN1E0C0
      port map(D => BITCNT_n3, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_14, E => N_93_mux, Q => 
        \BITCNT[3]_net_1\);
    
    SUPDATE_RNO : NOR3C
      port map(A => N_74_mux, B => m36_1, C => N_75_mux, Y => 
        N_SUPDATE_0_sqmuxa);
    
    SDIN_RNO_13 : NOR3B
      port map(A => \ALL81BITS[31]_net_1\, B => N_39, C => 
        \BITCNT[5]_net_1\, Y => N_108_mux);
    
    \ALL81BITS[46]\ : DFN1E1C0
      port map(D => PHASE_ADJ_160_L(0), CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_18, E => \SHIFT_SM_0[4]_net_1\, Q
         => \ALL81BITS[46]_net_1\);
    
    \ALL81BITS_RNO[73]\ : OR2
      port map(A => \ALL81BITS[73]_net_1\, B => 
        \SHIFT_SM[4]_net_1\, Y => \ALL81BITS_RNO[73]_net_1\);
    
    \BITCNT[6]\ : DFN1E0C0
      port map(D => BITCNT_n6, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_14, E => N_93_mux, Q => 
        \BITCNT[6]_net_1\);
    
    \ALL81BITS_RNO[39]\ : OR2
      port map(A => \ALL81BITS[39]_net_1\, B => 
        \SHIFT_SM_0[4]_net_1\, Y => N_23_0);
    
    SDIN : DFN1E0C0
      port map(D => N_SDIN, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_6, E => N_636, Q => AUX_SDIN);
    
    \ALL81BITS_RNO[40]\ : OR2
      port map(A => \ALL81BITS[40]_net_1\, B => 
        \SHIFT_SM_0[4]_net_1\, Y => N_22_0);
    
    \ALL81BITS_RNO[37]\ : OR2
      port map(A => \ALL81BITS[37]_net_1\, B => 
        \SHIFT_SM[4]_net_1\, Y => N_24_0);
    
    SDIN_RNO_15 : NOR3B
      port map(A => \BITCNT[1]_net_1\, B => \ALL81BITS[34]_net_1\, 
        C => \BITCNT[0]_net_1\, Y => N_106_mux);
    
    SDIN_RNO_1 : MX2
      port map(A => N_66, B => N_843, S => \BITCNT[3]_net_1\, Y
         => N_SDIN_2);
    
    \SHIFT_SM[2]\ : DFN1C0
      port map(D => \SHIFT_SM_ns[4]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_22, Q => \SHIFT_SM[2]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity MASTER_DES320M is

    port( PHASE_ADJ_160_L       : out   std_logic_vector(4 downto 0);
          ELK_RX_SER_WORD_0     : out   std_logic_vector(7 downto 0);
          TFC_RX_SER_WORD       : out   std_logic_vector(7 downto 0);
          BIT_OS_SEL            : out   std_logic_vector(2 downto 0);
          OP_MODE_c_0           : in    std_logic;
          BIT_OS_SEL_0          : out   std_logic_vector(2 downto 0);
          BIT_OS_SEL_1          : out   std_logic_vector(2 downto 0);
          BIT_OS_SEL_2          : out   std_logic_vector(2 downto 0);
          BIT_OS_SEL_3          : out   std_logic_vector(2 downto 0);
          BIT_OS_SEL_4          : out   std_logic_vector(2 downto 0);
          BIT_OS_SEL_5          : out   std_logic_vector(2 downto 0);
          BIT_OS_SEL_6          : out   std_logic_vector(2 downto 1);
          BIT_OS_SEL_7_0        : out   std_logic;
          P_MASTER_POR_B_c      : in    std_logic;
          P_MASTER_POR_B_c_23   : in    std_logic;
          P_MASTER_POR_B_c_34   : in    std_logic;
          CCC_160M_FXD          : in    std_logic;
          P_MASTER_POR_B_c_33   : in    std_logic;
          P_MASTER_POR_B_c_32_0 : in    std_logic;
          P_MASTER_POR_B_c_34_0 : in    std_logic;
          P_MASTER_POR_B_c_28   : in    std_logic;
          P_MASTER_POR_B_c_30   : in    std_logic;
          P_MASTER_POR_B_c_29   : in    std_logic;
          P_MASTER_POR_B_c_8    : in    std_logic;
          P_MASTER_POR_B_c_19   : in    std_logic;
          P_MASTER_POR_B_c_18   : in    std_logic;
          P_MASTER_POR_B_c_20   : in    std_logic;
          P_MASTER_POR_B_c_1    : in    std_logic;
          P_MASTER_POR_B_c_17   : in    std_logic;
          P_MASTER_POR_B_c_13   : in    std_logic;
          P_MASTER_POR_B_c_10   : in    std_logic;
          P_MASTER_POR_B_c_27   : in    std_logic;
          ALIGN_ACTIVE          : out   std_logic;
          P_MASTER_POR_B_c_7    : in    std_logic;
          P_MASTER_POR_B_c_11   : in    std_logic;
          P_MASTER_POR_B_c_12   : in    std_logic;
          P_MASTER_POR_B_c_14   : in    std_logic;
          P_MASTER_POR_B_c_16   : in    std_logic;
          P_MASTER_POR_B_c_15   : in    std_logic;
          P_MASTER_POR_B_c_21   : in    std_logic;
          P_MASTER_POR_B_c_9    : in    std_logic;
          P_MASTER_POR_B_c_3    : in    std_logic;
          P_MASTER_POR_B_c_2    : in    std_logic;
          P_MASTER_POR_B_c_4    : in    std_logic;
          P_MASTER_POR_B_c_6    : in    std_logic;
          P_MASTER_POR_B_c_5    : in    std_logic;
          P_MASTER_POR_B_c_24   : in    std_logic;
          CCC2_CONFIG_TRIG_i_0  : out   std_logic;
          P_MASTER_POR_B_c_32   : in    std_logic;
          P_MASTER_POR_B_c_26   : in    std_logic;
          P_MASTER_POR_B_c_31_0 : in    std_logic;
          CCC_160M_ADJ          : in    std_logic;
          CCC_MAIN_LOCK         : in    std_logic;
          ALL_PLL_LOCK_c        : out   std_logic;
          ELK0_IN_F             : in    std_logic;
          TFC_IN_F              : in    std_logic;
          ELK0_IN_R             : in    std_logic;
          TFC_IN_R              : in    std_logic;
          DCB_SALT_SEL_c        : in    std_logic;
          ELK0_SYNC_DET_1       : out   std_logic;
          TFC_SYNC_DET_1        : out   std_logic;
          CCC_RX_CLK_LOCK       : in    std_logic;
          P_MASTER_POR_B_c_24_0 : in    std_logic;
          P_MASTER_POR_B_c_17_0 : in    std_logic;
          P_MASTER_POR_B_c_16_0 : in    std_logic;
          P_MASTER_POR_B_c_27_1 : in    std_logic;
          P_MASTER_POR_B_c_27_0 : in    std_logic;
          CLK_40M_GL            : in    std_logic
        );

end MASTER_DES320M;

architecture DEF_ARCH of MASTER_DES320M is 

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component NOR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OA1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E0C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component NOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component AO1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO13
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO16
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XNOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XNOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component DFN1E1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

    signal \BEST_BIT_OS_VAL[0]_net_1\, \BIT_OS_SEL_1[0]_net_1\, 
        \BEST_BIT_OS_VAL[1]_net_1\, \BIT_OS_SEL_1[1]_net_1\, 
        \BEST_BIT_OS_VAL[2]_net_1\, \BIT_OS_SEL_1[2]_net_1\, 
        \INDEX_CNT_4[0]_net_1\, \N_INDEX_CNT[0]\, N_5149, 
        \INDEX_CNT_3[0]_net_1\, \INDEX_CNT_2[0]_net_1\, 
        \INDEX_CNT_1[0]_net_1\, \INDEX_CNT_0[0]_net_1\, 
        \INDEX_CNT_0[2]_net_1\, \N_INDEX_CNT[2]\, 
        \INDEX_CNT_2[3]_net_1\, \N_INDEX_CNT[3]\, 
        \INDEX_CNT_1[3]_net_1\, \INDEX_CNT_0[3]_net_1\, 
        \CLKPHASE_0[1]_net_1\, \TUNE_CLKPHASE_RNI79F03[1]_net_1\, 
        \CLKPHASE_1[2]_net_1\, \TUNE_CLKPHASE_RNIDA643[2]_net_1\, 
        \CLKPHASE_0[2]_net_1\, \CLKPHASE_2[3]_net_1\, 
        \TUNE_CLKPHASE_RNILF0P2[3]_net_1\, \CLKPHASE_1[3]_net_1\, 
        \CLKPHASE_0[3]_net_1\, \CLKPHASE_5[4]_net_1\, 
        \TUNE_CLKPHASE_RNITINS2[4]_net_1\, \CLKPHASE_4[4]_net_1\, 
        \CLKPHASE_3[4]_net_1\, \CLKPHASE_2[4]_net_1\, 
        \CLKPHASE_1[4]_net_1\, \CLKPHASE_0[4]_net_1\, 
        \DES_SM_1[8]_net_1\, \DES_SM_ns[0]\, \DES_SM_0[8]_net_1\, 
        \DES_SM_4[6]_net_1\, N_MAX_CNT_0_sqmuxa, 
        \DES_SM_3[6]_net_1\, \DES_SM_2[6]_net_1\, 
        \DES_SM_1[6]_net_1\, \DES_SM_0[6]_net_1\, N_4530_2, 
        N_4530_1, N_4530_0, N_5666_0, N_BIT_OS_VAL_3126, N_84, 
        N_BIT_OS_VAL_3130, N_781_0, N_360, N_437, N_206_0, N_445, 
        N_209_0, N_BIT_OS_VAL_14_18_3_0_a2_1, N_717_0, N_782_0, 
        un1_DES_SM_1034_i_o2_1, N_754, un1_DES_SM_1034_i_o2_2, 
        \N_SEQCNTS_1_0[4]\, I_12, \N_SEQCNTS_1_0[3]\, I_9, 
        \N_SEQCNTS_1_0[2]\, I_7, \N_SEQCNTS_1_0[1]\, I_5, 
        \N_SEQCNTS_1_0[0]\, \un39_n_seqcnts[0]\, 
        \DWACT_ADD_CI_0_g_array_2[0]\, 
        \DWACT_ADD_CI_0_g_array_1[0]\, 
        \DWACT_ADD_CI_0_pog_array_1[0]\, \DWACT_ADD_CI_0_TMP[0]\, 
        \CLKPHASE[1]_net_1\, \DWACT_ADD_CI_0_g_array_12[0]\, 
        \CLKPHASE[2]_net_1\, N_4, \un39_n_seqcnts[1]\, N_2, 
        \un39_n_seqcnts[3]\, \DWACT_FINC_E[0]\, N_4_0, 
        \INDEX_CNT[1]_net_1\, \INDEX_CNT[0]_net_1\, N_2_0, 
        \INDEX_CNT[3]_net_1\, \DWACT_FINC_E_0[0]\, N_5792, 
        \DES_SM[8]_net_1\, \DES_SM[4]_net_1\, 
        un1_N_CCC_RESET_EN_0_sqmuxa, N_5784_i, N_128, N_5724, 
        n_best_clkphase14, un1_N_CCC_RESET_EN_0_sqmuxa_0_0_a3_0, 
        N_759, \CLKPHASE_RNIPQFPE1[0]_net_1\, 
        un1_DES_SM_1034_i_a2_0_1, N_427, N_758, 
        \DES_SM_ns_0_i_0_a3_0_1[6]\, \DES_SM_ns_0_i_0_a3_0_0[6]\, 
        \WAITCNT[13]_net_1\, un1_DES_SM_471_i_0_0_0_1, 
        un1_DES_SM_471_i_0_0_0_a3_0, N_116, 
        un1_DES_SM_471_i_0_0_0_0, N_5783, \DES_SM[0]_net_1\, 
        N_5730, un1_DES_SM_471_i_0_0_a3_0_0, 
        \DES_SM_ns_0_0_0_a2_4[0]\, \DES_SM_ns_0_0_0_a2_1[0]\, 
        \DES_SM_ns_0_0_0_a2_0[0]\, \DES_SM_ns_0_0_0_a2_2[0]\, 
        \WAITCNT[11]_net_1\, \WAITCNT[9]_net_1\, 
        \WAITCNT[10]_net_1\, \WAITCNT[12]_net_1\, 
        \WAITCNT[8]_net_1\, \un107_bit_os_val[0]\, 
        \un107_bit_os_val[1]\, N_761, un1_DES_SM_1034_i_a2_3_2, 
        un1_DES_SM_1034_i_a2_4_2, un1_DES_SM_1034_i_a2_4_0, 
        \un107_bit_os_val[3]\, \DES_SM[6]_net_1\, 
        N_BIT_OS_VAL_3110, N_BIT_OS_VAL_14_18_3_0_a2_0, 
        N_BIT_OS_VAL_312, N_BIT_OS_VAL_316, 
        \N_RECD_SER_WORD_iv_5[0]\, \ARB_BYTE_m[2]\, 
        \ARB_BYTE_m[0]\, \N_RECD_SER_WORD_iv_3[0]\, 
        \ARB_BYTE[1]_net_1\, n_recd_ser_word165, \ARB_BYTE_m[3]\, 
        \N_RECD_SER_WORD_iv_1[0]\, n_recd_ser_word170, 
        \ARB_BYTE[6]_net_1\, \ARB_BYTE_m[7]\, 
        \N_RECD_SER_WORD_iv_0[0]\, n_recd_ser_word168, 
        \ARB_BYTE[4]_net_1\, \ARB_BYTE_m[5]\, 
        \N_RECD_SER_WORD_iv_5[1]\, \ARB_BYTE_m_0[3]\, 
        \ARB_BYTE_m_0[1]\, \N_RECD_SER_WORD_iv_3[1]\, 
        \ARB_BYTE[2]_net_1\, \ARB_BYTE_m_0[4]\, 
        \N_RECD_SER_WORD_iv_1[1]\, \ARB_BYTE[7]_net_1\, 
        \ARB_BYTE_m[8]\, \N_RECD_SER_WORD_iv_0[1]\, 
        \ARB_BYTE[5]_net_1\, \ARB_BYTE_m_0[6]\, 
        \N_RECD_SER_WORD_iv_5[6]\, \ARB_BYTE_m_4[8]\, 
        \ARB_BYTE_m_5[6]\, \N_RECD_SER_WORD_iv_3[6]\, 
        \ARB_BYTE_m_3[9]\, \N_RECD_SER_WORD_iv_1[6]\, 
        \ARB_BYTE[12]_net_1\, \ARB_BYTE_m[13]\, 
        \N_RECD_SER_WORD_iv_0[6]\, \ARB_BYTE[10]_net_1\, 
        \ARB_BYTE_m_1[11]\, \N_RECD_SER_WORD_iv_5[3]\, 
        \ARB_BYTE_m_2[5]\, \ARB_BYTE_m_2[3]\, 
        \N_RECD_SER_WORD_iv_3[3]\, \ARB_BYTE_m_2[6]\, 
        \N_RECD_SER_WORD_iv_1[3]\, \ARB_BYTE[9]_net_1\, 
        \ARB_BYTE_m[10]\, \N_RECD_SER_WORD_iv_0[3]\, 
        \ARB_BYTE_m_1[8]\, \N_RECD_SER_WORD_iv_5[7]\, 
        \ARB_BYTE_m_4[9]\, \ARB_BYTE_m_6[7]\, 
        \N_RECD_SER_WORD_iv_3[7]\, \ARB_BYTE[8]_net_1\, 
        \ARB_BYTE_m_3[10]\, \N_RECD_SER_WORD_iv_1[7]\, 
        \ARB_BYTE[13]_net_1\, \ARB_BYTE_m[14]\, 
        \N_RECD_SER_WORD_iv_0[7]\, \ARB_BYTE[11]_net_1\, 
        \ARB_BYTE_m_1[12]\, \N_RECD_SER_WORD_iv_5[2]\, 
        \ARB_BYTE_m_1[4]\, \ARB_BYTE_m_1[2]\, 
        \N_RECD_SER_WORD_iv_3[2]\, \ARB_BYTE[3]_net_1\, 
        \ARB_BYTE_m_1[5]\, \N_RECD_SER_WORD_iv_1[2]\, 
        \ARB_BYTE_m[9]\, \N_RECD_SER_WORD_iv_0[2]\, 
        \ARB_BYTE_m_1[7]\, \N_RECD_SER_WORD_iv_5[5]\, 
        \ARB_BYTE_m_4[7]\, \ARB_BYTE_m_4[5]\, 
        \N_RECD_SER_WORD_iv_3[5]\, \ARB_BYTE_m_3[8]\, 
        \N_RECD_SER_WORD_iv_1[5]\, \ARB_BYTE_m[12]\, 
        \N_RECD_SER_WORD_iv_0[5]\, \ARB_BYTE_m_1[10]\, 
        \N_RECD_SER_WORD_iv_5[4]\, \ARB_BYTE_m_3[6]\, 
        \ARB_BYTE_m_3[4]\, \N_RECD_SER_WORD_iv_3[4]\, 
        \ARB_BYTE_m_3[7]\, \N_RECD_SER_WORD_iv_1[4]\, 
        \ARB_BYTE_m[11]\, \N_RECD_SER_WORD_iv_0[4]\, 
        \ARB_BYTE_m_1[9]\, BIT_OS_CNT_6_n7_i_0, \BIT_OS_CNT_6[6]\, 
        N_387, \BIT_OS_CNT_6[7]\, BIT_OS_CNT_6_n5_i_0, 
        \BIT_OS_CNT_6[4]\, N_378, \BIT_OS_CNT_6[5]\, 
        n_recd_ser_word166_0, \BIT_OS_SEL[1]_net_1\, 
        \BIT_OS_SEL[0]_net_1\, n_recd_ser_word169_0, 
        \BIT_OS_SEL[2]_net_1\, n_recd_ser_word171_0, 
        \BIT_OS_SEL[3]_net_1\, n_recd_ser_word170_0, DES_SM_tr7_0, 
        \CLKPHASE[0]_net_1\, DES_SM_tr5_0_a3_3, DES_SM_tr5_0_a3_1, 
        \MAX_CNT[6]_net_1\, \MAX_CNT[7]_net_1\, DES_SM_tr5_0_a3_2, 
        \MAX_CNT[5]_net_1\, \MAX_CNT[4]_net_1\, \DES_SM[7]_net_1\, 
        \MAX_CNT[8]_net_1\, DES_SM_tr8_i_o2_1, 
        \INDEX_CNT[4]_net_1\, \INDEX_CNT[2]_net_1\, 
        \DES_SM_ns_i_a2_i_a3_0[1]\, N_70, 
        \DES_SM_ns_i_a2_0_0_a3_0_1[5]\, \DES_SM_i_0[5]\, 
        \WAITCNT[0]_net_1\, N_123, BIT_OS_CNT_1lde_0_a3_2, 
        N_560_2, BIT_OS_CNT_1lde_0_a3_1, \ARB_BYTE[0]_net_1\, 
        N_776, BIT_OS_CNT_5lde_0_a3_2, N_563_2, 
        BIT_OS_CNT_5lde_0_a3_1, N_772, BIT_OS_CNT_2lde_0_a3_1, 
        BIT_OS_CNT_4lde_0_a3_1, BIT_OS_CNT_7lde_0_a3_1, N_562_3, 
        BIT_OS_CNT_7lde_0_a3_0, BIT_OS_CNT_0lde_0_a3_1, N_559_1, 
        BIT_OS_CNT_0lde_0_a3_0, N_771, BIT_OS_CNT_6lde_0_a3_1, 
        BIT_OS_CNT_6lde_0_a3_0, N_BIT_OS_VAL_316lto8_0_o3_2, 
        \BIT_OS_CNT_1[6]\, \BIT_OS_CNT_1[4]\, \BIT_OS_CNT_1[5]\, 
        N_BIT_OS_VAL_316lto8_0_o3_1, \BIT_OS_CNT_1[8]\, 
        \BIT_OS_CNT_1[7]\, N_BIT_OS_VAL_3118lto8_0_o3_2, 
        \BIT_OS_CNT_4[4]\, \BIT_OS_CNT_4[6]\, \BIT_OS_CNT_4[7]\, 
        N_BIT_OS_VAL_3118lto8_0_o3_1, \BIT_OS_CNT_4[8]\, 
        \BIT_OS_CNT_4[5]\, BIT_OS_CNT_3lde_0_a3_3, 
        BIT_OS_CNT_3lde_0_a3_1, BIT_OS_CNT_3lde_0_a3_0, 
        un1_DES_SM_471_i_0_a2_0_0_a2_9, 
        un1_DES_SM_471_i_0_a2_0_0_a2_6, 
        un1_DES_SM_471_i_0_a2_0_0_a2_8, \WAITCNT[5]_net_1\, 
        un1_DES_SM_471_i_0_a2_0_0_a2_4, 
        un1_DES_SM_471_i_0_a2_0_0_a2_7, \WAITCNT[1]_net_1\, 
        \WAITCNT[7]_net_1\, un1_DES_SM_471_i_0_a2_0_0_a2_2, 
        \WAITCNT[4]_net_1\, \WAITCNT[3]_net_1\, 
        \WAITCNT[2]_net_1\, \WAITCNT[6]_net_1\, 
        N_BIT_OS_VAL_3126lto8_0_o3_0, \BIT_OS_CNT_6[8]\, 
        N_BIT_OS_VAL_3110lto8_2, \BIT_OS_CNT_2[4]\, 
        \BIT_OS_CNT_2[8]\, \BIT_OS_CNT_2[5]\, 
        N_BIT_OS_VAL_3110lto8_1, \BIT_OS_CNT_2[7]\, 
        \BIT_OS_CNT_2[6]\, N_BIT_OS_VAL_3122lto8_0_o3_2, 
        \BIT_OS_CNT_5[4]\, \BIT_OS_CNT_5[5]\, \BIT_OS_CNT_5[8]\, 
        N_BIT_OS_VAL_3122lto8_0_o3_1, \BIT_OS_CNT_5[7]\, 
        \BIT_OS_CNT_5[6]\, N_BIT_OS_VAL_3130lto8_2, 
        \BIT_OS_CNT_7[4]\, \BIT_OS_CNT_7[8]\, \BIT_OS_CNT_7[5]\, 
        N_BIT_OS_VAL_3130lto8_1, \BIT_OS_CNT_7[7]\, 
        \BIT_OS_CNT_7[6]\, N_BIT_OS_VAL_3114lto8_2, 
        \BIT_OS_CNT_3[4]\, \BIT_OS_CNT_3[8]\, \BIT_OS_CNT_3[5]\, 
        N_BIT_OS_VAL_3114lto8_1, \BIT_OS_CNT_3[7]\, 
        \BIT_OS_CNT_3[6]\, ELK0_SYNC_DET_1_3, 
        \ELK_RX_SER_WORD_0[7]\, \RECD_SER_WORD[3]_net_1\, 
        \ELK_RX_SER_WORD_0[5]\, ELK0_SYNC_DET_1_2, 
        \ELK_RX_SER_WORD_0[0]\, \ELK_RX_SER_WORD_0[6]\, 
        ELK0_SYNC_DET_1_1, \RECD_SER_WORD[1]_net_1\, 
        \RECD_SER_WORD[2]_net_1\, \ELK_RX_SER_WORD_0[4]\, 
        DES_SM_tr2_i_a3_6, DES_SM_tr2_i_a3_4, DES_SM_tr2_i_a3_5, 
        \MAX_CNT[2]_net_1\, DES_SM_tr2_i_a3_2, \MAX_CNT[1]_net_1\, 
        \MAX_CNT[3]_net_1\, \MAX_CNT[0]_net_1\, 
        N_BIT_OS_VAL_312lto8_0_o3_2, \BIT_OS_CNT_0[5]\, 
        \BIT_OS_CNT_0[6]\, \BIT_OS_CNT_0[7]\, 
        N_BIT_OS_VAL_312lto8_0_o3_1, \BIT_OS_CNT_0[4]\, 
        \BIT_OS_CNT_0[8]\, N_CONFIG_ONCE_TRIG_i_a3_0, 
        \DES_SM[1]_net_1\, TFC_SYNC_DET_1_4, TFC_SYNC_DET_1_2, 
        \RECD_SER_WORD[4]_net_1\, \RECD_SER_WORD[0]_net_1\, 
        TFC_SYNC_DET_1_1, \RECD_SER_WORD[5]_net_1\, 
        \RECD_SER_WORD[6]_net_1\, n_recd_ser_word165_2, 
        n_recd_ser_word168_2, N_5072, N_5072_2, N_215, N_750, 
        \BIT_OS_CNT_0[2]\, \BIT_OS_CNT_0[1]\, \BIT_OS_CNT_0[3]\, 
        n_recd_ser_word164, \N_TUNE_CLKPHASE_2[2]\, 
        \BEST_SEQCNT[3]_net_1\, \BEST_CLKPHASE[2]_net_1\, N86, 
        \N_RECD_SER_WORD[7]\, \N_RECD_SER_WORD[6]\, 
        \N_RECD_SER_WORD[5]\, \N_RECD_SER_WORD[4]\, 
        \N_RECD_SER_WORD[3]\, \N_RECD_SER_WORD[2]\, 
        \N_RECD_SER_WORD[1]\, \N_RECD_SER_WORD[0]\, N_5626, N_409, 
        N_4530, N_511, N_5627, N_384, N_5628, N_376, N_5632, 
        N_419, N_75, N_79, N_81, N_524, N_83, N_430, N_525, N_85, 
        \BIT_OS_CNT_6[0]\, \BIT_OS_CNT_6[1]\, N_77, N_73, N_107, 
        N_435, N_5639, N_404, N_111, N_390, N_113, N_383, N_5640, 
        N_377, N_117, N_372, N_119, N_368, \N_TUNE_CLKPHASE_2[3]\, 
        \BEST_SEQCNT[4]_net_1\, \BEST_CLKPHASE[3]_net_1\, 
        I2_un1_CO1, N_35, N_420, N_5620, N_410, N_5621, N_501, 
        N_5622, N_382, N_5623, N_379, N_45, N_504, N_47, N_429, 
        N_505, N_5624, \BIT_OS_CNT_4[0]\, \BIT_OS_CNT_4[1]\, 
        N_BIT_OS_VAL_3118, N_363, N_375, N_103, un1_DES_SM_19, 
        N_5638, N_370, N_535, N_5637, N_5636, N_5635, N_385, 
        N_5634, N_388, N_5633, N_405, N_89, N_422, 
        N_BIT_OS_VAL_3114, N_BIT_OS_VAL_3114lt8, 
        \BIT_OS_CNT_3[2]\, \BIT_OS_CNT_3[3]\, \BIT_OS_CNT_3[1]\, 
        N_BIT_OS_VAL_3130lt8, \BIT_OS_CNT_7[2]\, 
        \BIT_OS_CNT_7[3]\, \BIT_OS_CNT_7[1]\, 
        \TFC_RX_SER_WORD[7]\, N_359, N_139, \BIT_OS_CNT_1[0]\, 
        \BIT_OS_CNT_1[1]\, N_137, N_428, N_555, N_135, N_380, 
        N_554, N_133, N_131, N_381, N_129, N_403, N_551, N_127, 
        N_125, N_436, \un107_bit_os_val[2]\, N_782, N_762, N_433, 
        N_121, \BIT_OS_CNT_0[0]\, N_209, N_781, N_365, N_354, 
        N_34, N_5775, N_4539, N_32, N_5776, N_41, N_5772, N_37, 
        N_5774, N_5859, \N_TUNE_CLKPHASE_2[1]\, 
        \BEST_SEQCNT[2]_net_1\, \BEST_CLKPHASE[1]_net_1\, 
        I0_un1_CO1, N_39, N_5773, N_43, N_5718, N_5779, N_5807, 
        N_5719, N_5777, N_BIT_OS_VAL_3122, N_760, N_5631, 
        \BIT_OS_CNT_5[0]\, \BIT_OS_CNT_5[1]\, N_5630, 
        \BIT_OS_CNT_5[2]\, N_367, N_5629, \BIT_OS_CNT_5[3]\, 
        N_373, N_5625, N_53, N_421, N_BIT_OS_VAL_3110lt8, 
        \BIT_OS_CNT_2[2]\, \BIT_OS_CNT_2[3]\, \BIT_OS_CNT_2[1]\, 
        N_1151_tz, BIT_OS_CNT_3_n2, BIT_OS_CNT_3_n2_tz, 
        \BIT_OS_CNT_3[0]\, BIT_OS_CNT_3_n3, BIT_OS_CNT_3_c2, 
        BIT_OS_CNT_3_n4, BIT_OS_CNT_3_n4_tz, BIT_OS_CNT_3_n5, 
        BIT_OS_CNT_3_c4, BIT_OS_CNT_3_n6, BIT_OS_CNT_3_c5, 
        BIT_OS_CNT_3_n7, BIT_OS_CNT_3_c6, BIT_OS_CNT_3_n8, 
        BIT_OS_CNT_3_432_0, BIT_OS_CNT_7_n2, BIT_OS_CNT_7_c1, 
        BIT_OS_CNT_7_n3, BIT_OS_CNT_7_c2, BIT_OS_CNT_7_n4, 
        BIT_OS_CNT_7_c3, BIT_OS_CNT_7_n5, BIT_OS_CNT_7_c4, 
        BIT_OS_CNT_7_n6, BIT_OS_CNT_7_c5, BIT_OS_CNT_7_n7, 
        BIT_OS_CNT_7_c6, BIT_OS_CNT_7_n8, BIT_OS_CNT_7_360_0, 
        \DES_SM_RNO[0]_net_1\, BIT_OS_CNT_2_n2, BIT_OS_CNT_2_c1, 
        BIT_OS_CNT_2_n3, BIT_OS_CNT_2_c2, BIT_OS_CNT_2_n4, 
        BIT_OS_CNT_2_c3, BIT_OS_CNT_2_n5, BIT_OS_CNT_2_c4, 
        BIT_OS_CNT_2_n6, BIT_OS_CNT_2_c5, BIT_OS_CNT_2_n7, 
        BIT_OS_CNT_2_c6, BIT_OS_CNT_2_n8, BIT_OS_CNT_2_260_0, N90, 
        \N_BEST_BIT_OS_VAL[0]\, \N_BEST_BIT_OS_VAL_3[0]\, 
        \N_BEST_BIT_OS_VAL[1]\, \N_BEST_BIT_OS_VAL_3[1]\, 
        \N_BEST_BIT_OS_VAL[2]\, \N_BEST_BIT_OS_VAL_3[2]\, 
        \N_BEST_BIT_OS_VAL[3]\, \N_BEST_BIT_OS_VAL_3[3]\, 
        \N_BEST_SEQCNT[0]\, \un6_n_best_seqcnt[0]\, 
        \N_BEST_SEQCNT[1]\, \un6_n_best_seqcnt[1]\, 
        \N_BEST_SEQCNT[2]\, \un6_n_best_seqcnt[2]\, 
        \N_BEST_SEQCNT[3]\, \un6_n_best_seqcnt[3]\, 
        \N_BEST_SEQCNT[4]\, \un6_n_best_seqcnt[4]\, 
        \N_SEQCNTS_1[0]\, \N_SEQCNTS_1[1]\, \N_SEQCNTS_1[2]\, 
        \N_SEQCNTS_1[3]\, \N_SEQCNTS_1[4]\, N_3599, 
        \BIT_OS_VAL_31[0]\, \BIT_OS_VAL_15[0]\, N_3600, 
        \BIT_OS_VAL_31[1]\, \BIT_OS_VAL_15[1]\, N_3601, 
        \BIT_OS_VAL_31[2]\, \BIT_OS_VAL_15[2]\, N_3603, 
        \BIT_OS_VAL_7[0]\, \BIT_OS_VAL_23[0]\, N_3604, 
        \BIT_OS_VAL_7[1]\, \BIT_OS_VAL_23[1]\, N_3605, 
        \BIT_OS_VAL_7[2]\, \BIT_OS_VAL_23[2]\, N_3607, N_3608, 
        N_3609, N_3611, \BIT_OS_VAL_3[0]\, \BIT_OS_VAL_19[0]\, 
        N_3612, \BIT_OS_VAL_3[1]\, \BIT_OS_VAL_19[1]\, N_3613, 
        \BIT_OS_VAL_3[2]\, \BIT_OS_VAL_19[2]\, N_3615, 
        \BIT_OS_VAL_11[0]\, \BIT_OS_VAL_27[0]\, N_3616, 
        \BIT_OS_VAL_11[1]\, \BIT_OS_VAL_27[1]\, N_3617, 
        \BIT_OS_VAL_11[2]\, \BIT_OS_VAL_27[2]\, N_3619, 
        \CLKPHASE[3]_net_1\, N_3620, N_3621, N_3623, N_3625, 
        N_3627, \BIT_OS_VAL_1[0]\, \BIT_OS_VAL_17[0]\, N_3628, 
        \BIT_OS_VAL_1[1]\, \BIT_OS_VAL_17[1]\, N_3629, 
        \BIT_OS_VAL_1[2]\, \BIT_OS_VAL_17[2]\, N_3630, 
        \BIT_OS_VAL_1[3]\, \BIT_OS_VAL_17[3]\, N_3631, 
        \BIT_OS_VAL_9[0]\, \BIT_OS_VAL_25[0]\, N_3632, 
        \BIT_OS_VAL_9[1]\, \BIT_OS_VAL_25[1]\, N_3633, 
        \BIT_OS_VAL_9[2]\, \BIT_OS_VAL_25[2]\, N_3634, 
        \BIT_OS_VAL_9[3]\, \BIT_OS_VAL_25[3]\, N_3635, N_3636, 
        N_3637, N_3639, \BIT_OS_VAL_5[0]\, \BIT_OS_VAL_21[0]\, 
        N_3640, \BIT_OS_VAL_5[1]\, \BIT_OS_VAL_21[1]\, N_3641, 
        \BIT_OS_VAL_5[2]\, \BIT_OS_VAL_21[2]\, N_3642, 
        \BIT_OS_VAL_5[3]\, \BIT_OS_VAL_21[3]\, N_3643, 
        \BIT_OS_VAL_13[0]\, \BIT_OS_VAL_29[0]\, N_3644, 
        \BIT_OS_VAL_13[1]\, \BIT_OS_VAL_29[1]\, N_3645, 
        \BIT_OS_VAL_13[2]\, \BIT_OS_VAL_29[2]\, 
        \CLKPHASE[4]_net_1\, N_3646, \BIT_OS_VAL_13[3]\, 
        \BIT_OS_VAL_29[3]\, N_3647, N_3648, N_3649, N_3651, 
        N_3653, N_3655, N_3657, N_3659, \BIT_OS_VAL_0[0]\, 
        \BIT_OS_VAL_16[0]\, N_3661, \BIT_OS_VAL_0[2]\, 
        \BIT_OS_VAL_16[2]\, N_3663, \BIT_OS_VAL_8[0]\, 
        \BIT_OS_VAL_24[0]\, N_3665, \BIT_OS_VAL_8[2]\, 
        \BIT_OS_VAL_24[2]\, N_3667, N_3669, N_3671, 
        \BIT_OS_VAL_4[0]\, \BIT_OS_VAL_20[0]\, N_3673, 
        \BIT_OS_VAL_4[2]\, \BIT_OS_VAL_20[2]\, N_3675, 
        \BIT_OS_VAL_12[0]\, \BIT_OS_VAL_28[0]\, N_3677, 
        \BIT_OS_VAL_12[2]\, \BIT_OS_VAL_28[2]\, N_3678, 
        \BIT_OS_VAL_12[3]\, \BIT_OS_VAL_28[3]\, N_3679, N_3681, 
        N_3683, N_3685, N_3687, \BIT_OS_VAL_2[0]\, 
        \BIT_OS_VAL_18[0]\, N_3688, \BIT_OS_VAL_2[1]\, 
        \BIT_OS_VAL_18[1]\, N_3689, \BIT_OS_VAL_2[2]\, 
        \BIT_OS_VAL_18[2]\, N_3690, \BIT_OS_VAL_2[3]\, 
        \BIT_OS_VAL_18[3]\, N_3691, \BIT_OS_VAL_10[0]\, 
        \BIT_OS_VAL_26[0]\, N_3692, \BIT_OS_VAL_10[1]\, 
        \BIT_OS_VAL_26[1]\, N_3693, \BIT_OS_VAL_10[2]\, 
        \BIT_OS_VAL_26[2]\, N_3694, \BIT_OS_VAL_10[3]\, 
        \BIT_OS_VAL_26[3]\, N_3695, N_3696, N_3697, N_3698, 
        N_3699, \BIT_OS_VAL_6[0]\, \BIT_OS_VAL_22[0]\, N_3700, 
        \BIT_OS_VAL_6[1]\, \BIT_OS_VAL_22[1]\, N_3701, 
        \BIT_OS_VAL_6[2]\, \BIT_OS_VAL_22[2]\, N_3702, 
        \BIT_OS_VAL_6[3]\, \BIT_OS_VAL_22[3]\, N_3703, 
        \BIT_OS_VAL_14[0]\, \BIT_OS_VAL_30[0]\, N_3704, 
        \BIT_OS_VAL_14[1]\, \BIT_OS_VAL_30[1]\, N_3705, 
        \BIT_OS_VAL_14[2]\, \BIT_OS_VAL_30[2]\, N_3706, 
        \BIT_OS_VAL_14[3]\, \BIT_OS_VAL_30[3]\, N_3707, N_3708, 
        N_3709, N_3710, N_3711, N_3712, N_3713, N_3714, N_3715, 
        N_3717, N_3723, \SEQCNTS_31[0]\, \SEQCNTS_15[0]\, N_3724, 
        \SEQCNTS_31[1]\, \SEQCNTS_15[1]\, N_3725, \SEQCNTS_31[2]\, 
        \SEQCNTS_15[2]\, N_3726, \SEQCNTS_31[3]\, \SEQCNTS_15[3]\, 
        N_3727, \SEQCNTS_31[4]\, \SEQCNTS_15[4]\, N_3728, 
        \SEQCNTS_7[0]\, \SEQCNTS_23[0]\, N_3729, \SEQCNTS_7[1]\, 
        \SEQCNTS_23[1]\, N_3730, \SEQCNTS_7[2]\, \SEQCNTS_23[2]\, 
        N_3731, \SEQCNTS_7[3]\, \SEQCNTS_23[3]\, N_3732, 
        \SEQCNTS_7[4]\, \SEQCNTS_23[4]\, N_3733, N_3734, N_3735, 
        N_3736, N_3737, N_3738, \SEQCNTS_3[0]\, \SEQCNTS_19[0]\, 
        N_3739, \SEQCNTS_3[1]\, \SEQCNTS_19[1]\, N_3740, 
        \SEQCNTS_3[2]\, \SEQCNTS_19[2]\, N_3741, \SEQCNTS_3[3]\, 
        \SEQCNTS_19[3]\, N_3742, \SEQCNTS_3[4]\, \SEQCNTS_19[4]\, 
        N_3743, \SEQCNTS_11[0]\, \SEQCNTS_27[0]\, N_3744, 
        \SEQCNTS_11[1]\, \SEQCNTS_27[1]\, N_3745, \SEQCNTS_11[2]\, 
        \SEQCNTS_27[2]\, N_3746, \SEQCNTS_11[3]\, \SEQCNTS_27[3]\, 
        N_3747, \SEQCNTS_11[4]\, \SEQCNTS_27[4]\, N_3748, N_3749, 
        N_3750, N_3751, N_3752, N_3753, N_3754, N_3755, N_3756, 
        N_3757, N_3758, \SEQCNTS_1[0]\, \SEQCNTS_17[0]\, N_3759, 
        \SEQCNTS_1[1]\, \SEQCNTS_17[1]\, N_3760, \SEQCNTS_1[2]\, 
        \SEQCNTS_17[2]\, N_3761, \SEQCNTS_1[3]\, \SEQCNTS_17[3]\, 
        N_3762, \SEQCNTS_1[4]\, \SEQCNTS_17[4]\, N_3763, 
        \SEQCNTS_9[0]\, \SEQCNTS_25[0]\, N_3764, \SEQCNTS_9[1]\, 
        \SEQCNTS_25[1]\, N_3765, \SEQCNTS_9[2]\, \SEQCNTS_25[2]\, 
        N_3766, \SEQCNTS_9[3]\, \SEQCNTS_25[3]\, N_3767, 
        \SEQCNTS_9[4]\, \SEQCNTS_25[4]\, N_3768, N_3769, N_3770, 
        N_3771, N_3772, N_3773, \SEQCNTS_5[0]\, \SEQCNTS_21[0]\, 
        N_3774, \SEQCNTS_5[1]\, \SEQCNTS_21[1]\, N_3775, 
        \SEQCNTS_5[2]\, \SEQCNTS_21[2]\, N_3776, \SEQCNTS_5[3]\, 
        \SEQCNTS_21[3]\, N_3777, \SEQCNTS_5[4]\, \SEQCNTS_21[4]\, 
        N_3778, \SEQCNTS_13[0]\, \SEQCNTS_29[0]\, N_3779, 
        \SEQCNTS_13[1]\, \SEQCNTS_29[1]\, N_3780, \SEQCNTS_13[2]\, 
        \SEQCNTS_29[2]\, N_3781, \SEQCNTS_13[3]\, \SEQCNTS_29[3]\, 
        N_3782, \SEQCNTS_13[4]\, \SEQCNTS_29[4]\, N_3783, N_3784, 
        N_3785, N_3786, N_3787, N_3788, N_3789, N_3790, N_3791, 
        N_3792, N_3793, N_3794, N_3795, N_3796, N_3797, N_3803, 
        \SEQCNTS_8[0]\, \SEQCNTS_24[0]\, N_3804, \SEQCNTS_8[1]\, 
        \SEQCNTS_24[1]\, N_3805, \SEQCNTS_8[2]\, \SEQCNTS_24[2]\, 
        N_3806, \SEQCNTS_8[3]\, \SEQCNTS_24[3]\, N_3807, 
        \SEQCNTS_8[4]\, \SEQCNTS_24[4]\, N_3808, N_3798, N_3809, 
        N_3799, N_3810, N_3800, N_3811, N_3801, N_3812, N_3802, 
        N_3813, \SEQCNTS_4[0]\, \SEQCNTS_20[0]\, N_3814, 
        \SEQCNTS_4[1]\, \SEQCNTS_20[1]\, N_3815, \SEQCNTS_4[2]\, 
        \SEQCNTS_20[2]\, N_3816, \SEQCNTS_4[3]\, \SEQCNTS_20[3]\, 
        N_3817, \SEQCNTS_4[4]\, \SEQCNTS_20[4]\, N_3818, 
        \SEQCNTS_12[0]\, \SEQCNTS_28[0]\, N_3819, \SEQCNTS_12[1]\, 
        \SEQCNTS_28[1]\, N_3820, \SEQCNTS_12[2]\, \SEQCNTS_28[2]\, 
        N_3821, \SEQCNTS_12[3]\, \SEQCNTS_28[3]\, N_3822, 
        \SEQCNTS_12[4]\, \SEQCNTS_28[4]\, N_3823, N_3824, N_3825, 
        N_3826, N_3827, N_3828, N_3829, N_3830, N_3831, N_3832, 
        N_3833, \SEQCNTS_2[0]\, \SEQCNTS_18[0]\, N_3834, 
        \SEQCNTS_2[1]\, \SEQCNTS_18[1]\, N_3835, \SEQCNTS_2[2]\, 
        \SEQCNTS_18[2]\, N_3836, \SEQCNTS_2[3]\, \SEQCNTS_18[3]\, 
        N_3837, \SEQCNTS_2[4]\, \SEQCNTS_18[4]\, N_3838, 
        \SEQCNTS_10[0]\, \SEQCNTS_26[0]\, N_3839, \SEQCNTS_10[1]\, 
        \SEQCNTS_26[1]\, N_3840, \SEQCNTS_10[2]\, \SEQCNTS_26[2]\, 
        N_3841, \SEQCNTS_10[3]\, \SEQCNTS_26[3]\, N_3842, 
        \SEQCNTS_10[4]\, \SEQCNTS_26[4]\, N_3843, N_3844, N_3845, 
        N_3846, N_3847, N_3848, \SEQCNTS_6[0]\, \SEQCNTS_22[0]\, 
        N_3849, \SEQCNTS_6[1]\, \SEQCNTS_22[1]\, N_3850, 
        \SEQCNTS_6[2]\, \SEQCNTS_22[2]\, N_3851, \SEQCNTS_6[3]\, 
        \SEQCNTS_22[3]\, N_3852, \SEQCNTS_6[4]\, \SEQCNTS_22[4]\, 
        N_3853, \SEQCNTS_14[0]\, \SEQCNTS_30[0]\, N_3854, 
        \SEQCNTS_14[1]\, \SEQCNTS_30[1]\, N_3855, \SEQCNTS_14[2]\, 
        \SEQCNTS_30[2]\, N_3856, \SEQCNTS_14[3]\, \SEQCNTS_30[3]\, 
        N_3857, \SEQCNTS_14[4]\, \SEQCNTS_30[4]\, N_3858, N_3859, 
        N_3860, N_3861, N_3862, N_3863, N_3864, N_3865, N_3866, 
        N_3867, N_3868, N_3869, N_3870, N_3871, N_3872, 
        \un39_n_seqcnts[2]\, \un39_n_seqcnts[4]\, 
        n_recd_ser_word167_1, \ARB_BYTE[14]_net_1\, N_3878, 
        N_3879, N_3880, N_3881, N_3882, N_3883, N_3884, N_3885, 
        N_3886, N_3887, N_3888, N_3889, N_3890, N_3891, N_3892, 
        N_3893, N_3894, N_3895, N_3896, N_3897, N_3898, N_3899, 
        N_3900, N_3901, N_3902, N_3903, N_3904, N_3905, N_3906, 
        N_3907, N_3908, N_3909, N_3910, N_3911, N_3912, N_3913, 
        N_3914, N_3915, N_3916, N_3917, N_3918, N_3919, N_3920, 
        N_3921, N_3922, N_3923, N_3924, N_3925, N_3926, N_3927, 
        N_3928, N_3929, N_3930, N_3931, N_3932, N_3933, N_3934, 
        N_3935, \BIT_OS_VAL_4[1]\, N_3936, N_3937, 
        \BIT_OS_VAL_3[3]\, \BIT_OS_VAL_4[3]\, N_3938, N_3939, 
        \BIT_OS_VAL_12[1]\, N_3940, N_3941, \BIT_OS_VAL_11[3]\, 
        N_3942, N_3943, N_3944, N_3945, N_3946, N_3947, 
        \BIT_OS_VAL_8[1]\, N_3948, N_3949, \BIT_OS_VAL_7[3]\, 
        \BIT_OS_VAL_8[3]\, N_3950, N_3951, \BIT_OS_VAL_16[1]\, 
        N_3952, N_3953, \BIT_OS_VAL_15[3]\, \BIT_OS_VAL_16[3]\, 
        N_3954, N_3955, N_3956, N_3957, N_3958, N_3959, N_3960, 
        N_3961, N_3962, N_3963, \BIT_OS_VAL_20[1]\, N_3964, 
        N_3965, \BIT_OS_VAL_19[3]\, \BIT_OS_VAL_20[3]\, N_3966, 
        N_3967, \BIT_OS_VAL_28[1]\, N_3968, N_3969, 
        \BIT_OS_VAL_27[3]\, N_3970, N_3971, N_3972, N_3973, 
        N_3974, N_3975, \BIT_OS_VAL_24[1]\, N_3976, N_3977, 
        \BIT_OS_VAL_23[3]\, \BIT_OS_VAL_24[3]\, N_3978, N_3979, 
        \BIT_OS_VAL_0[1]\, N_3980, N_3981, \BIT_OS_VAL_31[3]\, 
        \BIT_OS_VAL_0[3]\, N_3982, N_3983, N_3984, N_3985, N_3986, 
        N_3987, N_3988, N_3989, N_3990, N_3991, N_3992, N_3993, 
        N_3998, N_3999, N_4000, N_4001, N_4002, N_4003, N_4004, 
        N_4005, N_4006, N_4007, N_4008, N_4009, N_4010, N_4011, 
        N_4012, N_4013, N_4014, N_4015, N_4016, N_4017, N_4018, 
        N_4019, N_4020, N_4021, N_4022, N_4023, N_4024, N_4025, 
        N_4026, N_4027, N_4028, N_4029, N_4030, N_4031, N_4032, 
        N_4033, N_4034, N_4035, N_4036, N_4037, N_4038, N_4039, 
        N_4040, N_4041, N_4042, N_4043, N_4044, N_4045, N_4046, 
        N_4047, N_4048, N_4049, N_4050, N_4051, N_4052, N_4053, 
        N_4054, N_4055, N_4056, N_4057, N_4058, N_4059, N_4060, 
        N_4061, N_4062, N_4063, N_4064, N_4065, N_4066, N_4067, 
        N_4068, N_4069, N_4070, N_4071, N_4072, N_4073, N_4074, 
        N_4075, N_4076, N_4077, N_4078, N_4079, N_4080, N_4081, 
        N_4082, N_4083, N_4084, N_4085, N_4086, N_4087, N_4088, 
        \SEQCNTS_16[0]\, N_4089, \SEQCNTS_16[1]\, N_4090, 
        \SEQCNTS_16[2]\, N_4091, \SEQCNTS_16[3]\, N_4092, 
        \SEQCNTS_16[4]\, N_4093, N_4094, N_4095, N_4096, N_4097, 
        N_4098, N_4099, N_4100, N_4101, N_4102, N_4103, N_4104, 
        N_4105, N_4106, N_4107, N_4108, N_4109, N_4110, N_4111, 
        N_4112, N_4113, N_4114, N_4115, N_4116, N_4117, N_4118, 
        N_4119, N_4120, N_4121, N_4122, N_4128, N_4123, N_4129, 
        N_4124, N_4130, N_4125, N_4131, N_4126, N_4132, N_4127, 
        N_4133, N_4134, N_4135, N_4136, N_4137, N_4138, N_4139, 
        N_4140, N_4141, N_4142, \DES_SM_RNO[4]_net_1\, 
        \BEST_SEQCNT[1]_net_1\, \BEST_CLKPHASE[0]_net_1\, 
        I0_un1_S, \N_BIT_OS_VAL_31_18[3]\, \un36_n_bit_os_val[0]\, 
        \N_BIT_OS_VAL_30_18[3]\, \un36_n_bit_os_val[1]\, 
        \N_BIT_OS_VAL_29_18[3]\, \un36_n_bit_os_val[2]\, 
        \N_BIT_OS_VAL_28_18[3]\, \un36_n_bit_os_val[3]\, 
        \N_BIT_OS_VAL_27_18[3]\, \un36_n_bit_os_val[4]\, 
        \N_BIT_OS_VAL_26_18[3]\, \un36_n_bit_os_val[5]\, 
        \N_BIT_OS_VAL_25_18[3]\, \un36_n_bit_os_val[6]\, 
        \N_BIT_OS_VAL_24_18[3]\, \un36_n_bit_os_val[7]\, 
        \N_BIT_OS_VAL_23_18[3]\, \un36_n_bit_os_val[8]\, 
        \N_BIT_OS_VAL_22_18[3]\, \un36_n_bit_os_val[9]\, 
        \N_BIT_OS_VAL_21_18[3]\, \un36_n_bit_os_val[10]\, 
        \N_BIT_OS_VAL_20_18[3]\, \un36_n_bit_os_val[11]\, 
        \N_BIT_OS_VAL_19_18[3]\, \un36_n_bit_os_val[12]\, 
        \N_BIT_OS_VAL_18_18[3]\, \un36_n_bit_os_val[13]\, 
        \N_BIT_OS_VAL_17_18[3]\, \un36_n_bit_os_val[14]\, 
        \N_BIT_OS_VAL_16_18[3]\, \un36_n_bit_os_val[15]\, 
        \N_BIT_OS_VAL_15_18[3]\, \un36_n_bit_os_val[16]\, 
        \N_BIT_OS_VAL_13_18[3]\, \un36_n_bit_os_val[18]\, 
        \N_BIT_OS_VAL_12_18[3]\, \un36_n_bit_os_val[19]\, 
        \N_BIT_OS_VAL_11_18[3]\, \un36_n_bit_os_val[20]\, 
        \N_BIT_OS_VAL_10_18[3]\, \un36_n_bit_os_val[21]\, 
        \N_BIT_OS_VAL_9_18[3]\, \un36_n_bit_os_val[22]\, 
        \N_BIT_OS_VAL_8_18[3]\, \un36_n_bit_os_val[23]\, 
        \N_BIT_OS_VAL_7_18[3]\, \un36_n_bit_os_val[24]\, 
        BIT_OS_CNT_0e, BIT_OS_CNT_2e, N_561_3, BIT_OS_CNT_3e, 
        BIT_OS_CNT_4e, BIT_OS_CNT_6e, N_159, N_161, N_163, N_165, 
        N_167, N_169, N_171, N_173, N_5641, N_177, N_179, N_213, 
        N_216, N_219, N_5666, N_222, N_225, N_228, N_231, N_234, 
        N_237, N_240, N_243, N_246, N_249, N_252, 
        \N_INDEX_CNT[4]\, I_12_0, I_9_0, I_7_0, \N_INDEX_CNT[1]\, 
        I_5_0, \N_BEST_CLKPHASE[4]\, \N_BEST_CLKPHASE[2]\, 
        \N_BEST_CLKPHASE[1]\, \N_BEST_CLKPHASE[0]\, N_5679, N_80, 
        N_5678, N_5677, N_5676, N_5663, N_5668, N_5675, N_5674, 
        N_90, N_5673, N_5672, \N_BIT_OS_VAL_0_18[0]\, N_5662, 
        N_206, \N_BIT_OS_VAL_1_18[0]\, N_5661, N_5660, 
        \N_BIT_OS_VAL_3_18[0]\, N_5659, \N_BIT_OS_VAL_4_18[0]\, 
        N_5658, \N_BIT_OS_VAL_6_18[0]\, N_5657, N_5656, N_5655, 
        N_5654, N_5653, N_5652, N_5651, N_5650, N_5649, 
        \DES_SM_RNO[5]_net_1\, \N_BIT_OS_VAL_0_18[3]\, 
        \N_BIT_OS_VAL_1_18[3]\, \N_BIT_OS_VAL_2_18[3]\, 
        \N_BIT_OS_VAL_3_18[3]\, \N_BIT_OS_VAL_4_18[3]\, 
        \N_BIT_OS_VAL_6_18[3]\, \N_BIT_OS_VAL_14_18[3]\, N_5712, 
        N_214, N_5711, N_212, N_204, N_211, 
        \un36_n_bit_os_val[26]\, N_344, N_342, N_340, N_338, 
        N_336, N_334, N_332, N_330, N_328, N_326, N_324, N_322, 
        N_320, N_318, N_316, N_314, N_717, N_312, N_310, N_308, 
        N_306, N_304, N_302, N_300, N_298, N_296, N_294, N_292, 
        N_290, N_288, N_286, N_284, N_282, \N_BIT_OS_VAL_5_18[1]\, 
        N_279, \N_BIT_OS_VAL_7_18[1]\, N_276, 
        \N_BIT_OS_VAL_8_18[1]\, N_273, \N_BIT_OS_VAL_9_18[1]\, 
        N_270, \N_BIT_OS_VAL_10_18[1]\, \N_BIT_OS_VAL_11_18[1]\, 
        N_264, \N_BIT_OS_VAL_12_18[1]\, N_261, 
        \N_BIT_OS_VAL_13_18[1]\, N_258, \N_BIT_OS_VAL_15_18[1]\, 
        N_255, \N_BIT_OS_VAL_16_18[1]\, \N_BIT_OS_VAL_17_18[1]\, 
        \N_BIT_OS_VAL_18_18[1]\, \N_BIT_OS_VAL_19_18[1]\, 
        \N_BIT_OS_VAL_20_18[1]\, \N_BIT_OS_VAL_21_18[1]\, 
        \N_BIT_OS_VAL_22_18[1]\, \N_BIT_OS_VAL_23_18[1]\, 
        \N_BIT_OS_VAL_24_18[1]\, \N_BIT_OS_VAL_25_18[1]\, 
        \N_BIT_OS_VAL_26_18[1]\, \N_BIT_OS_VAL_27_18[1]\, 
        \N_BIT_OS_VAL_28_18[1]\, \N_BIT_OS_VAL_29_18[1]\, 
        \N_BIT_OS_VAL_30_18[1]\, \N_BIT_OS_VAL_31_18[1]\, N_207, 
        N_205, N_203, N_201, N_199, N_197, N_195, N_193, N_191, 
        N_189, N_187, N_185, N_183, N_181, \N_BIT_OS_VAL_5_18[3]\, 
        \DES_SM_RNO[1]_net_1\, N_5813, \DES_SM[3]_net_1\, 
        \DES_SM_RNO[3]_net_1\, \BIT_OS_CNT_6[3]\, 
        \BIT_OS_CNT_6[2]\, N_527, N_547, N_3658, N_3718, N_3656, 
        N_3716, N_3686, N_3684, N_3670, N_3682, N_3668, N_3680, 
        N_3674, N_3672, N_3676, N_3662, N_3666, N_3660, N_3664, 
        N_3626, N_3654, N_3624, N_3652, N_3638, N_3650, N_3610, 
        N_3622, N_3614, N_3618, N_3602, N_3606, 
        \N_BEST_CLKPHASE[3]\, N_1, \BEST_CLKPHASE[4]_net_1\, 
        \BIT_OS_CNT_4[3]\, \BIT_OS_CNT_4[2]\, N_507, N_558, N_537, 
        \DES_SM[2]_net_1\, N_54, N_49, N_5619, BIT_OS_CNT_3_n1, 
        \BIT_OS_CNT_7[0]\, N_5615, BIT_OS_CNT_7_n1, BIT_OS_CNT_7e, 
        \RECD_SER_WORD[7]_net_1\, SER_RX_IN_R, SER_RX_IN_F, 
        \BIT_OS_CNT_1[2]\, \BIT_OS_CNT_1[3]\, N_557, N_82, N_267, 
        BIT_OS_CNT_1e, N_5790, N_5810, N_5811, N_5781, N_5812, 
        N_5782, WAITCNT_n12, N_5785, N_58, N_140, N_5787, N_5780, 
        WAITCNT_n13, N_36, N_142, \CLKPHASE_RNO[0]_net_1\, 
        \TUNE_CLKPHASE[0]_net_1\, N_5797, 
        \TUNE_CLKPHASE[4]_net_1\, N_5796, 
        \TUNE_CLKPHASE[3]_net_1\, N_5795, 
        \TUNE_CLKPHASE[2]_net_1\, N_5794, 
        \TUNE_CLKPHASE[1]_net_1\, N_5793, 
        \DES_SM_RNIL6CU[5]_net_1\, N_94, 
        \DWACT_ADD_CI_0_partial_sum[0]\, I_20, I_21, I_22, I_18, 
        BIT_OS_CNT_5e, N_517, \N_BIT_OS_VAL_14_18[0]\, 
        \N_BIT_OS_VAL_2_18[0]\, \BIT_OS_CNT_2[0]\, N_5610, 
        BIT_OS_CNT_2_n1, N_210, \ADJ_SER_IN_F_0DEL\, 
        \ADJ_SER_IN_R_0DEL\, \ADJ_SER_IN_F_1DEL\, 
        \ADJ_SER_IN_R_1DEL\, \BEST_BIT_OS_VAL[3]_net_1\, 
        \BEST_SEQCNT[0]_net_1\, \ARB_WRD_40M_FIXED[0]_net_1\, 
        \Q[0]_net_1\, \ARB_WRD_40M_FIXED[1]_net_1\, \Q[1]_net_1\, 
        \ARB_WRD_40M_FIXED[2]_net_1\, \Q[2]_net_1\, 
        \ARB_WRD_40M_FIXED[3]_net_1\, \Q[3]_net_1\, 
        \ARB_WRD_40M_FIXED[4]_net_1\, \Q[4]_net_1\, 
        \ARB_WRD_40M_FIXED[5]_net_1\, \Q[5]_net_1\, 
        \ARB_WRD_40M_FIXED[6]_net_1\, \Q[6]_net_1\, 
        \ARB_WRD_40M_FIXED[7]_net_1\, \Q[7]_net_1\, 
        \ARB_WRD_40M_FIXED[8]_net_1\, \Q[8]_net_1\, 
        \ARB_WRD_40M_FIXED[9]_net_1\, \Q[9]_net_1\, 
        \ARB_WRD_40M_FIXED[10]_net_1\, \Q[10]_net_1\, 
        \ARB_WRD_40M_FIXED[11]_net_1\, \Q[11]_net_1\, 
        \ARB_WRD_40M_FIXED[12]_net_1\, \Q[12]_net_1\, 
        \ARB_WRD_40M_FIXED[13]_net_1\, \Q[13]_net_1\, 
        \ARB_WRD_40M_FIXED[14]_net_1\, \Q[14]_net_1\, 
        \ADJ_Q[0]_net_1\, \ADJ_Q[1]_net_1\, \ADJ_Q[2]_net_1\, 
        \ADJ_Q[3]_net_1\, \ADJ_Q[4]_net_1\, \ADJ_Q[5]_net_1\, 
        \ADJ_Q[6]_net_1\, \ADJ_Q[7]_net_1\, \ADJ_Q[8]_net_1\, 
        \ADJ_Q[9]_net_1\, \ADJ_Q[10]_net_1\, \ADJ_Q[11]_net_1\, 
        \ADJ_Q[12]_net_1\, \ADJ_Q[13]_net_1\, \ADJ_Q[14]_net_1\, 
        N_3, N_11, N_10, N_9, N_6, N_8, N_7, N_5, N_2_1, N_3_0, 
        N_4_1, N_3_1, \GND\, \VCC\ : std_logic;

begin 

    ELK_RX_SER_WORD_0(7) <= \ELK_RX_SER_WORD_0[7]\;
    ELK_RX_SER_WORD_0(6) <= \ELK_RX_SER_WORD_0[6]\;
    ELK_RX_SER_WORD_0(5) <= \ELK_RX_SER_WORD_0[5]\;
    ELK_RX_SER_WORD_0(4) <= \ELK_RX_SER_WORD_0[4]\;
    ELK_RX_SER_WORD_0(0) <= \ELK_RX_SER_WORD_0[0]\;
    TFC_RX_SER_WORD(7) <= \TFC_RX_SER_WORD[7]\;
    BIT_OS_SEL(2) <= \BIT_OS_SEL[2]_net_1\;
    BIT_OS_SEL(1) <= \BIT_OS_SEL[1]_net_1\;
    BIT_OS_SEL(0) <= \BIT_OS_SEL[0]_net_1\;
    BIT_OS_SEL_1(2) <= \BIT_OS_SEL_1[2]_net_1\;
    BIT_OS_SEL_1(1) <= \BIT_OS_SEL_1[1]_net_1\;
    BIT_OS_SEL_1(0) <= \BIT_OS_SEL_1[0]_net_1\;

    \CLKPHASE_0_RNIG0T43[2]\ : MX2
      port map(A => N_3610, B => N_3622, S => 
        \CLKPHASE_0[2]_net_1\, Y => N_3626);
    
    \REG40M.BIT_OS_CNT_4_RNO[8]\ : XA1C
      port map(A => \BIT_OS_CNT_4[8]\, B => N_420, C => N_4530_0, 
        Y => N_35);
    
    \BEST_BIT_OS_VAL[1]\ : DFN1E1C0
      port map(D => \N_BEST_BIT_OS_VAL[1]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_14, E => 
        un1_N_CCC_RESET_EN_0_sqmuxa, Q => 
        \BEST_BIT_OS_VAL[1]_net_1\);
    
    \ARB_BYTE_RNI8GJU_0[1]\ : NOR3B
      port map(A => \ARB_BYTE[1]_net_1\, B => N_772, C => 
        \ARB_BYTE[4]_net_1\, Y => BIT_OS_CNT_7lde_0_a3_0);
    
    \REG40M.BIT_OS_VAL_23_RNO[0]\ : MX2
      port map(A => \BIT_OS_VAL_23[0]\, B => N_5666, S => 
        \un36_n_bit_os_val[8]\, Y => N_234);
    
    \RECD_SER_WORD_RNO_6[6]\ : OA1
      port map(A => \BIT_OS_SEL[3]_net_1\, B => 
        n_recd_ser_word164, C => \ARB_BYTE[6]_net_1\, Y => 
        \ARB_BYTE_m_5[6]\);
    
    \REG40M.BIT_OS_CNT_1_RNO[5]\ : XA1C
      port map(A => \BIT_OS_CNT_1[5]\, B => N_381, C => N_4530_1, 
        Y => N_131);
    
    \REG40M.BIT_OS_CNT_1_RNO_0[8]\ : OR2A
      port map(A => \BIT_OS_CNT_1[7]\, B => N_403, Y => N_436);
    
    \CLKPHASE_0[3]\ : DFN1C0
      port map(D => \TUNE_CLKPHASE_RNILF0P2[3]_net_1\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_24_0, Q => 
        \CLKPHASE_0[3]_net_1\);
    
    \REG40M.BIT_OS_CNT_2_RNIGPSV9[1]\ : OA1C
      port map(A => N_445, B => N_437, C => N_360, Y => N_206);
    
    un1_N_CCC_RESET_EN_0_sqmuxa_0_0_a3_RNO : NOR2B
      port map(A => \DES_SM[4]_net_1\, B => N_5730, Y => 
        un1_N_CCC_RESET_EN_0_sqmuxa_0_0_a3_0);
    
    \CLKPHASE_RNIP0JI_3[0]\ : NOR2B
      port map(A => N_212, B => N_5072_2, Y => 
        \un36_n_bit_os_val[9]\);
    
    \RECD_SER_WORD_RNO_3[1]\ : NOR3C
      port map(A => n_recd_ser_word167_1, B => 
        n_recd_ser_word171_0, C => \ARB_BYTE[8]_net_1\, Y => 
        \ARB_BYTE_m[8]\);
    
    \BEST_BIT_OS_VAL_RNO_16[2]\ : MX2
      port map(A => \BIT_OS_VAL_9[2]\, B => \BIT_OS_VAL_10[2]\, S
         => \INDEX_CNT_0[0]_net_1\, Y => N_3884);
    
    \DES_SM_RNO[5]\ : OR2A
      port map(A => \DES_SM[6]_net_1\, B => 
        \un36_n_bit_os_val[1]\, Y => \DES_SM_RNO[5]_net_1\);
    
    \REG40M.BIT_OS_VAL_31_RNO[1]\ : MX2B
      port map(A => \BIT_OS_VAL_31[1]\, B => N_206_0, S => 
        \un36_n_bit_os_val[0]\, Y => \N_BIT_OS_VAL_31_18[1]\);
    
    \REG40M.SEQCNTS_3[0]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[0]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_11, E => N_340, Q => \SEQCNTS_3[0]\);
    
    \REG40M.SEQCNTS_25_RNI553P[1]\ : MX2
      port map(A => \SEQCNTS_9[1]\, B => \SEQCNTS_25[1]\, S => 
        \CLKPHASE_3[4]_net_1\, Y => N_3764);
    
    \REG40M.SEQCNTS_22[3]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[3]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_5, E => N_302, Q => \SEQCNTS_22[3]\);
    
    \REG40M.SEQCNTS_10[4]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[4]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_18, E => N_326, Q => \SEQCNTS_10[4]\);
    
    \REG40M.BIT_OS_VAL_27_RNIK79C[1]\ : MX2
      port map(A => \BIT_OS_VAL_11[1]\, B => \BIT_OS_VAL_27[1]\, 
        S => \CLKPHASE_5[4]_net_1\, Y => N_3616);
    
    \CLKPHASE_0_RNIKNR71[3]\ : MX2
      port map(A => N_3758, B => N_3763, S => 
        \CLKPHASE_0[3]_net_1\, Y => N_3768);
    
    \BIT_OS_SEL_4[0]\ : DFN1C0
      port map(D => \BEST_BIT_OS_VAL[0]_net_1\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_27_0, Q => BIT_OS_SEL_4(0));
    
    \REG40M.BIT_OS_VAL_8_RNO[2]\ : MX2
      port map(A => \BIT_OS_VAL_8[2]\, B => N_781_0, S => 
        \un36_n_bit_os_val[23]\, Y => N_203);
    
    \REG40M.BIT_OS_VAL_20_RNI03HQ[3]\ : MX2
      port map(A => \BIT_OS_VAL_4[3]\, B => \BIT_OS_VAL_20[3]\, S
         => \CLKPHASE_2[4]_net_1\, Y => N_3674);
    
    \REG40M.SEQCNTS_4[1]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[1]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_13, E => N_338, Q => \SEQCNTS_4[1]\);
    
    \REG40M.BIT_OS_VAL_9_RNI2L9J[0]\ : MX2
      port map(A => \BIT_OS_VAL_9[0]\, B => \BIT_OS_VAL_25[0]\, S
         => \CLKPHASE_0[4]_net_1\, Y => N_3631);
    
    \REG40M.BIT_OS_CNT_0_RNO[7]\ : XA1C
      port map(A => \BIT_OS_CNT_0[7]\, B => N_404, C => N_4530_2, 
        Y => N_5639);
    
    \INDEX_CNT_RNIFNQEG[1]\ : MX2
      port map(A => N_4065, B => N_4140, S => 
        \INDEX_CNT[1]_net_1\, Y => \un6_n_best_seqcnt[2]\);
    
    \REG40M.SEQCNTS_15_RNI2NAD[4]\ : MX2
      port map(A => \SEQCNTS_15[4]\, B => \SEQCNTS_16[4]\, S => 
        \INDEX_CNT_0[0]_net_1\, Y => N_4092);
    
    \REG40M.BIT_OS_VAL_4[2]\ : DFN1E1C0
      port map(D => N_5651, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_21, E => \DES_SM[6]_net_1\, Q => 
        \BIT_OS_VAL_4[2]\);
    
    \BIT_OS_SEL_6[1]\ : DFN1C0
      port map(D => \BEST_BIT_OS_VAL[1]_net_1\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_27_0, Q => BIT_OS_SEL_6(1));
    
    \REG40M.BIT_OS_VAL_19_RNO[3]\ : MX2
      port map(A => \BIT_OS_VAL_19[3]\, B => N_209_0, S => 
        \un36_n_bit_os_val[12]\, Y => \N_BIT_OS_VAL_19_18[3]\);
    
    \REG40M.BIT_OS_CNT_1_RNO[0]\ : NOR2
      port map(A => \BIT_OS_CNT_1[0]\, B => N_4530, Y => N_557);
    
    \CLKPHASE_1_RNIPDI72[2]\ : MX2
      port map(A => N_3770, B => N_3785, S => 
        \CLKPHASE_1[2]_net_1\, Y => N_3790);
    
    \CLKPHASE_1_RNILS5B1[3]\ : MX2
      port map(A => N_3660, B => N_3664, S => 
        \CLKPHASE_1[3]_net_1\, Y => N_3668);
    
    \REG40M.SEQCNTS_7_RNIJJ051[3]\ : MX2
      port map(A => \SEQCNTS_7[3]\, B => \SEQCNTS_8[3]\, S => 
        \INDEX_CNT[0]_net_1\, Y => N_4086);
    
    \REG40M.BIT_OS_VAL_27[3]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_27_18[3]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_2, E => \DES_SM_0[6]_net_1\, Q
         => \BIT_OS_VAL_27[3]\);
    
    \CLKPHASE_RNI8UD7[2]\ : OR2A
      port map(A => \CLKPHASE[0]_net_1\, B => \CLKPHASE[2]_net_1\, 
        Y => N_5668);
    
    \BEST_BIT_OS_VAL_RNO_1[2]\ : MX2
      port map(A => N_3904, B => N_3928, S => 
        \INDEX_CNT[4]_net_1\, Y => N_3932);
    
    \REG40M.BIT_OS_VAL_20_RNO[0]\ : MX2
      port map(A => \BIT_OS_VAL_20[0]\, B => N_5666_0, S => 
        \un36_n_bit_os_val[11]\, Y => N_243);
    
    \CLKPHASE_RNIG15B[3]\ : OR3A
      port map(A => \CLKPHASE[3]_net_1\, B => \CLKPHASE[0]_net_1\, 
        C => \CLKPHASE[4]_net_1\, Y => N_5672);
    
    \RECD_SER_WORD_RNO_4[7]\ : NOR3C
      port map(A => n_recd_ser_word168_2, B => 
        n_recd_ser_word169_0, C => \ARB_BYTE[12]_net_1\, Y => 
        \ARB_BYTE_m_1[12]\);
    
    un1_CLKPHASE_I_16 : XOR2
      port map(A => \CLKPHASE[0]_net_1\, B => 
        \DES_SM_RNIL6CU[5]_net_1\, Y => 
        \DWACT_ADD_CI_0_partial_sum[0]\);
    
    \Q[7]\ : DFN1C0
      port map(D => \ADJ_Q[7]_net_1\, CLK => CCC_160M_FXD, CLR
         => P_MASTER_POR_B_c_34, Q => \Q[7]_net_1\);
    
    \REG40M.BIT_OS_VAL_5[1]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_5_18[1]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_1, E => \DES_SM_0[6]_net_1\, Q
         => \BIT_OS_VAL_5[1]\);
    
    \REG40M.BIT_OS_CNT_5_RNIGBFI1[6]\ : OR3B
      port map(A => \BIT_OS_CNT_5[5]\, B => \BIT_OS_CNT_5[6]\, C
         => N_384, Y => N_409);
    
    \MAX_CNT[2]\ : DFN1E0C0
      port map(D => N_5638, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_16, E => N_558, Q => \MAX_CNT[2]_net_1\);
    
    \INDEX_CNT_0_RNIAHTE3[2]\ : MX2
      port map(A => N_4116, B => N_4131, S => 
        \INDEX_CNT_0[2]_net_1\, Y => N_4136);
    
    \INDEX_CNT[2]\ : DFN1E0C0
      port map(D => \N_INDEX_CNT[2]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_17, E => N_5149, Q => 
        \INDEX_CNT[2]_net_1\);
    
    \BEST_BIT_OS_VAL_RNO[3]\ : NOR2A
      port map(A => \N_BEST_BIT_OS_VAL_3[3]\, B => 
        \DES_SM[8]_net_1\, Y => \N_BEST_BIT_OS_VAL[3]\);
    
    \RECD_SER_WORD_RNIKKBK[7]\ : NOR2B
      port map(A => \RECD_SER_WORD[7]_net_1\, B => DCB_SALT_SEL_c, 
        Y => \ELK_RX_SER_WORD_0[7]\);
    
    \REG40M.SEQCNTS_29_RNIBFG41[4]\ : MX2
      port map(A => N_4052, B => \SEQCNTS_29[4]\, S => 
        \INDEX_CNT_2[3]_net_1\, Y => N_4057);
    
    \ARB_BYTE[11]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[11]_net_1\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_32_0, Q => 
        \ARB_BYTE[11]_net_1\);
    
    \REG40M.BIT_OS_CNT_4_RNO_0[2]\ : AOI1
      port map(A => \BIT_OS_CNT_4[1]\, B => \BIT_OS_CNT_4[0]\, C
         => \BIT_OS_CNT_4[2]\, Y => N_505);
    
    \REG40M.BIT_OS_CNT_1_RNIABF8[4]\ : OR3
      port map(A => \BIT_OS_CNT_1[6]\, B => \BIT_OS_CNT_1[4]\, C
         => \BIT_OS_CNT_1[5]\, Y => N_BIT_OS_VAL_316lto8_0_o3_2);
    
    \REG40M.SEQCNTS_13_RNILGFE[2]\ : MX2
      port map(A => \SEQCNTS_13[2]\, B => \SEQCNTS_29[2]\, S => 
        \CLKPHASE_2[4]_net_1\, Y => N_3780);
    
    \DES_SM_0_RNI05GJ3[8]\ : AO1
      port map(A => DES_SM_tr2_i_a3_6, B => DES_SM_tr2_i_a3_5, C
         => \DES_SM_0[8]_net_1\, Y => un1_DES_SM_19);
    
    \WAITCNT_RNO[8]\ : NOR3A
      port map(A => N_5779, B => N_5807, C => N_4539, Y => N_5718);
    
    \MAX_CNT_RNO_0[2]\ : AOI1
      port map(A => \MAX_CNT[1]_net_1\, B => \MAX_CNT[0]_net_1\, 
        C => \MAX_CNT[2]_net_1\, Y => N_535);
    
    \REG40M.BIT_OS_CNT_7_RNIB4QI[6]\ : OR2
      port map(A => \BIT_OS_CNT_7[7]\, B => \BIT_OS_CNT_7[6]\, Y
         => N_BIT_OS_VAL_3130lto8_1);
    
    \REG40M.SEQCNTS_5[1]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[1]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_15, E => N_336, Q => \SEQCNTS_5[1]\);
    
    \REG40M.BIT_OS_VAL_1[2]\ : DFN1E1C0
      port map(D => N_5654, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_17_0, E => \DES_SM_3[6]_net_1\, Q => 
        \BIT_OS_VAL_1[2]\);
    
    \RECD_SER_WORD_RNO_5[5]\ : NOR3C
      port map(A => n_recd_ser_word165_2, B => 
        n_recd_ser_word166_0, C => \ARB_BYTE[7]_net_1\, Y => 
        \ARB_BYTE_m_4[7]\);
    
    \REG40M.BIT_OS_VAL_10_RNO[2]\ : MX2
      port map(A => \BIT_OS_VAL_10[2]\, B => N_781, S => 
        \un36_n_bit_os_val[21]\, Y => N_199);
    
    \CLKPHASE_RNIDPPFC[0]\ : MX2
      port map(A => N_BIT_OS_VAL_312, B => N_BIT_OS_VAL_316, S
         => \un107_bit_os_val[0]\, Y => N_1151_tz);
    
    \WAITCNT[2]\ : DFN1E0C0
      port map(D => N_41, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_9, E => N_5790, Q => \WAITCNT[2]_net_1\);
    
    \INDEX_CNT_RNI41T63[2]\ : MX2
      port map(A => N_4044, B => N_4054, S => 
        \INDEX_CNT[2]_net_1\, Y => N_4059);
    
    \REG40M.SEQCNTS_5[2]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[2]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_15, E => N_336, Q => \SEQCNTS_5[2]\);
    
    \REG40M.BIT_OS_VAL_5[3]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_5_18[3]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_1, E => \DES_SM_0[6]_net_1\, Q
         => \BIT_OS_VAL_5[3]\);
    
    \DES_SM_RNO[0]\ : AO1A
      port map(A => N_5859, B => \DES_SM[0]_net_1\, C => 
        \DES_SM[1]_net_1\, Y => \DES_SM_RNO[0]_net_1\);
    
    \BEST_BIT_OS_VAL_RNO_1[0]\ : MX2
      port map(A => N_3902, B => N_3926, S => 
        \INDEX_CNT[4]_net_1\, Y => N_3930);
    
    \BEST_BIT_OS_VAL_RNO_14[1]\ : MX2
      port map(A => N_3975, B => N_3979, S => 
        \INDEX_CNT_2[3]_net_1\, Y => N_3983);
    
    \REG40M.BIT_OS_VAL_11[3]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_11_18[3]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_8, E => \DES_SM_1[6]_net_1\, Q
         => \BIT_OS_VAL_11[3]\);
    
    \REG40M.BIT_OS_CNT_5_RNO[3]\ : XA1C
      port map(A => \BIT_OS_CNT_5[3]\, B => N_373, C => N_4530, Y
         => N_5629);
    
    \BEST_BIT_OS_VAL_RNO_9[3]\ : MX2
      port map(A => N_3909, B => N_3913, S => 
        \INDEX_CNT[3]_net_1\, Y => N_3917);
    
    \BEST_BIT_OS_VAL[0]\ : DFN1E1C0
      port map(D => \N_BEST_BIT_OS_VAL[0]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_13, E => 
        un1_N_CCC_RESET_EN_0_sqmuxa, Q => 
        \BEST_BIT_OS_VAL[0]_net_1\);
    
    un3_n_index_cnt_I_12 : XOR2
      port map(A => N_2_0, B => \INDEX_CNT[4]_net_1\, Y => I_12_0);
    
    \REG40M.BIT_OS_CNT_2[5]\ : DFN1E1C0
      port map(D => BIT_OS_CNT_2_n5, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_5, E => BIT_OS_CNT_2e, Q => 
        \BIT_OS_CNT_2[5]\);
    
    \RECD_SER_WORD_RNO_7[6]\ : AO1
      port map(A => n_recd_ser_word165, B => \ARB_BYTE[7]_net_1\, 
        C => \ARB_BYTE_m_3[9]\, Y => \N_RECD_SER_WORD_iv_3[6]\);
    
    \CLKPHASE_1_RNIOG4D[2]\ : NOR3B
      port map(A => \CLKPHASE_0[1]_net_1\, B => N_211, C => 
        \CLKPHASE_1[2]_net_1\, Y => \un36_n_bit_os_val[5]\);
    
    \REG40M.SEQCNTS_7_RNIFF051[1]\ : MX2
      port map(A => \SEQCNTS_7[1]\, B => \SEQCNTS_8[1]\, S => 
        \INDEX_CNT[0]_net_1\, Y => N_4084);
    
    \REG40M.SEQCNTS_11_RNIUAU81[4]\ : MX2
      port map(A => \SEQCNTS_11[4]\, B => \SEQCNTS_12[4]\, S => 
        \INDEX_CNT_4[0]_net_1\, Y => N_4077);
    
    \REG40M.BIT_OS_VAL_29_RNO[3]\ : MX2
      port map(A => \BIT_OS_VAL_29[3]\, B => N_209, S => 
        \un36_n_bit_os_val[2]\, Y => \N_BIT_OS_VAL_29_18[3]\);
    
    \RECD_SER_WORD_RNO_1[5]\ : AO1
      port map(A => \ARB_BYTE[9]_net_1\, B => n_recd_ser_word168, 
        C => \ARB_BYTE_m_1[10]\, Y => \N_RECD_SER_WORD_iv_0[5]\);
    
    \REG40M.BIT_OS_VAL_22[1]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_22_18[1]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_15, E => \DES_SM_3[6]_net_1\, Q
         => \BIT_OS_VAL_22[1]\);
    
    \INDEX_CNT_RNI273N4[2]\ : MX2
      port map(A => N_4081, B => N_4096, S => 
        \INDEX_CNT[2]_net_1\, Y => N_4101);
    
    \REG40M.BIT_OS_VAL_0_RNO[1]\ : MX2A
      port map(A => N_206, B => \BIT_OS_VAL_0[1]\, S => N_5679, Y
         => N_5662);
    
    \DES_SM_RNO_0[3]\ : NOR3B
      port map(A => \DES_SM_i_0[5]\, B => CCC_RX_CLK_LOCK, C => 
        \WAITCNT[0]_net_1\, Y => \DES_SM_ns_i_a2_0_0_a3_0_1[5]\);
    
    \ARB_BYTE[3]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[3]_net_1\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_27, Q => 
        \ARB_BYTE[3]_net_1\);
    
    \WAITCNT_RNIDH6C3[12]\ : OR2A
      port map(A => \WAITCNT[12]_net_1\, B => N_5785, Y => N_5787);
    
    \REG40M.BIT_OS_VAL_0[0]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_0_18[0]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_15, E => \DES_SM_2[6]_net_1\, Q
         => \BIT_OS_VAL_0[0]\);
    
    ADJ_SER_IN_F_0DEL : DFN1C0
      port map(D => SER_RX_IN_F, CLK => CCC_160M_ADJ, CLR => 
        P_MASTER_POR_B_c_31_0, Q => \ADJ_SER_IN_F_0DEL\);
    
    \INDEX_CNT_2_RNIVDAR1[3]\ : MX2
      port map(A => N_4087, B => N_4092, S => 
        \INDEX_CNT_2[3]_net_1\, Y => N_4097);
    
    \REG40M.SEQCNTS_19[1]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[1]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_11, E => N_308, Q => \SEQCNTS_19[1]\);
    
    \REG40M.SEQCNTS_18[0]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[0]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_8, E => N_310, Q => \SEQCNTS_18[0]\);
    
    \CLKPHASE_0_RNI8OLNH7_0[2]\ : AO1A
      port map(A => N_5678, B => N_782_0, C => N_717_0, Y => 
        N_342);
    
    \REG40M.BIT_OS_CNT_5[0]\ : DFN1E1C0
      port map(D => N_517, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_11, E => BIT_OS_CNT_5e, Q => 
        \BIT_OS_CNT_5[0]\);
    
    \REG40M.BIT_OS_CNT_1_RNO[8]\ : XA1C
      port map(A => \BIT_OS_CNT_1[8]\, B => N_436, C => N_4530_1, 
        Y => N_125);
    
    \WAITCNT_RNO[6]\ : XA1C
      port map(A => \WAITCNT[6]_net_1\, B => N_5776, C => N_4539, 
        Y => N_32);
    
    \REG40M.SEQCNTS_7[3]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[3]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_17_0, E => N_332, Q => \SEQCNTS_7[3]\);
    
    \REG40M.BIT_OS_VAL_3[3]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_3_18[3]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_19, E => \DES_SM_4[6]_net_1\, Q
         => \BIT_OS_VAL_3[3]\);
    
    \REG40M.BIT_OS_CNT_5_RNO_0[6]\ : OA1C
      port map(A => \BIT_OS_CNT_5[5]\, B => N_384, C => 
        \BIT_OS_CNT_5[6]\, Y => N_511);
    
    \REG40M.BIT_OS_VAL_10_RNO[3]\ : MX2
      port map(A => \BIT_OS_VAL_10[3]\, B => N_209_0, S => 
        \un36_n_bit_os_val[21]\, Y => \N_BIT_OS_VAL_10_18[3]\);
    
    \REG40M.BIT_OS_CNT_3_RNO[7]\ : XA1B
      port map(A => BIT_OS_CNT_3_c6, B => \BIT_OS_CNT_3[7]\, C
         => N_4530_1, Y => BIT_OS_CNT_3_n7);
    
    \RECD_SER_WORD_RNIIIBK_0[5]\ : NOR2A
      port map(A => \RECD_SER_WORD[5]_net_1\, B => DCB_SALT_SEL_c, 
        Y => TFC_RX_SER_WORD(5));
    
    \CLKPHASE_RNI9DM65[1]\ : MX2
      port map(A => N_3828, B => N_3863, S => \CLKPHASE[1]_net_1\, 
        Y => N_3868);
    
    \TUNE_CLKPHASE_RNITINS2[4]\ : AO1A
      port map(A => N_5780, B => \TUNE_CLKPHASE[4]_net_1\, C => 
        N_5796, Y => \TUNE_CLKPHASE_RNITINS2[4]_net_1\);
    
    \REG40M.BIT_OS_CNT_0_RNIVKBA[5]\ : OR2A
      port map(A => \BIT_OS_CNT_0[5]\, B => N_383, Y => N_390);
    
    \DES_SM[2]\ : DFN1C0
      port map(D => N_36, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_26, Q => \DES_SM[2]_net_1\);
    
    \CLKPHASE_2_RNI801I1[3]\ : MX2
      port map(A => N_3599, B => N_3603, S => 
        \CLKPHASE_2[3]_net_1\, Y => N_3607);
    
    \BIT_OS_SEL_0[0]\ : DFN1C0
      port map(D => \BEST_BIT_OS_VAL[0]_net_1\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_27_0, Q => BIT_OS_SEL_0(0));
    
    \REG40M.SEQCNTS_1_RNIGH6J[0]\ : MX2
      port map(A => \SEQCNTS_1[0]\, B => \SEQCNTS_2[0]\, S => 
        \INDEX_CNT_0[0]_net_1\, Y => N_3998);
    
    \REG40M.SEQCNTS_19_RNI0LGG[1]\ : MX2
      port map(A => \SEQCNTS_3[1]\, B => \SEQCNTS_19[1]\, S => 
        \CLKPHASE_1[4]_net_1\, Y => N_3739);
    
    \RECD_SER_WORD_RNO[1]\ : OR3
      port map(A => \N_RECD_SER_WORD_iv_1[1]\, B => 
        \N_RECD_SER_WORD_iv_0[1]\, C => \N_RECD_SER_WORD_iv_5[1]\, 
        Y => \N_RECD_SER_WORD[1]\);
    
    \REG40M.BIT_OS_VAL_19[2]\ : DFN1E1C0
      port map(D => N_183, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_20, E => \DES_SM[6]_net_1\, Q => 
        \BIT_OS_VAL_19[2]\);
    
    \REG40M.BIT_OS_VAL_10_RNO[1]\ : MX2B
      port map(A => \BIT_OS_VAL_10[1]\, B => N_206, S => 
        \un36_n_bit_os_val[21]\, Y => \N_BIT_OS_VAL_10_18[1]\);
    
    \REG40M.BIT_OS_CNT_4_RNO[6]\ : NOR3A
      port map(A => N_410, B => N_501, C => N_4530_0, Y => N_5621);
    
    \INDEX_CNT_RNILSDH8[4]\ : MX2
      port map(A => N_4100, B => N_4135, S => 
        \INDEX_CNT[4]_net_1\, Y => N_4140);
    
    \REG40M.SEQCNTS_2[3]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[3]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_10, E => N_342, Q => \SEQCNTS_2[3]\);
    
    \RECD_SER_WORD_RNO_2[1]\ : OR3
      port map(A => \ARB_BYTE_m_0[3]\, B => \ARB_BYTE_m_0[1]\, C
         => \N_RECD_SER_WORD_iv_3[1]\, Y => 
        \N_RECD_SER_WORD_iv_5[1]\);
    
    \RECD_SER_WORD_RNO_4[5]\ : NOR3C
      port map(A => n_recd_ser_word168_2, B => 
        n_recd_ser_word169_0, C => \ARB_BYTE[10]_net_1\, Y => 
        \ARB_BYTE_m_1[10]\);
    
    \REG40M.BIT_OS_VAL_20_RNO[2]\ : MX2
      port map(A => \BIT_OS_VAL_20[2]\, B => N_781_0, S => 
        \un36_n_bit_os_val[11]\, Y => N_181);
    
    \RECD_SER_WORD_RNO_8[1]\ : NOR3C
      port map(A => n_recd_ser_word165_2, B => 
        n_recd_ser_word167_1, C => \ARB_BYTE[4]_net_1\, Y => 
        \ARB_BYTE_m_0[4]\);
    
    \REG40M.SEQCNTS_15_RNISGAD[1]\ : MX2
      port map(A => \SEQCNTS_15[1]\, B => \SEQCNTS_16[1]\, S => 
        \INDEX_CNT_0[0]_net_1\, Y => N_4089);
    
    \RECD_SER_WORD_RNIDDBK_0[0]\ : NOR2A
      port map(A => \RECD_SER_WORD[0]_net_1\, B => DCB_SALT_SEL_c, 
        Y => TFC_RX_SER_WORD(0));
    
    \BEST_BIT_OS_VAL_RNO_24[3]\ : MX2
      port map(A => \BIT_OS_VAL_7[3]\, B => \BIT_OS_VAL_8[3]\, S
         => \INDEX_CNT_2[0]_net_1\, Y => N_3949);
    
    \BIT_OS_SEL_6[2]\ : DFN1C0
      port map(D => \BEST_BIT_OS_VAL[2]_net_1\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_27_0, Q => BIT_OS_SEL_6(2));
    
    \BEST_BIT_OS_VAL_RNO_29[1]\ : MX2
      port map(A => \BIT_OS_VAL_31[1]\, B => \BIT_OS_VAL_0[1]\, S
         => \INDEX_CNT_3[0]_net_1\, Y => N_3979);
    
    \REG40M.SEQCNTS_20_RNI3VMJ[3]\ : MX2
      port map(A => \SEQCNTS_19[3]\, B => \SEQCNTS_20[3]\, S => 
        \INDEX_CNT_4[0]_net_1\, Y => N_4106);
    
    \ARB_BYTE[9]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[9]_net_1\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_27_1, Q => 
        \ARB_BYTE[9]_net_1\);
    
    \REG40M.BIT_OS_VAL_29_RNI60FE[2]\ : MX2
      port map(A => \BIT_OS_VAL_13[2]\, B => \BIT_OS_VAL_29[2]\, 
        S => \CLKPHASE[4]_net_1\, Y => N_3645);
    
    \REG40M.SEQCNTS_30_RNITFVA[2]\ : MX2
      port map(A => \SEQCNTS_14[2]\, B => \SEQCNTS_30[2]\, S => 
        \CLKPHASE[4]_net_1\, Y => N_3855);
    
    \DES_SM_RNO[4]\ : AO1
      port map(A => N_5730, B => \DES_SM[4]_net_1\, C => N_5072, 
        Y => \DES_SM_RNO[4]_net_1\);
    
    \REG40M.SEQCNTS_6[3]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[3]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_16, E => N_334, Q => \SEQCNTS_6[3]\);
    
    \REG40M.SEQCNTS_12[4]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[4]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_21, E => N_322, Q => \SEQCNTS_12[4]\);
    
    \CLKPHASE_RNIAB7UH7[0]\ : AO1
      port map(A => \un36_n_bit_os_val[26]\, B => N_782_0, C => 
        N_717_0, Y => N_336);
    
    \REG40M.SEQCNTS_11_RNIO4U81[1]\ : MX2
      port map(A => \SEQCNTS_11[1]\, B => \SEQCNTS_12[1]\, S => 
        \INDEX_CNT_4[0]_net_1\, Y => N_4074);
    
    \CLKPHASE_0_RNIEDCJ5[1]\ : MX2
      port map(A => N_3684, B => N_3712, S => 
        \CLKPHASE_0[1]_net_1\, Y => N_3716);
    
    \REG40M.SEQCNTS_23_RNIQCAH[1]\ : MX2
      port map(A => \SEQCNTS_23[1]\, B => \SEQCNTS_24[1]\, S => 
        \INDEX_CNT_0[0]_net_1\, Y => N_4119);
    
    \BIT_OS_SEL_5[2]\ : DFN1C0
      port map(D => \BEST_BIT_OS_VAL[2]_net_1\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_27_0, Q => BIT_OS_SEL_5(2));
    
    \REG40M.SEQCNTS_26[4]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[4]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_12, E => N_294, Q => \SEQCNTS_26[4]\);
    
    \REG40M.SEQCNTS_15[0]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[0]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_4, E => N_316, Q => \SEQCNTS_15[0]\);
    
    \INDEX_CNT_RNI56ST1[3]\ : MX2
      port map(A => N_4103, B => N_4108, S => 
        \INDEX_CNT[3]_net_1\, Y => N_4113);
    
    \INDEX_CNT_1_RNIGSNV1[3]\ : MX2
      port map(A => N_4002, B => N_4007, S => 
        \INDEX_CNT_1[3]_net_1\, Y => N_4012);
    
    \REG40M.BIT_OS_VAL_27_RNIOB9C[3]\ : MX2
      port map(A => \BIT_OS_VAL_11[3]\, B => \BIT_OS_VAL_27[3]\, 
        S => \CLKPHASE_5[4]_net_1\, Y => N_3618);
    
    \INDEX_CNT_0_RNIS2TE3[2]\ : MX2
      port map(A => N_4114, B => N_4129, S => 
        \INDEX_CNT_0[2]_net_1\, Y => N_4134);
    
    \CLKPHASE_RNIG15B_0[0]\ : NOR2A
      port map(A => N_204, B => \CLKPHASE[0]_net_1\, Y => N_212);
    
    \BEST_SEQCNT[0]\ : DFN1E1C0
      port map(D => \N_BEST_SEQCNT[0]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_8, E => N_5724, Q => 
        \BEST_SEQCNT[0]_net_1\);
    
    \REG40M.BIT_OS_VAL_1_RNO[1]\ : MX2A
      port map(A => N_206_0, B => \BIT_OS_VAL_1[1]\, S => N_5676, 
        Y => N_5661);
    
    \RECD_SER_WORD_RNIGGBK[3]\ : NOR2B
      port map(A => \RECD_SER_WORD[3]_net_1\, B => DCB_SALT_SEL_c, 
        Y => ELK_RX_SER_WORD_0(3));
    
    \CLKPHASE_0_RNI30JF2[2]\ : MX2
      port map(A => N_3667, B => N_3679, S => 
        \CLKPHASE_0[2]_net_1\, Y => N_3683);
    
    \INDEX_CNT[4]\ : DFN1E0C0
      port map(D => \N_INDEX_CNT[4]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_17, E => N_5149, Q => 
        \INDEX_CNT[4]_net_1\);
    
    \REG40M.BIT_OS_VAL_20_RNO[3]\ : MX2
      port map(A => \BIT_OS_VAL_20[3]\, B => N_209, S => 
        \un36_n_bit_os_val[11]\, Y => \N_BIT_OS_VAL_20_18[3]\);
    
    \RECD_SER_WORD_RNIKKBK_0[7]\ : NOR2A
      port map(A => \RECD_SER_WORD[7]_net_1\, B => DCB_SALT_SEL_c, 
        Y => \TFC_RX_SER_WORD[7]\);
    
    \DES_SM_RNIU9F02[0]\ : NOR3A
      port map(A => I_22, B => \DES_SM_0[8]_net_1\, C => 
        \DES_SM[0]_net_1\, Y => N_5794);
    
    \REG40M.BIT_OS_CNT_5_RNID6KL[1]\ : NOR3C
      port map(A => \BIT_OS_CNT_5[2]\, B => \BIT_OS_CNT_5[1]\, C
         => \BIT_OS_CNT_5[3]\, Y => N_760);
    
    \REG40M.BIT_OS_CNT_1_RNO[7]\ : XA1C
      port map(A => \BIT_OS_CNT_1[7]\, B => N_403, C => N_4530_1, 
        Y => N_127);
    
    \ALIGN_ACTIVE\ : DFN1E1C0
      port map(D => OP_MODE_c_0, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_9, E => \DES_SM_0[8]_net_1\, Q => 
        ALIGN_ACTIVE);
    
    un1_CLKPHASE_I_21 : XOR2
      port map(A => \CLKPHASE[3]_net_1\, B => 
        \DWACT_ADD_CI_0_g_array_12[0]\, Y => I_21);
    
    \RECD_SER_WORD_RNIV92L2[1]\ : NOR3C
      port map(A => \TFC_RX_SER_WORD[7]\, B => TFC_SYNC_DET_1_1, 
        C => TFC_SYNC_DET_1_4, Y => TFC_SYNC_DET_1);
    
    \REG40M.SEQCNTS_20_RNI51NJ[4]\ : MX2
      port map(A => \SEQCNTS_19[4]\, B => \SEQCNTS_20[4]\, S => 
        \INDEX_CNT_4[0]_net_1\, Y => N_4107);
    
    \CLKPHASE_RNICU2EH7[2]\ : AO1
      port map(A => \un36_n_bit_os_val[15]\, B => N_782_0, C => 
        N_717, Y => N_314);
    
    \REG40M.BIT_OS_CNT_5_RNO[0]\ : NOR2
      port map(A => \BIT_OS_CNT_5[0]\, B => N_4530, Y => N_517);
    
    \REG40M.SEQCNTS_14[2]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[2]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_2, E => N_318, Q => \SEQCNTS_14[2]\);
    
    \REG40M.BIT_OS_VAL_20_RNO[1]\ : MX2B
      port map(A => \BIT_OS_VAL_20[1]\, B => N_206_0, S => 
        \un36_n_bit_os_val[11]\, Y => \N_BIT_OS_VAL_20_18[1]\);
    
    \REG40M.SEQCNTS_22_RNIVMMK[0]\ : MX2
      port map(A => \SEQCNTS_6[0]\, B => \SEQCNTS_22[0]\, S => 
        \CLKPHASE_5[4]_net_1\, Y => N_3848);
    
    \CLKPHASE_RNIP0JI_4[1]\ : NOR2B
      port map(A => N_5712, B => N_5711, Y => 
        \un36_n_bit_os_val[20]\);
    
    \REG40M.BIT_OS_VAL_16[0]\ : DFN1E1C0
      port map(D => N_255, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_16, E => \DES_SM_3[6]_net_1\, Q => 
        \BIT_OS_VAL_16[0]\);
    
    \REG40M.BIT_OS_VAL_14_RNO[2]\ : MX2
      port map(A => N_781_0, B => \BIT_OS_VAL_14[2]\, S => N_5673, 
        Y => N_5649);
    
    \RECD_SER_WORD_RNO_4[1]\ : NOR3C
      port map(A => n_recd_ser_word168_2, B => 
        n_recd_ser_word169_0, C => \ARB_BYTE[6]_net_1\, Y => 
        \ARB_BYTE_m_0[6]\);
    
    \CLKPHASE_RNIUHVV03[0]\ : AO1
      port map(A => un1_DES_SM_1034_i_a2_0_1, B => N_427, C => 
        N_758, Y => un1_DES_SM_1034_i_o2_1);
    
    \DES_SM_RNIUEK921[6]\ : NOR3C
      port map(A => \un107_bit_os_val[0]\, B => 
        \un107_bit_os_val[1]\, C => N_761, Y => 
        un1_DES_SM_1034_i_a2_0_1);
    
    \DES_SM_0_RNI3ECBA[8]\ : NOR2
      port map(A => \un39_n_seqcnts[0]\, B => \DES_SM_0[8]_net_1\, 
        Y => \N_SEQCNTS_1_0[0]\);
    
    \RECD_SER_WORD_RNO_6[7]\ : OA1
      port map(A => \BIT_OS_SEL[3]_net_1\, B => 
        n_recd_ser_word164, C => \ARB_BYTE[7]_net_1\, Y => 
        \ARB_BYTE_m_6[7]\);
    
    \DES_SM_0_RNIAB7UH7_2[8]\ : AO1
      port map(A => \un36_n_bit_os_val[19]\, B => N_782_0, C => 
        N_717_0, Y => N_322);
    
    \DES_SM_0_RNIII0V_2[8]\ : NOR2A
      port map(A => \DES_SM_0[8]_net_1\, B => \DES_SM_0[6]_net_1\, 
        Y => N_717_0);
    
    \REG40M.BIT_OS_CNT_4[7]\ : DFN1E1C0
      port map(D => N_5620, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_9, E => BIT_OS_CNT_4e, Q => 
        \BIT_OS_CNT_4[7]\);
    
    \REG40M.BIT_OS_VAL_30[1]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_30_18[1]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_18, E => \DES_SM_4[6]_net_1\, Q
         => \BIT_OS_VAL_30[1]\);
    
    \BEST_BIT_OS_VAL_RNO_18[3]\ : MX2
      port map(A => \BIT_OS_VAL_13[3]\, B => \BIT_OS_VAL_14[3]\, 
        S => \INDEX_CNT_2[0]_net_1\, Y => N_3897);
    
    \REG40M.SEQCNTS_27_RNIN0OU[3]\ : MX2
      port map(A => \SEQCNTS_27[3]\, B => \SEQCNTS_28[3]\, S => 
        \INDEX_CNT[0]_net_1\, Y => N_4111);
    
    \REG40M.BIT_OS_VAL_8_RNI5M6I[2]\ : MX2
      port map(A => \BIT_OS_VAL_8[2]\, B => \BIT_OS_VAL_24[2]\, S
         => \CLKPHASE_1[4]_net_1\, Y => N_3665);
    
    \REG40M.BIT_OS_CNT_2[8]\ : DFN1E1C0
      port map(D => BIT_OS_CNT_2_n8, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_6, E => BIT_OS_CNT_2e, Q => 
        \BIT_OS_CNT_2[8]\);
    
    \DES_SM_RNO_1[2]\ : AOI1
      port map(A => OP_MODE_c_0, B => \DES_SM_0[8]_net_1\, C => 
        \DES_SM[2]_net_1\, Y => N_142);
    
    \BEST_BIT_OS_VAL_RNO_7[2]\ : MX2
      port map(A => N_3880, B => N_3884, S => 
        \INDEX_CNT_0[3]_net_1\, Y => N_3888);
    
    \REG40M.BIT_OS_VAL_3_RNIA0D21[3]\ : MX2
      port map(A => \BIT_OS_VAL_3[3]\, B => \BIT_OS_VAL_19[3]\, S
         => \CLKPHASE_5[4]_net_1\, Y => N_3614);
    
    \REG40M.BIT_OS_VAL_21[3]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_21_18[3]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_14, E => \DES_SM_2[6]_net_1\, Q
         => \BIT_OS_VAL_21[3]\);
    
    \WAITCNT_RNIRKL51[5]\ : OR2A
      port map(A => \WAITCNT[5]_net_1\, B => N_5775, Y => N_5776);
    
    \REG40M.SEQCNTS_19[0]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[0]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_10, E => N_308, Q => \SEQCNTS_19[0]\);
    
    \REG40M.BIT_OS_VAL_18_RNO[0]\ : MX2
      port map(A => \BIT_OS_VAL_18[0]\, B => N_5666_0, S => 
        \un36_n_bit_os_val[13]\, Y => N_249);
    
    \REG40M.SEQCNTS_18[4]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[4]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_8, E => N_310, Q => \SEQCNTS_18[4]\);
    
    \BEST_BIT_OS_VAL_RNO_16[3]\ : MX2
      port map(A => \BIT_OS_VAL_9[3]\, B => \BIT_OS_VAL_10[3]\, S
         => \INDEX_CNT_0[0]_net_1\, Y => N_3885);
    
    \REG40M.SEQCNTS_21_RNIRB7G[2]\ : MX2
      port map(A => \SEQCNTS_21[2]\, B => \SEQCNTS_22[2]\, S => 
        \INDEX_CNT_3[0]_net_1\, Y => N_4050);
    
    \REG40M.BIT_OS_CNT_2[1]\ : DFN1E1C0
      port map(D => BIT_OS_CNT_2_n1, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_5, E => BIT_OS_CNT_2e, Q => 
        \BIT_OS_CNT_2[1]\);
    
    \REG40M.SEQCNTS_18[1]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[1]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_8, E => N_310, Q => \SEQCNTS_18[1]\);
    
    \REG40M.BIT_OS_VAL_15_RNO[0]\ : MX2
      port map(A => \BIT_OS_VAL_15[0]\, B => N_5666, S => 
        \un36_n_bit_os_val[16]\, Y => N_258);
    
    \CLKPHASE_2_RNI56621[3]\ : MX2
      port map(A => N_3801, B => N_3806, S => 
        \CLKPHASE_2[3]_net_1\, Y => N_3811);
    
    \REG40M.BIT_OS_VAL_9[3]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_9_18[3]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_6, E => \DES_SM_1[6]_net_1\, Q
         => \BIT_OS_VAL_9[3]\);
    
    \REG40M.BIT_OS_VAL_0_RNO[0]\ : MX2
      port map(A => N_5666, B => \BIT_OS_VAL_0[0]\, S => N_5679, 
        Y => \N_BIT_OS_VAL_0_18[0]\);
    
    \CLKPHASE_RNIP0JI_3[1]\ : NOR2B
      port map(A => N_5712, B => N_204, Y => 
        \un36_n_bit_os_val[12]\);
    
    \REG40M.SEQCNTS_16[2]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[2]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_5, E => N_314, Q => \SEQCNTS_16[2]\);
    
    \REG40M.BIT_OS_CNT_2_RNI18OB[2]\ : NOR2B
      port map(A => BIT_OS_CNT_2_c1, B => \BIT_OS_CNT_2[2]\, Y
         => BIT_OS_CNT_2_c2);
    
    \ARB_BYTE_RNIALHJ2[1]\ : AO1
      port map(A => BIT_OS_CNT_7lde_0_a3_1, B => 
        BIT_OS_CNT_7lde_0_a3_0, C => N_4530, Y => BIT_OS_CNT_7e);
    
    \REG40M.SEQCNTS_23_RNIUGAH[3]\ : MX2
      port map(A => \SEQCNTS_23[3]\, B => \SEQCNTS_24[3]\, S => 
        \INDEX_CNT_0[0]_net_1\, Y => N_4121);
    
    \DES_SM_0_RNIII0V_0[8]\ : OR2
      port map(A => \DES_SM_0[8]_net_1\, B => \DES_SM_0[6]_net_1\, 
        Y => N_4530_0);
    
    \MAX_CNT[1]\ : DFN1E0C0
      port map(D => N_103, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_16, E => N_558, Q => \MAX_CNT[1]_net_1\);
    
    \REG40M.BIT_OS_VAL_1_RNIRUGO[0]\ : MX2
      port map(A => \BIT_OS_VAL_1[0]\, B => \BIT_OS_VAL_17[0]\, S
         => \CLKPHASE_0[4]_net_1\, Y => N_3627);
    
    \REG40M.BIT_OS_CNT_0_RNID13C[6]\ : OR2A
      port map(A => \BIT_OS_CNT_0[6]\, B => N_390, Y => N_404);
    
    \BEST_BIT_OS_VAL_RNO_9[2]\ : MX2
      port map(A => N_3908, B => N_3912, S => 
        \INDEX_CNT[3]_net_1\, Y => N_3916);
    
    \DES_SM_RNIK7A3A[8]\ : NOR2
      port map(A => \un39_n_seqcnts[0]\, B => \DES_SM[8]_net_1\, 
        Y => \N_SEQCNTS_1[0]\);
    
    \CLKPHASE_1_RNI16F92[2]\ : MX2
      port map(A => N_3735, B => N_3750, S => 
        \CLKPHASE_1[2]_net_1\, Y => N_3755);
    
    \BIT_OS_SEL[2]\ : DFN1C0
      port map(D => \BEST_BIT_OS_VAL[2]_net_1\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_27_1, Q => \BIT_OS_SEL[2]_net_1\);
    
    \REG40M.BIT_OS_CNT_0[8]\ : DFN1E1C0
      port map(D => N_107, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_3, E => BIT_OS_CNT_0e, Q => 
        \BIT_OS_CNT_0[8]\);
    
    \CLKPHASE_0_RNIB8JF2[2]\ : MX2
      port map(A => N_3668, B => N_3680, S => 
        \CLKPHASE_0[2]_net_1\, Y => N_3684);
    
    \ADJ_Q[10]\ : DFN1C0
      port map(D => \ADJ_Q[8]_net_1\, CLK => CCC_160M_ADJ, CLR
         => P_MASTER_POR_B_c_26, Q => \ADJ_Q[10]_net_1\);
    
    \REG40M.BIT_OS_VAL_24_RNO[2]\ : MX2
      port map(A => \BIT_OS_VAL_24[2]\, B => N_781_0, S => 
        \un36_n_bit_os_val[7]\, Y => N_173);
    
    \BEST_BIT_OS_VAL_RNO_17[1]\ : MX2
      port map(A => \BIT_OS_VAL_5[1]\, B => \BIT_OS_VAL_6[1]\, S
         => \INDEX_CNT_1[0]_net_1\, Y => N_3891);
    
    \RECD_SER_WORD_RNO_1[2]\ : AO1
      port map(A => n_recd_ser_word168, B => \ARB_BYTE[6]_net_1\, 
        C => \ARB_BYTE_m_1[7]\, Y => \N_RECD_SER_WORD_iv_0[2]\);
    
    \REG40M.BIT_OS_VAL_29[2]\ : DFN1E1C0
      port map(D => N_163, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_4, E => \DES_SM_1[6]_net_1\, Q => 
        \BIT_OS_VAL_29[2]\);
    
    \REG40M.BIT_OS_VAL_1[1]\ : DFN1E1C0
      port map(D => N_5661, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_17, E => \DES_SM_3[6]_net_1\, Q => 
        \BIT_OS_VAL_1[1]\);
    
    \REG40M.BIT_OS_VAL_16[3]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_16_18[3]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_16_0, E => \DES_SM_3[6]_net_1\, Q
         => \BIT_OS_VAL_16[3]\);
    
    \MAX_CNT[7]\ : DFN1E0C0
      port map(D => N_5633, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_16, E => N_558, Q => \MAX_CNT[7]_net_1\);
    
    \BIT_OS_SEL[1]\ : DFN1C0
      port map(D => \BEST_BIT_OS_VAL[1]_net_1\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_27_1, Q => \BIT_OS_SEL[1]_net_1\);
    
    un41_n_seqcnts_I_9 : XOR2
      port map(A => N_3_1, B => \un39_n_seqcnts[3]\, Y => I_9);
    
    \CLKPHASE_0_RNI87AF[1]\ : OR3
      port map(A => N_5663, B => N_5668, C => 
        \CLKPHASE_0[1]_net_1\, Y => N_5676);
    
    \REG40M.SEQCNTS_31[3]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[3]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_10, E => N_284, Q => \SEQCNTS_31[3]\);
    
    \REG40M.BIT_OS_CNT_4_RNO[7]\ : XA1C
      port map(A => \BIT_OS_CNT_4[7]\, B => N_410, C => N_4530_0, 
        Y => N_5620);
    
    \REG40M.BIT_OS_CNT_3[7]\ : DFN1E1C0
      port map(D => BIT_OS_CNT_3_n7, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_7, E => BIT_OS_CNT_3e, Q => 
        \BIT_OS_CNT_3[7]\);
    
    \DES_SM_RNO[3]\ : AOI1
      port map(A => \DES_SM_ns_i_a2_0_0_a3_0_1[5]\, B => N_116, C
         => N_5813, Y => \DES_SM_RNO[3]_net_1\);
    
    \INDEX_CNT_2_RNI79CJ1[3]\ : MX2
      port map(A => N_4016, B => N_4021, S => 
        \INDEX_CNT_2[3]_net_1\, Y => N_4026);
    
    \REG40M.BIT_OS_CNT_5[1]\ : DFN1E1C0
      port map(D => N_5631, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_11, E => BIT_OS_CNT_5e, Q => 
        \BIT_OS_CNT_5[1]\);
    
    \REG40M.BIT_OS_CNT_0_RNIRL55[2]\ : OR2A
      port map(A => \BIT_OS_CNT_0[2]\, B => N_368, Y => N_372);
    
    \REG40M.BIT_OS_VAL_17[0]\ : DFN1E1C0
      port map(D => N_252, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_18, E => \DES_SM_3[6]_net_1\, Q => 
        \BIT_OS_VAL_17[0]\);
    
    \REG40M.BIT_OS_VAL_0_RNO[3]\ : MX2
      port map(A => N_209_0, B => \BIT_OS_VAL_0[3]\, S => N_5679, 
        Y => \N_BIT_OS_VAL_0_18[3]\);
    
    \CLKPHASE_0_RNIDOEH4[1]\ : MX2
      port map(A => N_3753, B => N_3788, S => 
        \CLKPHASE_0[1]_net_1\, Y => N_3793);
    
    \REG40M.SEQCNTS_25_RNI773P[2]\ : MX2
      port map(A => \SEQCNTS_9[2]\, B => \SEQCNTS_25[2]\, S => 
        \CLKPHASE_3[4]_net_1\, Y => N_3765);
    
    \REG40M.BIT_OS_VAL_28_RNO[0]\ : MX2
      port map(A => \BIT_OS_VAL_28[0]\, B => N_5666, S => 
        \un36_n_bit_os_val[3]\, Y => N_219);
    
    \REG40M.SEQCNTS_27[4]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[4]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_13, E => N_292, Q => \SEQCNTS_27[4]\);
    
    \RECD_SER_WORD[4]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[4]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_30, Q => \RECD_SER_WORD[4]_net_1\);
    
    \REG40M.BIT_OS_VAL_25_RNO[0]\ : MX2
      port map(A => \BIT_OS_VAL_25[0]\, B => N_5666, S => 
        \un36_n_bit_os_val[6]\, Y => N_228);
    
    \REG40M.BIT_OS_VAL_15_RNIL33S[3]\ : MX2
      port map(A => \BIT_OS_VAL_31[3]\, B => \BIT_OS_VAL_15[3]\, 
        S => \CLKPHASE_3[4]_net_1\, Y => N_3602);
    
    \REG40M.SEQCNTS_2[4]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[4]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_10, E => N_342, Q => \SEQCNTS_2[4]\);
    
    \CLKPHASE_0_RNI8OS43[2]\ : MX2
      port map(A => N_3609, B => N_3621, S => 
        \CLKPHASE_0[2]_net_1\, Y => N_3625);
    
    \REG40M.BIT_OS_CNT_7_RNO[6]\ : XA1B
      port map(A => BIT_OS_CNT_7_c5, B => \BIT_OS_CNT_7[6]\, C
         => N_4530_2, Y => BIT_OS_CNT_7_n6);
    
    \BIT_OS_SEL_0[2]\ : DFN1C0
      port map(D => \BEST_BIT_OS_VAL[2]_net_1\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_27_1, Q => BIT_OS_SEL_0(2));
    
    \BEST_BIT_OS_VAL_RNO[2]\ : NOR2A
      port map(A => \N_BEST_BIT_OS_VAL_3[2]\, B => 
        \DES_SM[8]_net_1\, Y => \N_BEST_BIT_OS_VAL[2]\);
    
    \REG40M.SEQCNTS_28_RNIOHCT[4]\ : MX2
      port map(A => \SEQCNTS_12[4]\, B => \SEQCNTS_28[4]\, S => 
        \CLKPHASE_3[4]_net_1\, Y => N_3822);
    
    \REG40M.BIT_OS_VAL_13[2]\ : DFN1E1C0
      port map(D => N_193, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_12, E => \DES_SM_2[6]_net_1\, Q => 
        \BIT_OS_VAL_13[2]\);
    
    \REG40M.BIT_OS_CNT_3_RNO_0[4]\ : AX1C
      port map(A => \BIT_OS_CNT_3[3]\, B => BIT_OS_CNT_3_c2, C
         => \BIT_OS_CNT_3[4]\, Y => BIT_OS_CNT_3_n4_tz);
    
    \MAX_CNT_RNIOFHN1[4]\ : NOR3A
      port map(A => DES_SM_tr2_i_a3_4, B => \MAX_CNT[6]_net_1\, C
         => \MAX_CNT[4]_net_1\, Y => DES_SM_tr2_i_a3_6);
    
    \Q[3]\ : DFN1C0
      port map(D => \ADJ_Q[3]_net_1\, CLK => CCC_160M_FXD, CLR
         => P_MASTER_POR_B_c_34, Q => \Q[3]_net_1\);
    
    \INDEX_CNT_RNI3M821[1]\ : OR3B
      port map(A => \INDEX_CNT[4]_net_1\, B => 
        \INDEX_CNT[2]_net_1\, C => \INDEX_CNT[1]_net_1\, Y => 
        DES_SM_tr8_i_o2_1);
    
    \CLKPHASE_2_RNIS9FE1[3]\ : MX2
      port map(A => N_3629, B => N_3633, S => 
        \CLKPHASE_2[3]_net_1\, Y => N_3637);
    
    \DES_SM_0_RNIAB7UH7[8]\ : AO1A
      port map(A => N_5677, B => N_782_0, C => N_717_0, Y => 
        N_334);
    
    \CLKPHASE_RNIG15B_0[3]\ : NOR3B
      port map(A => \CLKPHASE[3]_net_1\, B => \CLKPHASE[4]_net_1\, 
        C => \CLKPHASE[0]_net_1\, Y => N_211);
    
    \REG40M.SEQCNTS_22_RNI5TMK[3]\ : MX2
      port map(A => \SEQCNTS_6[3]\, B => \SEQCNTS_22[3]\, S => 
        \CLKPHASE_5[4]_net_1\, Y => N_3851);
    
    \REG40M.SEQCNTS_15_RNIUIAD[2]\ : MX2
      port map(A => \SEQCNTS_15[2]\, B => \SEQCNTS_16[2]\, S => 
        \INDEX_CNT_0[0]_net_1\, Y => N_4090);
    
    \BEST_BIT_OS_VAL_RNO_18[1]\ : MX2
      port map(A => \BIT_OS_VAL_13[1]\, B => \BIT_OS_VAL_14[1]\, 
        S => \INDEX_CNT_2[0]_net_1\, Y => N_3895);
    
    \REG40M.BIT_OS_CNT_2_RNIRBER[6]\ : NOR2B
      port map(A => BIT_OS_CNT_2_c5, B => \BIT_OS_CNT_2[6]\, Y
         => BIT_OS_CNT_2_c6);
    
    \REG40M.BIT_OS_CNT_0[1]\ : DFN1E1C0
      port map(D => N_121, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_2, E => BIT_OS_CNT_0e, Q => 
        \BIT_OS_CNT_0[1]\);
    
    \ARB_WRD_40M_FIXED[10]\ : DFN1C0
      port map(D => \Q[10]_net_1\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_28, Q => \ARB_WRD_40M_FIXED[10]_net_1\);
    
    \BEST_BIT_OS_VAL_RNO_12[0]\ : MX2
      port map(A => N_3946, B => N_3950, S => 
        \INDEX_CNT_0[3]_net_1\, Y => N_3954);
    
    \REG40M.SEQCNTS_31[1]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[1]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_10, E => N_284, Q => \SEQCNTS_31[1]\);
    
    \RECD_SER_WORD_RNO[3]\ : OR3
      port map(A => \N_RECD_SER_WORD_iv_1[3]\, B => 
        \N_RECD_SER_WORD_iv_0[3]\, C => \N_RECD_SER_WORD_iv_5[3]\, 
        Y => \N_RECD_SER_WORD[3]\);
    
    \CLKPHASE_1_RNIHLE92[2]\ : MX2
      port map(A => N_3733, B => N_3748, S => 
        \CLKPHASE_1[2]_net_1\, Y => N_3753);
    
    \MAX_CNT[4]\ : DFN1E0C0
      port map(D => N_5636, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_16, E => N_558, Q => \MAX_CNT[4]_net_1\);
    
    \BEST_BIT_OS_VAL_RNO_17[3]\ : MX2
      port map(A => \BIT_OS_VAL_5[3]\, B => \BIT_OS_VAL_6[3]\, S
         => \INDEX_CNT_2[0]_net_1\, Y => N_3893);
    
    \WAITCNT[5]\ : DFN1E0C0
      port map(D => N_34, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_9, E => N_5790, Q => \WAITCNT[5]_net_1\);
    
    \Q[6]\ : DFN1C0
      port map(D => \ADJ_Q[6]_net_1\, CLK => CCC_160M_FXD, CLR
         => P_MASTER_POR_B_c_34, Q => \Q[6]_net_1\);
    
    \CLKPHASE_RNIPSLVG1[0]\ : NOR3C
      port map(A => N_762, B => \un107_bit_os_val[2]\, C => N_433, 
        Y => N_754);
    
    \REG40M.BIT_OS_VAL_17_RNO[1]\ : MX2B
      port map(A => \BIT_OS_VAL_17[1]\, B => N_206, S => 
        \un36_n_bit_os_val[14]\, Y => \N_BIT_OS_VAL_17_18[1]\);
    
    \REG40M.BIT_OS_VAL_26[0]\ : DFN1E1C0
      port map(D => N_225, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_21, E => \DES_SM[6]_net_1\, Q => 
        \BIT_OS_VAL_26[0]\);
    
    \REG40M.SEQCNTS_26[1]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[1]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_12, E => N_294, Q => \SEQCNTS_26[1]\);
    
    \REG40M.SEQCNTS_11[0]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[0]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_20, E => N_324, Q => \SEQCNTS_11[0]\);
    
    \Q[9]\ : DFN1C0
      port map(D => \ADJ_Q[9]_net_1\, CLK => CCC_160M_FXD, CLR
         => P_MASTER_POR_B_c_34, Q => \Q[9]_net_1\);
    
    \REG40M.BIT_OS_CNT_4[0]\ : DFN1E1C0
      port map(D => N_507, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_9, E => BIT_OS_CNT_4e, Q => 
        \BIT_OS_CNT_4[0]\);
    
    \CLKPHASE_0_RNIPHUQH7[1]\ : AO1
      port map(A => \un36_n_bit_os_val[22]\, B => N_782_0, C => 
        N_717_0, Y => N_328);
    
    \BEST_CLKPHASE[1]\ : DFN1E1C0
      port map(D => \N_BEST_CLKPHASE[1]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_10, E => un1_N_CCC_RESET_EN_0_sqmuxa, 
        Q => \BEST_CLKPHASE[1]_net_1\);
    
    \REG40M.BIT_OS_CNT_5[2]\ : DFN1E1C0
      port map(D => N_5630, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_11, E => BIT_OS_CNT_5e, Q => 
        \BIT_OS_CNT_5[2]\);
    
    \Q[5]\ : DFN1C0
      port map(D => \ADJ_Q[5]_net_1\, CLK => CCC_160M_FXD, CLR
         => P_MASTER_POR_B_c_34, Q => \Q[5]_net_1\);
    
    un3_n_index_cnt_I_7 : XOR2
      port map(A => N_4_0, B => \INDEX_CNT[2]_net_1\, Y => I_7_0);
    
    \REG40M.BIT_OS_VAL_7_RNI8R9J[3]\ : MX2
      port map(A => \BIT_OS_VAL_7[3]\, B => \BIT_OS_VAL_23[3]\, S
         => \CLKPHASE_4[4]_net_1\, Y => N_3606);
    
    \RECD_SER_WORD_RNO_3[5]\ : NOR3C
      port map(A => n_recd_ser_word167_1, B => 
        n_recd_ser_word171_0, C => \ARB_BYTE[12]_net_1\, Y => 
        \ARB_BYTE_m[12]\);
    
    \WAITCNT_RNO[1]\ : XA1B
      port map(A => \WAITCNT[0]_net_1\, B => \WAITCNT[1]_net_1\, 
        C => N_4539, Y => N_43);
    
    \REG40M.BIT_OS_VAL_8[3]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_8_18[3]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_5, E => \DES_SM_1[6]_net_1\, Q
         => \BIT_OS_VAL_8[3]\);
    
    \BIT_OS_SEL_3[2]\ : DFN1C0
      port map(D => \BEST_BIT_OS_VAL[2]_net_1\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_27_0, Q => BIT_OS_SEL_3(2));
    
    \REG40M.SEQCNTS_17_RNI0HAE[2]\ : MX2
      port map(A => \SEQCNTS_1[2]\, B => \SEQCNTS_17[2]\, S => 
        \CLKPHASE_3[4]_net_1\, Y => N_3760);
    
    \ARB_BYTE_RNICT161_1[1]\ : NOR3A
      port map(A => N_563_2, B => \ARB_BYTE[4]_net_1\, C => 
        \ARB_BYTE[1]_net_1\, Y => BIT_OS_CNT_4lde_0_a3_1);
    
    \REG40M.BIT_OS_CNT_5_RNIRBDE[0]\ : OR2B
      port map(A => \BIT_OS_CNT_5[1]\, B => \BIT_OS_CNT_5[0]\, Y
         => N_367);
    
    \RECD_SER_WORD_RNO_6[5]\ : OA1
      port map(A => \BIT_OS_SEL[3]_net_1\, B => 
        n_recd_ser_word164, C => \ARB_BYTE[5]_net_1\, Y => 
        \ARB_BYTE_m_4[5]\);
    
    \DES_SM_0_RNIII0V_1[8]\ : OR2
      port map(A => \DES_SM_0[8]_net_1\, B => \DES_SM_0[6]_net_1\, 
        Y => N_4530_1);
    
    \CLKPHASE_2_RNIEEBG1[3]\ : MX2
      port map(A => N_3816, B => N_3821, S => 
        \CLKPHASE_2[3]_net_1\, Y => N_3826);
    
    un1_CLKPHASE_I_1 : AND2
      port map(A => \CLKPHASE[0]_net_1\, B => 
        \DES_SM_RNIL6CU[5]_net_1\, Y => \DWACT_ADD_CI_0_TMP[0]\);
    
    \REG40M.BIT_OS_VAL_1[3]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_1_18[3]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_17_0, E => \DES_SM_3[6]_net_1\, Q
         => \BIT_OS_VAL_1[3]\);
    
    \BEST_BIT_OS_VAL_RNO_21[0]\ : MX2
      port map(A => \BIT_OS_VAL_21[0]\, B => \BIT_OS_VAL_22[0]\, 
        S => \INDEX_CNT[0]_net_1\, Y => N_3918);
    
    \REG40M.BIT_OS_VAL_7_RNO[1]\ : MX2B
      port map(A => \BIT_OS_VAL_7[1]\, B => N_206, S => 
        \un36_n_bit_os_val[24]\, Y => \N_BIT_OS_VAL_7_18[1]\);
    
    \REG40M.SEQCNTS_22[2]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[2]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_5, E => N_302, Q => \SEQCNTS_22[2]\);
    
    \ARB_BYTE[0]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[0]_net_1\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_27, Q => 
        \ARB_BYTE[0]_net_1\);
    
    \BEST_BIT_OS_VAL_RNO_18[2]\ : MX2
      port map(A => \BIT_OS_VAL_13[2]\, B => \BIT_OS_VAL_14[2]\, 
        S => \INDEX_CNT_2[0]_net_1\, Y => N_3896);
    
    \REG40M.BIT_OS_VAL_19_RNO[1]\ : MX2B
      port map(A => \BIT_OS_VAL_19[1]\, B => N_206, S => 
        \un36_n_bit_os_val[12]\, Y => \N_BIT_OS_VAL_19_18[1]\);
    
    \REG40M.SEQCNTS_7[2]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[2]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_17_0, E => N_332, Q => \SEQCNTS_7[2]\);
    
    \REG40M.BIT_OS_CNT_6_RNO_0[5]\ : OA1C
      port map(A => \BIT_OS_CNT_6[4]\, B => N_378, C => 
        \BIT_OS_CNT_6[5]\, Y => BIT_OS_CNT_6_n5_i_0);
    
    \REG40M.SEQCNTS_16_RNI6IH7[3]\ : NOR2B
      port map(A => \SEQCNTS_16[3]\, B => \CLKPHASE[4]_net_1\, Y
         => N_3801);
    
    \RECD_SER_WORD_RNO_8[4]\ : NOR3C
      port map(A => n_recd_ser_word165_2, B => 
        n_recd_ser_word167_1, C => \ARB_BYTE[7]_net_1\, Y => 
        \ARB_BYTE_m_3[7]\);
    
    \REG40M.BIT_OS_CNT_7_RNO[3]\ : XA1B
      port map(A => BIT_OS_CNT_7_c2, B => \BIT_OS_CNT_7[3]\, C
         => N_4530_2, Y => BIT_OS_CNT_7_n3);
    
    \ADJ_Q[8]\ : DFN1C0
      port map(D => \ADJ_Q[6]_net_1\, CLK => CCC_160M_ADJ, CLR
         => P_MASTER_POR_B_c_34_0, Q => \ADJ_Q[8]_net_1\);
    
    \REG40M.BIT_OS_VAL_7[1]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_7_18[1]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_3, E => \DES_SM_0[6]_net_1\, Q
         => \BIT_OS_VAL_7[1]\);
    
    \REG40M.BIT_OS_VAL_4_RNO[0]\ : MX2
      port map(A => N_5666_0, B => \BIT_OS_VAL_4[0]\, S => N_5674, 
        Y => \N_BIT_OS_VAL_4_18[0]\);
    
    \CLKPHASE_1_RNI195K1[3]\ : MX2
      port map(A => N_3687, B => N_3691, S => 
        \CLKPHASE_1[3]_net_1\, Y => N_3695);
    
    \REG40M.BIT_OS_VAL_5_RNI3G0G[2]\ : MX2
      port map(A => \BIT_OS_VAL_5[2]\, B => \BIT_OS_VAL_21[2]\, S
         => \CLKPHASE_5[4]_net_1\, Y => N_3641);
    
    \REG40M.BIT_OS_VAL_18_RNO[2]\ : MX2
      port map(A => \BIT_OS_VAL_18[2]\, B => N_781_0, S => 
        \un36_n_bit_os_val[13]\, Y => N_185);
    
    \REG40M.BIT_OS_CNT_2_RNO[4]\ : XA1B
      port map(A => BIT_OS_CNT_2_c3, B => \BIT_OS_CNT_2[4]\, C
         => N_4530_0, Y => BIT_OS_CNT_2_n4);
    
    \INDEX_CNT_RNIBLSEG[1]\ : MX2
      port map(A => N_4067, B => N_4142, S => 
        \INDEX_CNT[1]_net_1\, Y => \un6_n_best_seqcnt[4]\);
    
    \BEST_BIT_OS_VAL_RNO_16[1]\ : MX2
      port map(A => \BIT_OS_VAL_9[1]\, B => \BIT_OS_VAL_10[1]\, S
         => \INDEX_CNT_0[0]_net_1\, Y => N_3883);
    
    un41_n_seqcnts_I_11 : NOR2B
      port map(A => \un39_n_seqcnts[3]\, B => \DWACT_FINC_E[0]\, 
        Y => N_2);
    
    \REG40M.BIT_OS_VAL_27_RNO[1]\ : MX2B
      port map(A => \BIT_OS_VAL_27[1]\, B => N_206_0, S => 
        \un36_n_bit_os_val[4]\, Y => \N_BIT_OS_VAL_27_18[1]\);
    
    \INDEX_CNT_2_RNI35CJ1[3]\ : MX2
      port map(A => N_4015, B => N_4020, S => 
        \INDEX_CNT_2[3]_net_1\, Y => N_4025);
    
    \TUNE_CLKPHASE[1]\ : DFN1E1C0
      port map(D => \N_TUNE_CLKPHASE_2[1]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_12, E => \DES_SM[1]_net_1\, Q => 
        \TUNE_CLKPHASE[1]_net_1\);
    
    \RECD_SER_WORD_RNO_2[6]\ : OR3
      port map(A => \ARB_BYTE_m_4[8]\, B => \ARB_BYTE_m_5[6]\, C
         => \N_RECD_SER_WORD_iv_3[6]\, Y => 
        \N_RECD_SER_WORD_iv_5[6]\);
    
    \REG40M.BIT_OS_CNT_3[6]\ : DFN1E1C0
      port map(D => BIT_OS_CNT_3_n6, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_7, E => BIT_OS_CNT_3e, Q => 
        \BIT_OS_CNT_3[6]\);
    
    \RECD_SER_WORD_RNO_1[4]\ : AO1
      port map(A => \ARB_BYTE[8]_net_1\, B => n_recd_ser_word168, 
        C => \ARB_BYTE_m_1[9]\, Y => \N_RECD_SER_WORD_iv_0[4]\);
    
    \CLKPHASE_RNID3E7[3]\ : OR2
      port map(A => \CLKPHASE[3]_net_1\, B => \CLKPHASE[4]_net_1\, 
        Y => N_5663);
    
    \REG40M.BIT_OS_VAL_26[3]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_26_18[3]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_21, E => \DES_SM[6]_net_1\, Q => 
        \BIT_OS_VAL_26[3]\);
    
    \RECD_SER_WORD_RNO_0[7]\ : AO1
      port map(A => \ARB_BYTE[13]_net_1\, B => n_recd_ser_word170, 
        C => \ARB_BYTE_m[14]\, Y => \N_RECD_SER_WORD_iv_1[7]\);
    
    \CLKPHASE_0_RNIHE401[3]\ : MX2
      port map(A => N_3849, B => N_3854, S => 
        \CLKPHASE_0[3]_net_1\, Y => N_3859);
    
    \REG40M.BIT_OS_VAL_9_RNI6P9J[2]\ : MX2
      port map(A => \BIT_OS_VAL_9[2]\, B => \BIT_OS_VAL_25[2]\, S
         => \CLKPHASE_0[4]_net_1\, Y => N_3633);
    
    \REG40M.BIT_OS_VAL_3_RNO[1]\ : MX2A
      port map(A => N_206, B => \BIT_OS_VAL_3[1]\, S => N_5675, Y
         => N_5659);
    
    \DES_SM_1_RNIEL3O2[8]\ : NOR3B
      port map(A => N_5730, B => I_9_0, C => \DES_SM_1[8]_net_1\, 
        Y => \N_INDEX_CNT[3]\);
    
    \REG40M.BIT_OS_CNT_5_RNO[4]\ : XA1C
      port map(A => \BIT_OS_CNT_5[4]\, B => N_376, C => N_4530, Y
         => N_5628);
    
    \ARB_BYTE_RNI8S9F[3]\ : NOR2A
      port map(A => \ARB_BYTE[5]_net_1\, B => \ARB_BYTE[3]_net_1\, 
        Y => BIT_OS_CNT_3lde_0_a3_1);
    
    \BEST_BIT_OS_VAL_RNO_23[0]\ : MX2
      port map(A => \BIT_OS_VAL_11[0]\, B => \BIT_OS_VAL_12[0]\, 
        S => \INDEX_CNT_1[0]_net_1\, Y => N_3938);
    
    \RECD_SER_WORD_RNO_7[4]\ : AO1
      port map(A => n_recd_ser_word165, B => \ARB_BYTE[5]_net_1\, 
        C => \ARB_BYTE_m_3[7]\, Y => \N_RECD_SER_WORD_iv_3[4]\);
    
    \REG40M.BIT_OS_VAL_27[0]\ : DFN1E1C0
      port map(D => N_222, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_1, E => \DES_SM_0[6]_net_1\, Q => 
        \BIT_OS_VAL_27[0]\);
    
    \RECD_SER_WORD_RNO_3[6]\ : NOR3C
      port map(A => n_recd_ser_word167_1, B => 
        n_recd_ser_word171_0, C => \ARB_BYTE[13]_net_1\, Y => 
        \ARB_BYTE_m[13]\);
    
    \REG40M.SEQCNTS_8[4]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[4]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_19, E => N_330, Q => \SEQCNTS_8[4]\);
    
    \REG40M.BIT_OS_CNT_4[2]\ : DFN1E1C0
      port map(D => N_47, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_9, E => BIT_OS_CNT_4e, Q => 
        \BIT_OS_CNT_4[2]\);
    
    \CLKPHASE_0_RNIRDOR[3]\ : MX2
      port map(A => N_3723, B => N_3728, S => 
        \CLKPHASE_0[3]_net_1\, Y => N_3733);
    
    \WAITCNT[1]\ : DFN1E0C0
      port map(D => N_43, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_9, E => N_5790, Q => \WAITCNT[1]_net_1\);
    
    \REG40M.BIT_OS_CNT_7[3]\ : DFN1E1C0
      port map(D => BIT_OS_CNT_7_n3, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_14, E => BIT_OS_CNT_7e, Q => 
        \BIT_OS_CNT_7[3]\);
    
    \REG40M.SEQCNTS_28_RNIIBCT[1]\ : MX2
      port map(A => \SEQCNTS_12[1]\, B => \SEQCNTS_28[1]\, S => 
        \CLKPHASE_3[4]_net_1\, Y => N_3819);
    
    \REG40M.SEQCNTS_26[0]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[0]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_12, E => N_294, Q => \SEQCNTS_26[0]\);
    
    \REG40M.BIT_OS_VAL_18[2]\ : DFN1E1C0
      port map(D => N_185, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_19, E => \DES_SM_4[6]_net_1\, Q => 
        \BIT_OS_VAL_18[2]\);
    
    \REG40M.BIT_OS_CNT_6_RNO_0[7]\ : OA1C
      port map(A => \BIT_OS_CNT_6[6]\, B => N_387, C => 
        \BIT_OS_CNT_6[7]\, Y => BIT_OS_CNT_6_n7_i_0);
    
    \CLKPHASE_0_RNIE9411[3]\ : MX2
      port map(A => N_3640, B => N_3644, S => 
        \CLKPHASE_0[3]_net_1\, Y => N_3648);
    
    \ARB_BYTE[8]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[8]_net_1\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_27, Q => 
        \ARB_BYTE[8]_net_1\);
    
    \BIT_OS_SEL_5[1]\ : DFN1C0
      port map(D => \BEST_BIT_OS_VAL[1]_net_1\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_27_0, Q => BIT_OS_SEL_5(1));
    
    \WAITCNT_RNO[3]\ : XA1C
      port map(A => \WAITCNT[3]_net_1\, B => N_5773, C => N_4539, 
        Y => N_39);
    
    \WAITCNT[13]\ : DFN1E0C0
      port map(D => WAITCNT_n13, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_21, E => N_5790, Q => 
        \WAITCNT[13]_net_1\);
    
    \REG40M.BIT_OS_VAL_20_RNIQSGQ[0]\ : MX2
      port map(A => \BIT_OS_VAL_4[0]\, B => \BIT_OS_VAL_20[0]\, S
         => \CLKPHASE_2[4]_net_1\, Y => N_3671);
    
    \Q[2]\ : DFN1C0
      port map(D => \ADJ_Q[2]_net_1\, CLK => CCC_160M_FXD, CLR
         => P_MASTER_POR_B_c_34, Q => \Q[2]_net_1\);
    
    \BEST_BIT_OS_VAL_RNO_5[0]\ : MX2
      port map(A => N_3942, B => N_3954, S => 
        \INDEX_CNT_0[2]_net_1\, Y => N_3958);
    
    \REG40M.BIT_OS_VAL_29_RNO[1]\ : MX2B
      port map(A => \BIT_OS_VAL_29[1]\, B => N_206_0, S => 
        \un36_n_bit_os_val[2]\, Y => \N_BIT_OS_VAL_29_18[1]\);
    
    \RECD_SER_WORD_RNI31VH1[3]\ : NOR3B
      port map(A => \ELK_RX_SER_WORD_0[7]\, B => 
        \RECD_SER_WORD[3]_net_1\, C => \ELK_RX_SER_WORD_0[5]\, Y
         => ELK0_SYNC_DET_1_3);
    
    \REG40M.BIT_OS_VAL_23[2]\ : DFN1E1C0
      port map(D => N_5641, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_17_0, E => \DES_SM_3[6]_net_1\, Q => 
        \BIT_OS_VAL_23[2]\);
    
    \ARB_BYTE[5]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[5]_net_1\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_27, Q => 
        \ARB_BYTE[5]_net_1\);
    
    un3_n_index_cnt_I_9 : XOR2
      port map(A => N_3, B => \INDEX_CNT[3]_net_1\, Y => I_9_0);
    
    \REG40M.SEQCNTS_17[0]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[0]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_6, E => N_312, Q => \SEQCNTS_17[0]\);
    
    \REG40M.BIT_OS_CNT_6_RNO[6]\ : XA1C
      port map(A => N_387, B => \BIT_OS_CNT_6[6]\, C => N_4530_2, 
        Y => N_75);
    
    \CLKPHASE_0_RNIUSBJ5[1]\ : MX2
      port map(A => N_3683, B => N_3711, S => 
        \CLKPHASE_0[1]_net_1\, Y => N_3715);
    
    \REG40M.SEQCNTS_17_RNI6B3M[2]\ : MX2
      port map(A => \SEQCNTS_17[2]\, B => \SEQCNTS_18[2]\, S => 
        \INDEX_CNT_4[0]_net_1\, Y => N_4035);
    
    \DES_SM[1]\ : DFN1C0
      port map(D => \DES_SM_RNO[1]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_26, Q => \DES_SM[1]_net_1\);
    
    \CLKPHASE_0_RNIFHGK5[1]\ : MX2
      port map(A => N_3686, B => N_3714, S => 
        \CLKPHASE_0[1]_net_1\, Y => N_3718);
    
    \REG40M.BIT_OS_VAL_28_RNO[2]\ : MX2
      port map(A => \BIT_OS_VAL_28[2]\, B => N_781, S => 
        \un36_n_bit_os_val[3]\, Y => N_165);
    
    \CLKPHASE_RNID3E7_2[3]\ : NOR2A
      port map(A => \CLKPHASE[3]_net_1\, B => \CLKPHASE[4]_net_1\, 
        Y => N_5711);
    
    \REG40M.BIT_OS_VAL_6[2]\ : DFN1E1C0
      port map(D => N_5650, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_2, E => \DES_SM_0[6]_net_1\, Q => 
        \BIT_OS_VAL_6[2]\);
    
    \BEST_BIT_OS_VAL_RNO_23[1]\ : MX2
      port map(A => \BIT_OS_VAL_11[1]\, B => \BIT_OS_VAL_12[1]\, 
        S => \INDEX_CNT_1[0]_net_1\, Y => N_3939);
    
    \INDEX_CNT_2[3]\ : DFN1E0C0
      port map(D => \N_INDEX_CNT[3]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_17_0, E => N_5149, Q => 
        \INDEX_CNT_2[3]_net_1\);
    
    \REG40M.BIT_OS_VAL_8[1]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_8_18[1]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_5, E => \DES_SM_1[6]_net_1\, Q
         => \BIT_OS_VAL_8[1]\);
    
    \INDEX_CNT_RNIH4Q77[4]\ : MX2
      port map(A => N_4028, B => N_4058, S => 
        \INDEX_CNT[4]_net_1\, Y => N_4063);
    
    \DES_SM_RNO_2[2]\ : NOR2B
      port map(A => CCC_RX_CLK_LOCK, B => \WAITCNT[13]_net_1\, Y
         => \DES_SM_ns_0_i_0_a3_0_0[6]\);
    
    \REG40M.BIT_OS_CNT_6_RNIC0F22[7]\ : OR3B
      port map(A => \BIT_OS_CNT_6[6]\, B => \BIT_OS_CNT_6[7]\, C
         => N_387, Y => N_419);
    
    \INDEX_CNT_RNIJREH8[4]\ : MX2
      port map(A => N_4102, B => N_4137, S => 
        \INDEX_CNT[4]_net_1\, Y => N_4142);
    
    \WAITCNT[6]\ : DFN1E0C0
      port map(D => N_32, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_9, E => N_5790, Q => \WAITCNT[6]_net_1\);
    
    \REG40M.BIT_OS_CNT_1_RNICFJM[4]\ : OR3A
      port map(A => N_359, B => N_BIT_OS_VAL_316lto8_0_o3_2, C
         => N_BIT_OS_VAL_316lto8_0_o3_1, Y => N_BIT_OS_VAL_316);
    
    \INDEX_CNT_RNILMST1[3]\ : MX2
      port map(A => N_4107, B => N_4112, S => 
        \INDEX_CNT[3]_net_1\, Y => N_4117);
    
    \REG40M.BIT_OS_CNT_0_RNO[2]\ : XA1C
      port map(A => \BIT_OS_CNT_0[2]\, B => N_368, C => N_4530_2, 
        Y => N_119);
    
    \REG40M.SEQCNTS_24_RNI860O[3]\ : MX2
      port map(A => \SEQCNTS_8[3]\, B => \SEQCNTS_24[3]\, S => 
        \CLKPHASE_4[4]_net_1\, Y => N_3806);
    
    \CLKPHASE_1_RNIGC5U[3]\ : MX2
      port map(A => N_3777, B => N_3782, S => 
        \CLKPHASE_1[3]_net_1\, Y => N_3787);
    
    \REG40M.BIT_OS_CNT_1_RNO_0[3]\ : NOR2A
      port map(A => N_428, B => \BIT_OS_CNT_1[3]\, Y => N_554);
    
    \RECD_SER_WORD[2]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[2]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_29, Q => \RECD_SER_WORD[2]_net_1\);
    
    \CLKPHASE_RNICU2EH7_0[0]\ : AO1
      port map(A => \un36_n_bit_os_val[2]\, B => N_782, C => 
        N_717, Y => N_288);
    
    \REG40M.SEQCNTS_19[3]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[3]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_11, E => N_308, Q => \SEQCNTS_19[3]\);
    
    \REG40M.BIT_OS_VAL_1_RNO[0]\ : MX2
      port map(A => N_5666_0, B => \BIT_OS_VAL_1[0]\, S => N_5676, 
        Y => \N_BIT_OS_VAL_1_18[0]\);
    
    \REG40M.BIT_OS_CNT_3[1]\ : DFN1E1C0
      port map(D => BIT_OS_CNT_3_n1, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_7, E => BIT_OS_CNT_3e, Q => 
        \BIT_OS_CNT_3[1]\);
    
    \INDEX_CNT_RNICB083[2]\ : MX2
      port map(A => N_4045, B => N_4055, S => 
        \INDEX_CNT[2]_net_1\, Y => N_4060);
    
    \BEST_BIT_OS_VAL_RNO_26[0]\ : MX2
      port map(A => \BIT_OS_VAL_19[0]\, B => \BIT_OS_VAL_20[0]\, 
        S => \INDEX_CNT_1[0]_net_1\, Y => N_3962);
    
    \REG40M.BIT_OS_CNT_1_RNI12L5[8]\ : OR2
      port map(A => \BIT_OS_CNT_1[8]\, B => \BIT_OS_CNT_1[7]\, Y
         => N_BIT_OS_VAL_316lto8_0_o3_1);
    
    \REG40M.BIT_OS_VAL_0[3]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_0_18[3]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_15, E => \DES_SM_3[6]_net_1\, Q
         => \BIT_OS_VAL_0[3]\);
    
    \REG40M.BIT_OS_CNT_4_RNI9MPA1[6]\ : OR3B
      port map(A => \BIT_OS_CNT_4[5]\, B => \BIT_OS_CNT_4[6]\, C
         => N_382, Y => N_410);
    
    \PHASE_ADJ[4]\ : DFN1C0
      port map(D => \CLKPHASE[4]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c, Q => PHASE_ADJ_160_L(4));
    
    \BEST_BIT_OS_VAL_RNO_15[2]\ : MX2
      port map(A => \BIT_OS_VAL_1[2]\, B => \BIT_OS_VAL_2[2]\, S
         => \INDEX_CNT_0[0]_net_1\, Y => N_3880);
    
    \SYNC_SM.n_best_clkphase14_0_I_11\ : OA1
      port map(A => N_11, B => N_10, C => N_9, Y => 
        n_best_clkphase14);
    
    \REG40M.BIT_OS_VAL_13_RNO[3]\ : MX2
      port map(A => \BIT_OS_VAL_13[3]\, B => N_209, S => 
        \un36_n_bit_os_val[18]\, Y => \N_BIT_OS_VAL_13_18[3]\);
    
    \TUNE_CLKPHASE[2]\ : DFN1E1C0
      port map(D => \N_TUNE_CLKPHASE_2[2]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_12, E => \DES_SM[1]_net_1\, Q => 
        \TUNE_CLKPHASE[2]_net_1\);
    
    \SYNC_SM.n_best_clkphase14_0_I_2\ : OR2A
      port map(A => \BEST_SEQCNT[2]_net_1\, B => 
        \un6_n_best_seqcnt[2]\, Y => N_3_0);
    
    \REG40M.SEQCNTS_14[3]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[3]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_2, E => N_318, Q => \SEQCNTS_14[3]\);
    
    \REG40M.BIT_OS_CNT_2[3]\ : DFN1E1C0
      port map(D => BIT_OS_CNT_2_n3, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_5, E => BIT_OS_CNT_2e, Q => 
        \BIT_OS_CNT_2[3]\);
    
    \REG40M.SEQCNTS_17[1]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[1]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_7, E => N_312, Q => \SEQCNTS_17[1]\);
    
    \REG40M.BIT_OS_CNT_3_RNIHB3U[5]\ : NOR2B
      port map(A => BIT_OS_CNT_3_c4, B => \BIT_OS_CNT_3[5]\, Y
         => BIT_OS_CNT_3_c5);
    
    \REG40M.SEQCNTS_27_RNILUNU[2]\ : MX2
      port map(A => \SEQCNTS_27[2]\, B => \SEQCNTS_28[2]\, S => 
        \INDEX_CNT[0]_net_1\, Y => N_4110);
    
    \INDEX_CNT_RNID7BG2[3]\ : MX2
      port map(A => N_4070, B => N_4075, S => 
        \INDEX_CNT[3]_net_1\, Y => N_4080);
    
    \REG40M.SEQCNTS_24_RNI420O[1]\ : MX2
      port map(A => \SEQCNTS_8[1]\, B => \SEQCNTS_24[1]\, S => 
        \CLKPHASE_4[4]_net_1\, Y => N_3804);
    
    \REG40M.BIT_OS_VAL_6[1]\ : DFN1E1C0
      port map(D => N_5657, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_2, E => \DES_SM_0[6]_net_1\, Q => 
        \BIT_OS_VAL_6[1]\);
    
    \REG40M.BIT_OS_VAL_28_RNIHUV8[1]\ : MX2
      port map(A => \BIT_OS_VAL_12[1]\, B => \BIT_OS_VAL_28[1]\, 
        S => \CLKPHASE_0[4]_net_1\, Y => N_3676);
    
    \MAX_CNT_RNID37M[4]\ : NOR2
      port map(A => \MAX_CNT[5]_net_1\, B => \MAX_CNT[4]_net_1\, 
        Y => DES_SM_tr5_0_a3_2);
    
    \BIT_OS_SEL_1_RNII4DE1[0]\ : NOR3B
      port map(A => \BIT_OS_SEL_1[0]_net_1\, B => 
        n_recd_ser_word165_2, C => \BIT_OS_SEL_1[1]_net_1\, Y => 
        n_recd_ser_word165);
    
    \REG40M.SEQCNTS_17_RNI2JAE[3]\ : MX2
      port map(A => \SEQCNTS_1[3]\, B => \SEQCNTS_17[3]\, S => 
        \CLKPHASE_3[4]_net_1\, Y => N_3761);
    
    \REG40M.BIT_OS_VAL_16_RNO[1]\ : MX2B
      port map(A => \BIT_OS_VAL_16[1]\, B => N_206_0, S => 
        \un36_n_bit_os_val[15]\, Y => \N_BIT_OS_VAL_16_18[1]\);
    
    \REG40M.BIT_OS_CNT_4_RNO[5]\ : XA1C
      port map(A => \BIT_OS_CNT_4[5]\, B => N_382, C => N_4530_0, 
        Y => N_5622);
    
    \REG40M.BIT_OS_CNT_2_RNI16R7[6]\ : OR2
      port map(A => \BIT_OS_CNT_2[7]\, B => \BIT_OS_CNT_2[6]\, Y
         => N_BIT_OS_VAL_3110lto8_1);
    
    \BIT_OS_SEL_RNIPOQF[3]\ : NOR2
      port map(A => \BIT_OS_SEL[3]_net_1\, B => 
        \BIT_OS_SEL[0]_net_1\, Y => n_recd_ser_word170_0);
    
    un41_n_seqcnts_I_5 : XOR2
      port map(A => \un39_n_seqcnts[0]\, B => \un39_n_seqcnts[1]\, 
        Y => I_5);
    
    \DES_SM_4[6]\ : DFN1C0
      port map(D => N_MAX_CNT_0_sqmuxa, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_27_1, Q => \DES_SM_4[6]_net_1\);
    
    \CLKPHASE_0_RNIE8RD2[2]\ : MX2
      port map(A => N_3637, B => N_3649, S => 
        \CLKPHASE_0[2]_net_1\, Y => N_3653);
    
    \REG40M.BIT_OS_CNT_3_RNO[3]\ : XA1B
      port map(A => BIT_OS_CNT_3_c2, B => \BIT_OS_CNT_3[3]\, C
         => N_4530_1, Y => BIT_OS_CNT_3_n3);
    
    \PHASE_ADJ[2]\ : DFN1C0
      port map(D => \CLKPHASE[2]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c, Q => PHASE_ADJ_160_L(2));
    
    \DES_SM_RNIL6CU[5]\ : OR3A
      port map(A => \DES_SM_i_0[5]\, B => \DES_SM_0[8]_net_1\, C
         => \DES_SM[0]_net_1\, Y => \DES_SM_RNIL6CU[5]_net_1\);
    
    \REG40M.BIT_OS_CNT_4_RNIATAI[3]\ : OR3C
      port map(A => \BIT_OS_CNT_4[1]\, B => \BIT_OS_CNT_4[2]\, C
         => \BIT_OS_CNT_4[3]\, Y => N_363);
    
    \INDEX_CNT_1_RNIHG2O1[3]\ : MX2
      port map(A => N_4035, B => N_4040, S => 
        \INDEX_CNT_1[3]_net_1\, Y => N_4045);
    
    \CLKPHASE_2_RNI2EEB1[3]\ : MX2
      port map(A => N_3699, B => N_3703, S => 
        \CLKPHASE_2[3]_net_1\, Y => N_3707);
    
    \BEST_BIT_OS_VAL_RNO_26[2]\ : MX2
      port map(A => \BIT_OS_VAL_19[2]\, B => \BIT_OS_VAL_20[2]\, 
        S => \INDEX_CNT_1[0]_net_1\, Y => N_3964);
    
    \REG40M.SEQCNTS_4[3]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[3]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_13, E => N_338, Q => \SEQCNTS_4[3]\);
    
    \REG40M.BIT_OS_VAL_19[1]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_19_18[1]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_20, E => \DES_SM[6]_net_1\, Q => 
        \BIT_OS_VAL_19[1]\);
    
    \REG40M.BIT_OS_CNT_0_RNO[4]\ : XA1C
      port map(A => \BIT_OS_CNT_0[4]\, B => N_377, C => N_4530_2, 
        Y => N_5640);
    
    \REG40M.BIT_OS_VAL_23_RNO[3]\ : MX2
      port map(A => \BIT_OS_VAL_23[3]\, B => N_209_0, S => 
        \un36_n_bit_os_val[8]\, Y => \N_BIT_OS_VAL_23_18[3]\);
    
    \CLKPHASE_RNIAB7UH7_0[0]\ : AO1
      port map(A => \un36_n_bit_os_val[18]\, B => N_782_0, C => 
        N_717_0, Y => N_320);
    
    \REG40M.SEQCNTS_1_RNIJM9K[1]\ : MX2
      port map(A => \SEQCNTS_1[1]\, B => \SEQCNTS_2[1]\, S => 
        \INDEX_CNT_1[0]_net_1\, Y => N_3999);
    
    \REG40M.BIT_OS_CNT_5[8]\ : DFN1E1C0
      port map(D => N_53, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_11, E => BIT_OS_CNT_5e, Q => 
        \BIT_OS_CNT_5[8]\);
    
    \BIT_OS_SEL_RNIRQQF_0[3]\ : NOR2
      port map(A => \BIT_OS_SEL[3]_net_1\, B => 
        \BIT_OS_SEL[2]_net_1\, Y => n_recd_ser_word165_2);
    
    \REG40M.SEQCNTS_15_RNIGUS9[3]\ : MX2
      port map(A => \SEQCNTS_31[3]\, B => \SEQCNTS_15[3]\, S => 
        \CLKPHASE_0[4]_net_1\, Y => N_3726);
    
    \CLKPHASE_RNI9VD7[2]\ : OR2A
      port map(A => \CLKPHASE[2]_net_1\, B => \CLKPHASE[1]_net_1\, 
        Y => N_90);
    
    \REG40M.BIT_OS_VAL_30_RNIFPSP[1]\ : MX2
      port map(A => \BIT_OS_VAL_14[1]\, B => \BIT_OS_VAL_30[1]\, 
        S => \CLKPHASE_3[4]_net_1\, Y => N_3704);
    
    \REG40M.BIT_OS_CNT_5_RNO[8]\ : XA1C
      port map(A => \BIT_OS_CNT_5[8]\, B => N_421, C => N_4530, Y
         => N_53);
    
    \RECD_SER_WORD_RNO_8[0]\ : NOR3C
      port map(A => n_recd_ser_word165_2, B => 
        n_recd_ser_word167_1, C => \ARB_BYTE[3]_net_1\, Y => 
        \ARB_BYTE_m[3]\);
    
    \ADJ_Q[14]\ : DFN1C0
      port map(D => \ADJ_Q[12]_net_1\, CLK => CCC_160M_ADJ, CLR
         => P_MASTER_POR_B_c_26, Q => \ADJ_Q[14]_net_1\);
    
    \BEST_BIT_OS_VAL_RNO_0[3]\ : MX2
      port map(A => N_3933, B => N_3993, S => 
        \INDEX_CNT[1]_net_1\, Y => \N_BEST_BIT_OS_VAL_3[3]\);
    
    \REG40M.BIT_OS_VAL_28[2]\ : DFN1E1C0
      port map(D => N_165, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_2, E => \DES_SM_0[6]_net_1\, Q => 
        \BIT_OS_VAL_28[2]\);
    
    \RECD_SER_WORD_RNO_6[0]\ : OA1
      port map(A => \BIT_OS_SEL[3]_net_1\, B => 
        n_recd_ser_word164, C => \ARB_BYTE[0]_net_1\, Y => 
        \ARB_BYTE_m[0]\);
    
    \REG40M.BIT_OS_VAL_18[3]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_18_18[3]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_19, E => \DES_SM_4[6]_net_1\, Q
         => \BIT_OS_VAL_18[3]\);
    
    \INDEX_CNT_2_RNIFT9R1[3]\ : MX2
      port map(A => N_4083, B => N_4088, S => 
        \INDEX_CNT_2[3]_net_1\, Y => N_4093);
    
    \CLKPHASE_2_RNI89621[3]\ : MX2
      port map(A => N_3802, B => N_3807, S => 
        \CLKPHASE_2[3]_net_1\, Y => N_3812);
    
    \REG40M.BIT_OS_CNT_2_RNO[0]\ : NOR2
      port map(A => \BIT_OS_CNT_2[0]\, B => N_4530, Y => N_5610);
    
    \CLKPHASE_1_RNIHO5B1[3]\ : MX2
      port map(A => N_3659, B => N_3663, S => 
        \CLKPHASE_1[3]_net_1\, Y => N_3667);
    
    \INDEX_CNT_2_RNIN5AR1[3]\ : MX2
      port map(A => N_4085, B => N_4090, S => 
        \INDEX_CNT_2[3]_net_1\, Y => N_4095);
    
    \INDEX_CNT_RNIDEST1[3]\ : MX2
      port map(A => N_4105, B => N_4110, S => 
        \INDEX_CNT[3]_net_1\, Y => N_4115);
    
    \REG40M.BIT_OS_VAL_14[1]\ : DFN1E1C0
      port map(D => N_5656, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_13, E => \DES_SM_2[6]_net_1\, Q => 
        \BIT_OS_VAL_14[1]\);
    
    \REG40M.BIT_OS_CNT_4_RNO[4]\ : XA1C
      port map(A => \BIT_OS_CNT_4[4]\, B => N_379, C => N_4530_0, 
        Y => N_5623);
    
    \SYNC_SM.n_best_clkphase14_0_I_10\ : OA1A
      port map(A => N_6, B => N_8, C => N_7, Y => N_11);
    
    \REG40M.SEQCNTS_18_RNI7UJH[4]\ : MX2
      port map(A => \SEQCNTS_2[4]\, B => \SEQCNTS_18[4]\, S => 
        \CLKPHASE_4[4]_net_1\, Y => N_3837);
    
    \REG40M.BIT_OS_VAL_26_RNO[1]\ : MX2B
      port map(A => \BIT_OS_VAL_26[1]\, B => N_206, S => 
        \un36_n_bit_os_val[5]\, Y => \N_BIT_OS_VAL_26_18[1]\);
    
    \REG40M.BIT_OS_CNT_2_RNO[1]\ : XA1B
      port map(A => \BIT_OS_CNT_2[1]\, B => \BIT_OS_CNT_2[0]\, C
         => N_4530_0, Y => BIT_OS_CNT_2_n1);
    
    \REG40M.BIT_OS_CNT_6[1]\ : DFN1E1C0
      port map(D => N_85, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_12, E => BIT_OS_CNT_6e, Q => 
        \BIT_OS_CNT_6[1]\);
    
    \RECD_SER_WORD_RNO_8[7]\ : NOR3C
      port map(A => n_recd_ser_word165_2, B => 
        n_recd_ser_word167_1, C => \ARB_BYTE[10]_net_1\, Y => 
        \ARB_BYTE_m_3[10]\);
    
    \CLKPHASE_0_RNI3P0G2[2]\ : MX2
      port map(A => N_3845, B => N_3860, S => 
        \CLKPHASE_0[2]_net_1\, Y => N_3865);
    
    \REG40M.BIT_OS_CNT_2_RNI4BOB[1]\ : NOR3C
      port map(A => \BIT_OS_CNT_2[2]\, B => \BIT_OS_CNT_2[3]\, C
         => \BIT_OS_CNT_2[1]\, Y => N_BIT_OS_VAL_3110lt8);
    
    \ARB_BYTE[4]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[4]_net_1\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_27, Q => 
        \ARB_BYTE[4]_net_1\);
    
    \REG40M.SEQCNTS_23[4]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[4]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_6, E => N_300, Q => \SEQCNTS_23[4]\);
    
    \REG40M.SEQCNTS_3_RNISDVR[2]\ : MX2
      port map(A => \SEQCNTS_3[2]\, B => \SEQCNTS_4[2]\, S => 
        \INDEX_CNT_4[0]_net_1\, Y => N_4070);
    
    \REG40M.SEQCNTS_2[1]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[1]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_10, E => N_342, Q => \SEQCNTS_2[1]\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \SYNC_SM.n_best_clkphase14_0_I_1\ : OR2A
      port map(A => \un6_n_best_seqcnt[1]\, B => 
        \BEST_SEQCNT[1]_net_1\, Y => N_2_1);
    
    \REG40M.BIT_OS_CNT_6_RNI9UJG[7]\ : OR2
      port map(A => \BIT_OS_CNT_6[7]\, B => \BIT_OS_CNT_6[6]\, Y
         => N_354);
    
    \BEST_BIT_OS_VAL_RNO_10[1]\ : MX2
      port map(A => N_3919, B => \BIT_OS_VAL_29[1]\, S => 
        \INDEX_CNT[3]_net_1\, Y => N_3923);
    
    \REG40M.SEQCNTS_27_RNIL83Q[4]\ : MX2
      port map(A => \SEQCNTS_11[4]\, B => \SEQCNTS_27[4]\, S => 
        \CLKPHASE_2[4]_net_1\, Y => N_3747);
    
    \REG40M.BIT_OS_CNT_0_RNO[0]\ : NOR2
      port map(A => \BIT_OS_CNT_0[0]\, B => N_4530, Y => N_547);
    
    \CLKPHASE_RNIP0JI_9[0]\ : OR2A
      port map(A => N_5072_2, B => N_80, Y => N_5677);
    
    \REG40M.BIT_OS_VAL_1_RNO[3]\ : MX2
      port map(A => N_209, B => \BIT_OS_VAL_1[3]\, S => N_5676, Y
         => \N_BIT_OS_VAL_1_18[3]\);
    
    \INDEX_CNT_RNI2Q0A7[4]\ : MX2
      port map(A => N_4029, B => N_4059, S => 
        \INDEX_CNT[4]_net_1\, Y => N_4064);
    
    \REG40M.BIT_OS_CNT_1_RNI12F8[3]\ : OR3C
      port map(A => \BIT_OS_CNT_1[1]\, B => \BIT_OS_CNT_1[2]\, C
         => \BIT_OS_CNT_1[3]\, Y => N_359);
    
    \BEST_BIT_OS_VAL_RNO_24[1]\ : MX2
      port map(A => \BIT_OS_VAL_7[1]\, B => \BIT_OS_VAL_8[1]\, S
         => \INDEX_CNT_2[0]_net_1\, Y => N_3947);
    
    \REG40M.SEQCNTS_3_RNIUFVR[3]\ : MX2
      port map(A => \SEQCNTS_3[3]\, B => \SEQCNTS_4[3]\, S => 
        \INDEX_CNT_4[0]_net_1\, Y => N_4071);
    
    \WAITCNT[0]\ : DFN1E0C0
      port map(D => N_94, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_9, E => N_5790, Q => \WAITCNT[0]_net_1\);
    
    \REG40M.BIT_OS_VAL_0_RNI02EN[3]\ : MX2
      port map(A => \BIT_OS_VAL_0[3]\, B => \BIT_OS_VAL_16[3]\, S
         => \CLKPHASE_1[4]_net_1\, Y => N_3662);
    
    \RECD_SER_WORD_RNO_2[3]\ : OR3
      port map(A => \ARB_BYTE_m_2[5]\, B => \ARB_BYTE_m_2[3]\, C
         => \N_RECD_SER_WORD_iv_3[3]\, Y => 
        \N_RECD_SER_WORD_iv_5[3]\);
    
    \CLKPHASE_RNIVR8M2[2]\ : MX2
      port map(A => N_3812, B => N_3827, S => \CLKPHASE[2]_net_1\, 
        Y => N_3832);
    
    \DES_SM_RNICG0P1[0]\ : NOR3A
      port map(A => I_20, B => \DES_SM_1[8]_net_1\, C => 
        \DES_SM[0]_net_1\, Y => N_5796);
    
    \BIT_OS_SEL_RNIRQQF[3]\ : NOR2A
      port map(A => \BIT_OS_SEL[2]_net_1\, B => 
        \BIT_OS_SEL[3]_net_1\, Y => n_recd_ser_word171_0);
    
    \SYNC_SM.n_best_clkphase14_0_I_4\ : OR2A
      port map(A => \un6_n_best_seqcnt[4]\, B => 
        \BEST_SEQCNT[4]_net_1\, Y => N_5);
    
    \CLKPHASE_RNIV1AH1[3]\ : MX2
      port map(A => N_3612, B => N_3616, S => \CLKPHASE[3]_net_1\, 
        Y => N_3620);
    
    \REG40M.BIT_OS_VAL_9_RNI4N9J[1]\ : MX2
      port map(A => \BIT_OS_VAL_9[1]\, B => \BIT_OS_VAL_25[1]\, S
         => \CLKPHASE_0[4]_net_1\, Y => N_3632);
    
    \REG40M.SEQCNTS_12[1]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[1]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_21, E => N_322, Q => \SEQCNTS_12[1]\);
    
    \MAX_CNT_RNIKBHN1[4]\ : OR2A
      port map(A => \MAX_CNT[4]_net_1\, B => N_375, Y => N_385);
    
    \REG40M.BIT_OS_CNT_2_RNO[5]\ : XA1B
      port map(A => BIT_OS_CNT_2_c4, B => \BIT_OS_CNT_2[5]\, C
         => N_4530_0, Y => BIT_OS_CNT_2_n5);
    
    \REG40M.SEQCNTS_11[3]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[3]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_20, E => N_324, Q => \SEQCNTS_11[3]\);
    
    \CLKPHASE_RNI49DI1[3]\ : MX2
      port map(A => N_3613, B => N_3617, S => \CLKPHASE[3]_net_1\, 
        Y => N_3621);
    
    \REG40M.BIT_OS_VAL_7_RNI6P9J[2]\ : MX2
      port map(A => \BIT_OS_VAL_7[2]\, B => \BIT_OS_VAL_23[2]\, S
         => \CLKPHASE_4[4]_net_1\, Y => N_3605);
    
    \MAX_CNT_RNIGTDB3[4]\ : NOR3B
      port map(A => DES_SM_tr5_0_a3_3, B => DES_SM_tr5_0_a3_2, C
         => N_375, Y => N_MAX_CNT_0_sqmuxa);
    
    \INDEX_CNT_0_RNI65MN3[2]\ : MX2
      port map(A => N_4009, B => N_4024, S => 
        \INDEX_CNT_0[2]_net_1\, Y => N_4029);
    
    \BEST_CLKPHASE_RNO[4]\ : NOR2A
      port map(A => I_12_0, B => \DES_SM_1[8]_net_1\, Y => 
        \N_BEST_CLKPHASE[4]\);
    
    \REG40M.SEQCNTS_20_RNIVEAG[2]\ : MX2
      port map(A => \SEQCNTS_4[2]\, B => \SEQCNTS_20[2]\, S => 
        \CLKPHASE_5[4]_net_1\, Y => N_3815);
    
    \CLKPHASE_RNIDRVLE[0]\ : MX2
      port map(A => N_BIT_OS_VAL_3118, B => N_BIT_OS_VAL_3122, S
         => \un107_bit_os_val[0]\, Y => N_433);
    
    \CLKPHASE_4[4]\ : DFN1C0
      port map(D => \TUNE_CLKPHASE_RNITINS2[4]_net_1\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_24_0, Q => 
        \CLKPHASE_4[4]_net_1\);
    
    \BEST_BIT_OS_VAL_RNO_3[1]\ : MX2
      port map(A => N_3887, B => N_3899, S => 
        \INDEX_CNT_0[2]_net_1\, Y => N_3903);
    
    \REG40M.BIT_OS_CNT_2_RNIFMOB[8]\ : OR3
      port map(A => \BIT_OS_CNT_2[4]\, B => \BIT_OS_CNT_2[8]\, C
         => \BIT_OS_CNT_2[5]\, Y => N_BIT_OS_VAL_3110lto8_2);
    
    \CLKPHASE_0_RNIB11G2[2]\ : MX2
      port map(A => N_3846, B => N_3861, S => 
        \CLKPHASE_0[2]_net_1\, Y => N_3866);
    
    \MAX_CNT_RNO[8]\ : XA1C
      port map(A => \MAX_CNT[8]_net_1\, B => N_422, C => 
        un1_DES_SM_19, Y => N_89);
    
    \REG40M.BIT_OS_VAL_12[0]\ : DFN1E1C0
      port map(D => N_264, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_10, E => \DES_SM_1[6]_net_1\, Q => 
        \BIT_OS_VAL_12[0]\);
    
    \REG40M.BIT_OS_VAL_2_RNO[3]\ : MX2
      port map(A => N_209, B => \BIT_OS_VAL_2[3]\, S => N_5678, Y
         => \N_BIT_OS_VAL_2_18[3]\);
    
    \REG40M.BIT_OS_CNT_1_RNO_0[2]\ : AOI1
      port map(A => \BIT_OS_CNT_1[1]\, B => \BIT_OS_CNT_1[0]\, C
         => \BIT_OS_CNT_1[2]\, Y => N_555);
    
    \BEST_BIT_OS_VAL_RNO_15[1]\ : MX2
      port map(A => \BIT_OS_VAL_1[1]\, B => \BIT_OS_VAL_2[1]\, S
         => \INDEX_CNT_0[0]_net_1\, Y => N_3879);
    
    \WAITCNT_RNIU8DL[9]\ : NOR2
      port map(A => \WAITCNT[9]_net_1\, B => \WAITCNT[10]_net_1\, 
        Y => \DES_SM_ns_0_0_0_a2_1[0]\);
    
    \REG40M.BIT_OS_VAL_0_RNIQRDN[0]\ : MX2
      port map(A => \BIT_OS_VAL_0[0]\, B => \BIT_OS_VAL_16[0]\, S
         => \CLKPHASE_1[4]_net_1\, Y => N_3659);
    
    \WAITCNT_RNICVHC[2]\ : NOR2B
      port map(A => \WAITCNT[2]_net_1\, B => \WAITCNT[6]_net_1\, 
        Y => un1_DES_SM_471_i_0_a2_0_0_a2_2);
    
    \REG40M.BIT_OS_VAL_16[1]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_16_18[1]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_16_0, E => \DES_SM_3[6]_net_1\, Q
         => \BIT_OS_VAL_16[1]\);
    
    \CLKPHASE_0_RNIND1C_0[2]\ : NOR3A
      port map(A => \CLKPHASE_0[1]_net_1\, B => 
        \CLKPHASE_0[2]_net_1\, C => N_5672, Y => 
        \un36_n_bit_os_val[21]\);
    
    \CLKPHASE_RNO_0[0]\ : NOR3
      port map(A => \DES_SM_1[8]_net_1\, B => \DES_SM[0]_net_1\, 
        C => \DWACT_ADD_CI_0_partial_sum[0]\, Y => N_5797);
    
    \REG40M.BIT_OS_VAL_12_RNO[2]\ : MX2
      port map(A => \BIT_OS_VAL_12[2]\, B => N_781, S => 
        \un36_n_bit_os_val[19]\, Y => N_195);
    
    \REG40M.SEQCNTS_5[0]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[0]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_15, E => N_336, Q => \SEQCNTS_5[0]\);
    
    \REG40M.BIT_OS_VAL_28_RNIL209[3]\ : MX2
      port map(A => \BIT_OS_VAL_12[3]\, B => \BIT_OS_VAL_28[3]\, 
        S => \CLKPHASE_0[4]_net_1\, Y => N_3678);
    
    \REG40M.BIT_OS_CNT_2[4]\ : DFN1E1C0
      port map(D => BIT_OS_CNT_2_n4, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_5, E => BIT_OS_CNT_2e, Q => 
        \BIT_OS_CNT_2[4]\);
    
    \ADJ_Q[1]\ : DFN1C0
      port map(D => \ADJ_SER_IN_F_1DEL\, CLK => CCC_160M_ADJ, CLR
         => P_MASTER_POR_B_c_34_0, Q => \ADJ_Q[1]_net_1\);
    
    \REG40M.BIT_OS_VAL_11[0]\ : DFN1E1C0
      port map(D => N_267, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_8, E => \DES_SM_1[6]_net_1\, Q => 
        \BIT_OS_VAL_11[0]\);
    
    \RECD_SER_WORD_RNO_3[2]\ : NOR3C
      port map(A => n_recd_ser_word167_1, B => 
        n_recd_ser_word171_0, C => \ARB_BYTE[9]_net_1\, Y => 
        \ARB_BYTE_m[9]\);
    
    \RECD_SER_WORD_RNO_2[4]\ : OR3
      port map(A => \ARB_BYTE_m_3[6]\, B => \ARB_BYTE_m_3[4]\, C
         => \N_RECD_SER_WORD_iv_3[4]\, Y => 
        \N_RECD_SER_WORD_iv_5[4]\);
    
    \WAITCNT_RNO[0]\ : NOR2
      port map(A => \WAITCNT[0]_net_1\, B => N_4539, Y => N_94);
    
    \ARB_WRD_40M_FIXED[4]\ : DFN1C0
      port map(D => \Q[4]_net_1\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_26, Q => \ARB_WRD_40M_FIXED[4]_net_1\);
    
    \ARB_BYTE_RNI8GJU[1]\ : NOR3B
      port map(A => \ARB_BYTE[1]_net_1\, B => N_771, C => 
        \ARB_BYTE[4]_net_1\, Y => BIT_OS_CNT_0lde_0_a3_0);
    
    \REG40M.SEQCNTS_18_RNIVLJH[0]\ : MX2
      port map(A => \SEQCNTS_2[0]\, B => \SEQCNTS_18[0]\, S => 
        \CLKPHASE_4[4]_net_1\, Y => N_3833);
    
    \REG40M.BIT_OS_CNT_7[8]\ : DFN1E1C0
      port map(D => BIT_OS_CNT_7_n8, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_14, E => BIT_OS_CNT_7e, Q => 
        \BIT_OS_CNT_7[8]\);
    
    \DES_SM_RNI48SIB[6]\ : NOR2A
      port map(A => \DES_SM[6]_net_1\, B => \un107_bit_os_val[3]\, 
        Y => N_761);
    
    \REG40M.SEQCNTS_13[1]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[1]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_1, E => N_320, Q => \SEQCNTS_13[1]\);
    
    \RECD_SER_WORD_RNO_1[3]\ : AO1
      port map(A => n_recd_ser_word168, B => \ARB_BYTE[7]_net_1\, 
        C => \ARB_BYTE_m_1[8]\, Y => \N_RECD_SER_WORD_iv_0[3]\);
    
    \REG40M.BIT_OS_CNT_7_RNIS08B2[1]\ : OR3
      port map(A => N_BIT_OS_VAL_3130lt8, B => 
        N_BIT_OS_VAL_3130lto8_1, C => N_BIT_OS_VAL_3130lto8_2, Y
         => N_BIT_OS_VAL_3130);
    
    \RECD_SER_WORD_RNO_4[6]\ : NOR3C
      port map(A => n_recd_ser_word168_2, B => 
        n_recd_ser_word169_0, C => \ARB_BYTE[11]_net_1\, Y => 
        \ARB_BYTE_m_1[11]\);
    
    \WAITCNT_RNO[7]\ : XA1C
      port map(A => \WAITCNT[7]_net_1\, B => N_5777, C => N_4539, 
        Y => N_5719);
    
    \CLKPHASE_RNIP0JI_10[0]\ : OR2
      port map(A => N_80, B => N_90, Y => N_5674);
    
    \REG40M.BIT_OS_VAL_12_RNO[0]\ : MX2
      port map(A => \BIT_OS_VAL_12[0]\, B => N_5666, S => 
        \un36_n_bit_os_val[19]\, Y => N_264);
    
    \REG40M.BIT_OS_CNT_2_RNILPQ7[0]\ : NOR2B
      port map(A => \BIT_OS_CNT_2[0]\, B => \BIT_OS_CNT_2[1]\, Y
         => BIT_OS_CNT_2_c1);
    
    \INDEX_CNT_RNITIK4G[1]\ : MX2
      port map(A => N_4063, B => N_4138, S => 
        \INDEX_CNT[1]_net_1\, Y => \un6_n_best_seqcnt[0]\);
    
    \REG40M.SEQCNTS_11[1]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[1]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_20, E => N_324, Q => \SEQCNTS_11[1]\);
    
    \REG40M.BIT_OS_VAL_29[1]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_29_18[1]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_4, E => \DES_SM_1[6]_net_1\, Q
         => \BIT_OS_VAL_29[1]\);
    
    \WAITCNT_RNIAC8U[11]\ : NOR2
      port map(A => \WAITCNT[11]_net_1\, B => \WAITCNT[13]_net_1\, 
        Y => \DES_SM_ns_0_0_0_a2_2[0]\);
    
    \REG40M.SEQCNTS_17[3]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[3]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_7, E => N_312, Q => \SEQCNTS_17[3]\);
    
    \CLKPHASE_0_RNIBUOR[3]\ : MX2
      port map(A => N_3727, B => N_3732, S => 
        \CLKPHASE_0[3]_net_1\, Y => N_3737);
    
    \REG40M.BIT_OS_CNT_2_RNO[8]\ : XA1B
      port map(A => BIT_OS_CNT_2_260_0, B => \BIT_OS_CNT_2[8]\, C
         => N_4530_0, Y => BIT_OS_CNT_2_n8);
    
    \REG40M.SEQCNTS_20[0]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[0]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_2, E => N_306, Q => \SEQCNTS_20[0]\);
    
    \REG40M.SEQCNTS_17_RNI4LAE[4]\ : MX2
      port map(A => \SEQCNTS_1[4]\, B => \SEQCNTS_17[4]\, S => 
        \CLKPHASE_3[4]_net_1\, Y => N_3762);
    
    \REG40M.BIT_OS_VAL_20_RNISUGQ[1]\ : MX2
      port map(A => \BIT_OS_VAL_4[1]\, B => \BIT_OS_VAL_20[1]\, S
         => \CLKPHASE_2[4]_net_1\, Y => N_3672);
    
    \INDEX_CNT_RNO[1]\ : NOR3B
      port map(A => N_5730, B => I_5_0, C => \DES_SM_1[8]_net_1\, 
        Y => \N_INDEX_CNT[1]\);
    
    \REG40M.SEQCNTS_26_RNIH43Q[2]\ : MX2
      port map(A => \SEQCNTS_10[2]\, B => \SEQCNTS_26[2]\, S => 
        \CLKPHASE_4[4]_net_1\, Y => N_3840);
    
    \WAITCNT_RNI4KCV[4]\ : OR2A
      port map(A => \WAITCNT[4]_net_1\, B => N_5774, Y => N_5775);
    
    \WAITCNT_RNI8B2T2[11]\ : OR2A
      port map(A => \WAITCNT[11]_net_1\, B => N_5782, Y => N_5785);
    
    \REG40M.BIT_OS_VAL_9[0]\ : DFN1E1C0
      port map(D => N_273, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_6, E => \DES_SM_1[6]_net_1\, Q => 
        \BIT_OS_VAL_9[0]\);
    
    \REG40M.SEQCNTS_13[0]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[0]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_1, E => N_320, Q => \SEQCNTS_13[0]\);
    
    \REG40M.SEQCNTS_10_RNICTH31[2]\ : MX2
      port map(A => \SEQCNTS_9[2]\, B => \SEQCNTS_10[2]\, S => 
        \INDEX_CNT_1[0]_net_1\, Y => N_4005);
    
    \REG40M.BIT_OS_CNT_6[7]\ : DFN1E1C0
      port map(D => N_73, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_12, E => BIT_OS_CNT_6e, Q => 
        \BIT_OS_CNT_6[7]\);
    
    \DES_SM_0_RNIAB7UH7_0[8]\ : AO1A
      port map(A => N_5673, B => N_782_0, C => N_717_0, Y => 
        N_318);
    
    \CLKPHASE_0_RNIPM6J5[1]\ : MX2
      port map(A => N_3626, B => N_3654, S => 
        \CLKPHASE_0[1]_net_1\, Y => N_3658);
    
    \REG40M.BIT_OS_VAL_11_RNO[1]\ : MX2B
      port map(A => \BIT_OS_VAL_11[1]\, B => N_206_0, S => 
        \un36_n_bit_os_val[20]\, Y => \N_BIT_OS_VAL_11_18[1]\);
    
    \REG40M.SEQCNTS_28_RNIMFCT[3]\ : MX2
      port map(A => \SEQCNTS_12[3]\, B => \SEQCNTS_28[3]\, S => 
        \CLKPHASE_3[4]_net_1\, Y => N_3821);
    
    un3_n_index_cnt_I_10 : AND3
      port map(A => \INDEX_CNT_3[0]_net_1\, B => 
        \INDEX_CNT[1]_net_1\, C => \INDEX_CNT[2]_net_1\, Y => 
        \DWACT_FINC_E_0[0]\);
    
    \REG40M.BIT_OS_CNT_0_RNI00B4B_0[1]\ : NOR2A
      port map(A => N_BIT_OS_VAL_14_18_3_0_a2_1, B => N_781, Y
         => N_209);
    
    \INDEX_CNT_RNIHIST1[3]\ : MX2
      port map(A => N_4106, B => N_4111, S => 
        \INDEX_CNT[3]_net_1\, Y => N_4116);
    
    \BEST_SEQCNT[3]\ : DFN1E1C0
      port map(D => \N_BEST_SEQCNT[3]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_9, E => N_5724, Q => 
        \BEST_SEQCNT[3]_net_1\);
    
    \REG40M.BIT_OS_VAL_31_RNO[3]\ : MX2
      port map(A => \BIT_OS_VAL_31[3]\, B => N_209_0, S => 
        \un36_n_bit_os_val[0]\, Y => \N_BIT_OS_VAL_31_18[3]\);
    
    \REG40M.BIT_OS_VAL_19_RNO[0]\ : MX2
      port map(A => \BIT_OS_VAL_19[0]\, B => N_5666, S => 
        \un36_n_bit_os_val[12]\, Y => N_246);
    
    CONFIG_ONCE_TRIG : DFN1P0
      port map(D => N_58, CLK => CLK_40M_GL, PRE => 
        P_MASTER_POR_B_c_24, Q => CCC2_CONFIG_TRIG_i_0);
    
    \REG40M.BIT_OS_VAL_8[2]\ : DFN1E1C0
      port map(D => N_203, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_5, E => \DES_SM_1[6]_net_1\, Q => 
        \BIT_OS_VAL_8[2]\);
    
    \REG40M.BIT_OS_VAL_28[3]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_28_18[3]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_2, E => \DES_SM_0[6]_net_1\, Q
         => \BIT_OS_VAL_28[3]\);
    
    \REG40M.BIT_OS_CNT_0[6]\ : DFN1E1C0
      port map(D => N_111, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_3, E => BIT_OS_CNT_0e, Q => 
        \BIT_OS_CNT_0[6]\);
    
    \WAITCNT_RNIV9DL[8]\ : NOR2B
      port map(A => \WAITCNT[12]_net_1\, B => \WAITCNT[8]_net_1\, 
        Y => un1_DES_SM_471_i_0_a2_0_0_a2_4);
    
    \REG40M.SEQCNTS_10_RNIG1I31[4]\ : MX2
      port map(A => \SEQCNTS_9[4]\, B => \SEQCNTS_10[4]\, S => 
        \INDEX_CNT_1[0]_net_1\, Y => N_4007);
    
    \REG40M.BIT_OS_CNT_5_RNO[6]\ : NOR3A
      port map(A => N_409, B => N_4530, C => N_511, Y => N_5626);
    
    \ARB_BYTE_RNIALHJ2_0[1]\ : AO1
      port map(A => BIT_OS_CNT_2lde_0_a3_1, B => N_561_3, C => 
        N_4530, Y => BIT_OS_CNT_2e);
    
    \REG40M.BIT_OS_VAL_4_RNO[1]\ : MX2A
      port map(A => N_206_0, B => \BIT_OS_VAL_4[1]\, S => N_5674, 
        Y => N_5658);
    
    \REG40M.SEQCNTS_26_RNIL83Q[4]\ : MX2
      port map(A => \SEQCNTS_10[4]\, B => \SEQCNTS_26[4]\, S => 
        \CLKPHASE_4[4]_net_1\, Y => N_3842);
    
    \RECD_SER_WORD_RNO_5[6]\ : NOR3C
      port map(A => n_recd_ser_word165_2, B => 
        n_recd_ser_word166_0, C => \ARB_BYTE[8]_net_1\, Y => 
        \ARB_BYTE_m_4[8]\);
    
    \REG40M.BIT_OS_CNT_1[2]\ : DFN1E1C0
      port map(D => N_137, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_4, E => BIT_OS_CNT_1e, Q => 
        \BIT_OS_CNT_1[2]\);
    
    \REG40M.BIT_OS_VAL_24[1]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_24_18[1]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_18, E => \DES_SM_4[6]_net_1\, Q
         => \BIT_OS_VAL_24[1]\);
    
    \REG40M.BIT_OS_VAL_12_RNO[1]\ : MX2B
      port map(A => \BIT_OS_VAL_12[1]\, B => N_206_0, S => 
        \un36_n_bit_os_val[19]\, Y => \N_BIT_OS_VAL_12_18[1]\);
    
    \CLKPHASE_2_RNI0EFE1[3]\ : MX2
      port map(A => N_3630, B => N_3634, S => 
        \CLKPHASE_2[3]_net_1\, Y => N_3638);
    
    \REG40M.SEQCNTS_12[3]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[3]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_21, E => N_322, Q => \SEQCNTS_12[3]\);
    
    \REG40M.BIT_OS_VAL_22_RNO[2]\ : MX2
      port map(A => \BIT_OS_VAL_22[2]\, B => N_781_0, S => 
        \un36_n_bit_os_val[9]\, Y => N_177);
    
    \REG40M.SEQCNTS_17_RNIAF3M[4]\ : MX2
      port map(A => \SEQCNTS_17[4]\, B => \SEQCNTS_18[4]\, S => 
        \INDEX_CNT_4[0]_net_1\, Y => N_4037);
    
    \REG40M.BIT_OS_VAL_9_RNO[0]\ : MX2
      port map(A => \BIT_OS_VAL_9[0]\, B => N_5666, S => 
        \un36_n_bit_os_val[22]\, Y => N_273);
    
    \CLKPHASE_0[4]\ : DFN1C0
      port map(D => \TUNE_CLKPHASE_RNITINS2[4]_net_1\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_24_0, Q => 
        \CLKPHASE_0[4]_net_1\);
    
    \CLKPHASE_1_RNI1U4C1[3]\ : MX2
      port map(A => N_3738, B => N_3743, S => 
        \CLKPHASE_1[3]_net_1\, Y => N_3748);
    
    \CLKPHASE_0_RNI87AF_0[1]\ : NOR3A
      port map(A => N_5711, B => \CLKPHASE_0[1]_net_1\, C => 
        N_5668, Y => \un36_n_bit_os_val[22]\);
    
    \BEST_BIT_OS_VAL_RNO_6[2]\ : MX2
      port map(A => N_3972, B => N_3984, S => 
        \INDEX_CNT[2]_net_1\, Y => N_3988);
    
    \REG40M.BIT_OS_VAL_31[3]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_31_18[3]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_20, E => \DES_SM[6]_net_1\, Q => 
        \BIT_OS_VAL_31[3]\);
    
    \MAX_CNT_RNO[0]\ : NOR2
      port map(A => \MAX_CNT[0]_net_1\, B => un1_DES_SM_19, Y => 
        N_537);
    
    \SYNC_SM.n_best_clkphase14_0_I_5\ : AO1C
      port map(A => \un6_n_best_seqcnt[1]\, B => 
        \BEST_SEQCNT[1]_net_1\, C => N_4_1, Y => N_6);
    
    \DES_SM_RNO_0[2]\ : AOI1B
      port map(A => OP_MODE_c_0, B => \DES_SM_0[8]_net_1\, C => 
        \DES_SM_ns_0_i_0_a3_0_0[6]\, Y => 
        \DES_SM_ns_0_i_0_a3_0_1[6]\);
    
    \DES_SM_RNI1EH11_0[0]\ : AOI1
      port map(A => N_5783, B => CCC_RX_CLK_LOCK, C => 
        \DES_SM[0]_net_1\, Y => un1_DES_SM_471_i_0_0_0_0);
    
    \REG40M.BIT_OS_CNT_1_RNIAB9B[0]\ : OR2A
      port map(A => \BIT_OS_CNT_1[0]\, B => N_359, Y => N_380);
    
    \CLKPHASE_3[4]\ : DFN1C0
      port map(D => \TUNE_CLKPHASE_RNITINS2[4]_net_1\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_24_0, Q => 
        \CLKPHASE_3[4]_net_1\);
    
    \PHASE_ADJ[3]\ : DFN1C0
      port map(D => \CLKPHASE[3]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c, Q => PHASE_ADJ_160_L(3));
    
    \BEST_BIT_OS_VAL_RNO_28[3]\ : MX2
      port map(A => \BIT_OS_VAL_23[3]\, B => \BIT_OS_VAL_24[3]\, 
        S => \INDEX_CNT_2[0]_net_1\, Y => N_3977);
    
    \WAITCNT_RNO[11]\ : XA1C
      port map(A => \WAITCNT[11]_net_1\, B => N_5782, C => N_4539, 
        Y => N_5812);
    
    \REG40M.BIT_OS_VAL_22_RNO[0]\ : MX2
      port map(A => \BIT_OS_VAL_22[0]\, B => N_5666_0, S => 
        \un36_n_bit_os_val[9]\, Y => N_237);
    
    \MAX_CNT_RNIUAEC1[2]\ : NOR3B
      port map(A => \MAX_CNT[2]_net_1\, B => DES_SM_tr2_i_a3_2, C
         => \MAX_CNT[8]_net_1\, Y => DES_SM_tr2_i_a3_5);
    
    \CLKPHASE_1_RNISRMG2[2]\ : MX2
      port map(A => N_3670, B => N_3682, S => 
        \CLKPHASE_1[2]_net_1\, Y => N_3686);
    
    \INDEX_CNT_0_RNIN78A1[3]\ : MX2
      port map(A => N_4122, B => N_4127, S => 
        \INDEX_CNT_0[3]_net_1\, Y => N_4132);
    
    \CLKPHASE_0_RNIF0NJ4[1]\ : MX2
      port map(A => N_3757, B => N_3792, S => 
        \CLKPHASE_0[1]_net_1\, Y => N_3797);
    
    \REG40M.BIT_OS_VAL_9[1]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_9_18[1]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_6, E => \DES_SM_1[6]_net_1\, Q
         => \BIT_OS_VAL_9[1]\);
    
    \BEST_BIT_OS_VAL_RNO_26[3]\ : MX2
      port map(A => \BIT_OS_VAL_19[3]\, B => \BIT_OS_VAL_20[3]\, 
        S => \INDEX_CNT_1[0]_net_1\, Y => N_3965);
    
    \REG40M.BIT_OS_CNT_6[8]\ : DFN1E1C0
      port map(D => N_5632, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_12, E => BIT_OS_CNT_6e, Q => 
        \BIT_OS_CNT_6[8]\);
    
    \REG40M.SEQCNTS_21_RNI1D4E[4]\ : MX2
      port map(A => \SEQCNTS_5[4]\, B => \SEQCNTS_21[4]\, S => 
        \CLKPHASE_1[4]_net_1\, Y => N_3777);
    
    \CLKPHASE_0_RNIVCP33[2]\ : MX2
      port map(A => N_3608, B => N_3620, S => 
        \CLKPHASE_0[2]_net_1\, Y => N_3624);
    
    \REG40M.BIT_OS_CNT_7_RNIJO6S[1]\ : NOR3C
      port map(A => \BIT_OS_CNT_7[2]\, B => \BIT_OS_CNT_7[3]\, C
         => \BIT_OS_CNT_7[1]\, Y => N_BIT_OS_VAL_3130lt8);
    
    \REG40M.SEQCNTS_6[2]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[2]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_16, E => N_334, Q => \SEQCNTS_6[2]\);
    
    \REG40M.BIT_OS_VAL_21_RNO[1]\ : MX2B
      port map(A => \BIT_OS_VAL_21[1]\, B => N_206, S => 
        \un36_n_bit_os_val[10]\, Y => \N_BIT_OS_VAL_21_18[1]\);
    
    \REG40M.BIT_OS_CNT_6_RNIS8GMA[7]\ : AO1A
      port map(A => N_BIT_OS_VAL_3126, B => N_84, C => 
        N_BIT_OS_VAL_3130, Y => N_5666);
    
    \BEST_CLKPHASE[4]\ : DFN1E1C0
      port map(D => \N_BEST_CLKPHASE[4]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_10, E => un1_N_CCC_RESET_EN_0_sqmuxa, 
        Q => \BEST_CLKPHASE[4]_net_1\);
    
    \BEST_BIT_OS_VAL_RNO_2[1]\ : MX2
      port map(A => N_3959, B => N_3987, S => 
        \INDEX_CNT[4]_net_1\, Y => N_3991);
    
    \REG40M.BIT_OS_VAL_14_RNO[1]\ : MX2A
      port map(A => N_206_0, B => \BIT_OS_VAL_14[1]\, S => N_5673, 
        Y => N_5656);
    
    \REG40M.BIT_OS_VAL_29_RNO[0]\ : MX2
      port map(A => \BIT_OS_VAL_29[0]\, B => N_5666_0, S => 
        \un36_n_bit_os_val[2]\, Y => N_216);
    
    \REG40M.BIT_OS_VAL_0[2]\ : DFN1E1C0
      port map(D => N_5655, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_15, E => \DES_SM_3[6]_net_1\, Q => 
        \BIT_OS_VAL_0[2]\);
    
    \CLKPHASE_0_RNI25V31[3]\ : MX2
      port map(A => N_3672, B => N_3676, S => 
        \CLKPHASE_0[3]_net_1\, Y => N_3680);
    
    \DES_SM_RNICU2EH7_0[8]\ : AO1
      port map(A => \un36_n_bit_os_val[4]\, B => N_782, C => 
        N_717, Y => N_292);
    
    \ADJ_Q[2]\ : DFN1C0
      port map(D => \ADJ_Q[0]_net_1\, CLK => CCC_160M_ADJ, CLR
         => P_MASTER_POR_B_c_34_0, Q => \ADJ_Q[2]_net_1\);
    
    \MAX_CNT_RNO[1]\ : XA1B
      port map(A => \MAX_CNT[0]_net_1\, B => \MAX_CNT[1]_net_1\, 
        C => un1_DES_SM_19, Y => N_103);
    
    \ARB_WRD_40M_FIXED[0]\ : DFN1C0
      port map(D => \Q[0]_net_1\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_26, Q => \ARB_WRD_40M_FIXED[0]_net_1\);
    
    \REG40M.SEQCNTS_1[4]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[4]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_8, E => N_344, Q => \SEQCNTS_1[4]\);
    
    \REG40M.BIT_OS_VAL_22_RNO[1]\ : MX2B
      port map(A => \BIT_OS_VAL_22[1]\, B => N_206_0, S => 
        \un36_n_bit_os_val[9]\, Y => \N_BIT_OS_VAL_22_18[1]\);
    
    \REG40M.BIT_OS_VAL_22[0]\ : DFN1E1C0
      port map(D => N_237, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_15, E => \DES_SM_3[6]_net_1\, Q => 
        \BIT_OS_VAL_22[0]\);
    
    \REG40M.BIT_OS_VAL_18_RNO[3]\ : MX2
      port map(A => \BIT_OS_VAL_18[3]\, B => N_209, S => 
        \un36_n_bit_os_val[13]\, Y => \N_BIT_OS_VAL_18_18[3]\);
    
    \REG40M.BIT_OS_CNT_2_RNIGPSV9_0[1]\ : OA1C
      port map(A => N_445, B => N_437, C => N_360, Y => N_206_0);
    
    \REG40M.SEQCNTS_23_RNI0JAH[4]\ : MX2
      port map(A => \SEQCNTS_23[4]\, B => \SEQCNTS_24[4]\, S => 
        \INDEX_CNT_0[0]_net_1\, Y => N_4122);
    
    \REG40M.SEQCNTS_15_RNII0T9[4]\ : MX2
      port map(A => \SEQCNTS_31[4]\, B => \SEQCNTS_15[4]\, S => 
        \CLKPHASE_0[4]_net_1\, Y => N_3727);
    
    \INDEX_CNT_1[0]\ : DFN1E0C0
      port map(D => \N_INDEX_CNT[0]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_16_0, E => N_5149, Q => 
        \INDEX_CNT_1[0]_net_1\);
    
    \INDEX_CNT_0_RNILRSE3[2]\ : MX2
      port map(A => N_4113, B => N_4128, S => 
        \INDEX_CNT_0[2]_net_1\, Y => N_4133);
    
    \BEST_BIT_OS_VAL_RNO_27[1]\ : MX2
      port map(A => \BIT_OS_VAL_27[1]\, B => \BIT_OS_VAL_28[1]\, 
        S => \INDEX_CNT_1[0]_net_1\, Y => N_3967);
    
    \REG40M.BIT_OS_VAL_26[1]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_26_18[1]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_21, E => \DES_SM[6]_net_1\, Q => 
        \BIT_OS_VAL_26[1]\);
    
    \CLKPHASE_2_RNIAMEB1[3]\ : MX2
      port map(A => N_3701, B => N_3705, S => 
        \CLKPHASE_2[3]_net_1\, Y => N_3709);
    
    \Q[8]\ : DFN1C0
      port map(D => \ADJ_Q[8]_net_1\, CLK => CCC_160M_FXD, CLR
         => P_MASTER_POR_B_c_34, Q => \Q[8]_net_1\);
    
    \CLKPHASE_5[4]\ : DFN1C0
      port map(D => \TUNE_CLKPHASE_RNITINS2[4]_net_1\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_24_0, Q => 
        \CLKPHASE_5[4]_net_1\);
    
    \RECD_SER_WORD_RNO_7[5]\ : AO1
      port map(A => n_recd_ser_word165, B => \ARB_BYTE[6]_net_1\, 
        C => \ARB_BYTE_m_3[8]\, Y => \N_RECD_SER_WORD_iv_3[5]\);
    
    \REG40M.SEQCNTS_2[0]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[0]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_10, E => N_342, Q => \SEQCNTS_2[0]\);
    
    \CLKPHASE_0_RNIPHUQH7_0[1]\ : AO1A
      port map(A => N_5676, B => N_782_0, C => N_717_0, Y => 
        N_344);
    
    \BEST_BIT_OS_VAL_RNO_6[3]\ : MX2
      port map(A => N_3973, B => N_3985, S => 
        \INDEX_CNT[2]_net_1\, Y => N_3989);
    
    \WAITCNT_RNI6TGO1[8]\ : OR3B
      port map(A => \WAITCNT[7]_net_1\, B => \WAITCNT[8]_net_1\, 
        C => N_5777, Y => N_5779);
    
    \REG40M.BIT_OS_VAL_21[0]\ : DFN1E1C0
      port map(D => N_240, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_14, E => \DES_SM_2[6]_net_1\, Q => 
        \BIT_OS_VAL_21[0]\);
    
    \CLKPHASE_RNIP0JI_1[1]\ : NOR3A
      port map(A => N_204, B => \CLKPHASE[1]_net_1\, C => N_5668, 
        Y => \un36_n_bit_os_val[14]\);
    
    \REG40M.BIT_OS_CNT_7[4]\ : DFN1E1C0
      port map(D => BIT_OS_CNT_7_n4, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_14, E => BIT_OS_CNT_7e, Q => 
        \BIT_OS_CNT_7[4]\);
    
    \REG40M.BIT_OS_VAL_0[1]\ : DFN1E1C0
      port map(D => N_5662, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_15, E => \DES_SM_3[6]_net_1\, Q => 
        \BIT_OS_VAL_0[1]\);
    
    \REG40M.BIT_OS_CNT_5_RNO[7]\ : XA1C
      port map(A => \BIT_OS_CNT_5[7]\, B => N_409, C => N_4530, Y
         => N_5625);
    
    \BEST_BIT_OS_VAL_RNO_3[2]\ : MX2
      port map(A => N_3888, B => N_3900, S => 
        \INDEX_CNT_0[2]_net_1\, Y => N_3904);
    
    \INDEX_CNT_2[0]\ : DFN1E0C0
      port map(D => \N_INDEX_CNT[0]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_16_0, E => N_5149, Q => 
        \INDEX_CNT_2[0]_net_1\);
    
    \ADJ_Q[13]\ : DFN1C0
      port map(D => \ADJ_Q[11]_net_1\, CLK => CCC_160M_ADJ, CLR
         => P_MASTER_POR_B_c_26, Q => \ADJ_Q[13]_net_1\);
    
    \BEST_BIT_OS_VAL_RNO_13[3]\ : MX2
      port map(A => N_3965, B => N_3969, S => 
        \INDEX_CNT_1[3]_net_1\, Y => N_3973);
    
    \CLKPHASE_RNICU2EH7_0[2]\ : AO1
      port map(A => \un36_n_bit_os_val[7]\, B => N_782, C => 
        N_717, Y => N_298);
    
    \REG40M.SEQCNTS_13_RNIO84B[0]\ : MX2
      port map(A => \SEQCNTS_13[0]\, B => \SEQCNTS_14[0]\, S => 
        \INDEX_CNT_2[0]_net_1\, Y => N_4018);
    
    \REG40M.BIT_OS_CNT_2_RNIS7JJ[4]\ : NOR2B
      port map(A => BIT_OS_CNT_2_c3, B => \BIT_OS_CNT_2[4]\, Y
         => BIT_OS_CNT_2_c4);
    
    \CLKPHASE_0_RNIC89K5[1]\ : MX2
      port map(A => N_3624, B => N_3652, S => 
        \CLKPHASE_0[1]_net_1\, Y => N_3656);
    
    \REG40M.BIT_OS_VAL_24_RNO[1]\ : MX2B
      port map(A => \BIT_OS_VAL_24[1]\, B => N_206_0, S => 
        \un36_n_bit_os_val[7]\, Y => \N_BIT_OS_VAL_24_18[1]\);
    
    \INDEX_CNT_1_RNIUT8I1[3]\ : MX2
      port map(A => N_4014, B => N_4019, S => 
        \INDEX_CNT_1[3]_net_1\, Y => N_4024);
    
    \REG40M.BIT_OS_VAL_6[3]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_6_18[3]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_2, E => \DES_SM_0[6]_net_1\, Q
         => \BIT_OS_VAL_6[3]\);
    
    \DES_SM_RNIP9OS1[0]\ : NOR3A
      port map(A => I_18, B => \DES_SM_0[8]_net_1\, C => 
        \DES_SM[0]_net_1\, Y => N_5793);
    
    \REG40M.BIT_OS_VAL_3_RNO[2]\ : MX2
      port map(A => N_781, B => \BIT_OS_VAL_3[2]\, S => N_5675, Y
         => N_5652);
    
    \REG40M.BIT_OS_CNT_2[6]\ : DFN1E1C0
      port map(D => BIT_OS_CNT_2_n6, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_5, E => BIT_OS_CNT_2e, Q => 
        \BIT_OS_CNT_2[6]\);
    
    \REG40M.BIT_OS_CNT_1[1]\ : DFN1E1C0
      port map(D => N_139, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_4, E => BIT_OS_CNT_1e, Q => 
        \BIT_OS_CNT_1[1]\);
    
    \CLKPHASE_1_RNI5D5K1[3]\ : MX2
      port map(A => N_3688, B => N_3692, S => 
        \CLKPHASE_1[3]_net_1\, Y => N_3696);
    
    \REG40M.SEQCNTS_5_RNI2O5U[4]\ : MX2
      port map(A => \SEQCNTS_5[4]\, B => \SEQCNTS_6[4]\, S => 
        \INDEX_CNT_2[0]_net_1\, Y => N_4017);
    
    \INDEX_CNT_RNINTCH8[4]\ : MX2
      port map(A => N_4098, B => N_4133, S => 
        \INDEX_CNT[4]_net_1\, Y => N_4138);
    
    \REG40M.BIT_OS_VAL_3_RNO[3]\ : MX2
      port map(A => N_209, B => \BIT_OS_VAL_3[3]\, S => N_5675, Y
         => \N_BIT_OS_VAL_3_18[3]\);
    
    \REG40M.BIT_OS_CNT_4_RNI4OTG1[4]\ : OR3A
      port map(A => N_363, B => N_BIT_OS_VAL_3118lto8_0_o3_2, C
         => N_BIT_OS_VAL_3118lto8_0_o3_1, Y => N_BIT_OS_VAL_3118);
    
    \REG40M.SEQCNTS_27_RNIJ63Q[3]\ : MX2
      port map(A => \SEQCNTS_11[3]\, B => \SEQCNTS_27[3]\, S => 
        \CLKPHASE_2[4]_net_1\, Y => N_3746);
    
    \REG40M.SEQCNTS_24[0]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[0]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_8, E => N_298, Q => \SEQCNTS_24[0]\);
    
    \BEST_BIT_OS_VAL_RNO_19[2]\ : MX2
      port map(A => \BIT_OS_VAL_17[2]\, B => \BIT_OS_VAL_18[2]\, 
        S => \INDEX_CNT_3[0]_net_1\, Y => N_3908);
    
    \WAITCNT[8]\ : DFN1E0C0
      port map(D => N_5718, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_9, E => N_5790, Q => \WAITCNT[8]_net_1\);
    
    \REG40M.BIT_OS_VAL_8_RNI3K6I[1]\ : MX2
      port map(A => \BIT_OS_VAL_8[1]\, B => \BIT_OS_VAL_24[1]\, S
         => \CLKPHASE_1[4]_net_1\, Y => N_3664);
    
    \RECD_SER_WORD_RNO_6[3]\ : OA1
      port map(A => \BIT_OS_SEL[3]_net_1\, B => 
        n_recd_ser_word164, C => \ARB_BYTE[3]_net_1\, Y => 
        \ARB_BYTE_m_2[3]\);
    
    \BEST_BIT_OS_VAL_RNO_28[1]\ : MX2
      port map(A => \BIT_OS_VAL_23[1]\, B => \BIT_OS_VAL_24[1]\, 
        S => \INDEX_CNT_2[0]_net_1\, Y => N_3975);
    
    \REG40M.SEQCNTS_20[1]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[1]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_2, E => N_306, Q => \SEQCNTS_20[1]\);
    
    \REG40M.BIT_OS_VAL_28_RNO[3]\ : MX2
      port map(A => \BIT_OS_VAL_28[3]\, B => N_209_0, S => 
        \un36_n_bit_os_val[3]\, Y => \N_BIT_OS_VAL_28_18[3]\);
    
    \BEST_BIT_OS_VAL_RNO_22[0]\ : MX2
      port map(A => \BIT_OS_VAL_3[0]\, B => \BIT_OS_VAL_4[0]\, S
         => \INDEX_CNT_0[0]_net_1\, Y => N_3934);
    
    \ARB_BYTE_RNI82M33[2]\ : AO1
      port map(A => BIT_OS_CNT_5lde_0_a3_2, B => 
        BIT_OS_CNT_5lde_0_a3_1, C => N_4530_2, Y => BIT_OS_CNT_5e);
    
    \REG40M.SEQCNTS_3_RNIO9VR[0]\ : MX2
      port map(A => \SEQCNTS_3[0]\, B => \SEQCNTS_4[0]\, S => 
        \INDEX_CNT_4[0]_net_1\, Y => N_4068);
    
    \BEST_BIT_OS_VAL_RNO_27[3]\ : MX2
      port map(A => \BIT_OS_VAL_27[3]\, B => \BIT_OS_VAL_28[3]\, 
        S => \INDEX_CNT_1[0]_net_1\, Y => N_3969);
    
    \ADJ_Q[9]\ : DFN1C0
      port map(D => \ADJ_Q[7]_net_1\, CLK => CCC_160M_ADJ, CLR
         => P_MASTER_POR_B_c_34_0, Q => \ADJ_Q[9]_net_1\);
    
    \REG40M.BIT_OS_VAL_8_RNO[0]\ : MX2
      port map(A => \BIT_OS_VAL_8[0]\, B => N_5666_0, S => 
        \un36_n_bit_os_val[23]\, Y => N_276);
    
    \BEST_CLKPHASE_RNO[3]\ : NOR2A
      port map(A => I_9_0, B => \DES_SM_1[8]_net_1\, Y => 
        \N_BEST_CLKPHASE[3]\);
    
    \BEST_BIT_OS_VAL_RNO_11[3]\ : MX2
      port map(A => N_3937, B => N_3941, S => 
        \INDEX_CNT_0[3]_net_1\, Y => N_3945);
    
    \Q[4]\ : DFN1C0
      port map(D => \ADJ_Q[4]_net_1\, CLK => CCC_160M_FXD, CLR
         => P_MASTER_POR_B_c_34, Q => \Q[4]_net_1\);
    
    \REG40M.BIT_OS_VAL_4[1]\ : DFN1E1C0
      port map(D => N_5658, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_20, E => \DES_SM[6]_net_1\, Q => 
        \BIT_OS_VAL_4[1]\);
    
    \REG40M.BIT_OS_CNT_4[6]\ : DFN1E1C0
      port map(D => N_5621, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_9, E => BIT_OS_CNT_4e, Q => 
        \BIT_OS_CNT_4[6]\);
    
    \REG40M.SEQCNTS_17_RNIUEAE[1]\ : MX2
      port map(A => \SEQCNTS_1[1]\, B => \SEQCNTS_17[1]\, S => 
        \CLKPHASE_3[4]_net_1\, Y => N_3759);
    
    \CLKPHASE_RNID3E7_1[3]\ : NOR2A
      port map(A => \CLKPHASE[4]_net_1\, B => \CLKPHASE[3]_net_1\, 
        Y => N_204);
    
    \REG40M.BIT_OS_CNT_7_RNO[4]\ : XA1B
      port map(A => BIT_OS_CNT_7_c3, B => \BIT_OS_CNT_7[4]\, C
         => N_4530_2, Y => BIT_OS_CNT_7_n4);
    
    \CLKPHASE_1_RNIC85U[3]\ : MX2
      port map(A => N_3776, B => N_3781, S => 
        \CLKPHASE_1[3]_net_1\, Y => N_3786);
    
    \BEST_BIT_OS_VAL_RNO_17[0]\ : MX2
      port map(A => \BIT_OS_VAL_5[0]\, B => \BIT_OS_VAL_6[0]\, S
         => \INDEX_CNT_1[0]_net_1\, Y => N_3890);
    
    \REG40M.SEQCNTS_13_RNIVH7C[3]\ : MX2
      port map(A => \SEQCNTS_13[3]\, B => \SEQCNTS_14[3]\, S => 
        \INDEX_CNT_3[0]_net_1\, Y => N_4021);
    
    \REG40M.SEQCNTS_16[4]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[4]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_5, E => N_314, Q => \SEQCNTS_16[4]\);
    
    \REG40M.SEQCNTS_10_RNIEVH31[3]\ : MX2
      port map(A => \SEQCNTS_9[3]\, B => \SEQCNTS_10[3]\, S => 
        \INDEX_CNT_1[0]_net_1\, Y => N_4006);
    
    \BEST_BIT_OS_VAL_RNO_17[2]\ : MX2
      port map(A => \BIT_OS_VAL_5[2]\, B => \BIT_OS_VAL_6[2]\, S
         => \INDEX_CNT_1[0]_net_1\, Y => N_3892);
    
    \REG40M.BIT_OS_CNT_6[0]\ : DFN1E1C0
      port map(D => N_527, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_12, E => BIT_OS_CNT_6e, Q => 
        \BIT_OS_CNT_6[0]\);
    
    \MAX_CNT[0]\ : DFN1E0C0
      port map(D => N_537, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_15, E => N_558, Q => \MAX_CNT[0]_net_1\);
    
    \CLKPHASE_1_RNI525C1[3]\ : MX2
      port map(A => N_3739, B => N_3744, S => 
        \CLKPHASE_1[3]_net_1\, Y => N_3749);
    
    \REG40M.BIT_OS_VAL_11[2]\ : DFN1E1C0
      port map(D => N_197, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_8, E => \DES_SM_1[6]_net_1\, Q => 
        \BIT_OS_VAL_11[2]\);
    
    \REG40M.SEQCNTS_29[2]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[2]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_16_0, E => N_288, Q => \SEQCNTS_29[2]\);
    
    \REG40M.BIT_OS_VAL_4[0]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_4_18[0]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_20, E => \DES_SM[6]_net_1\, Q => 
        \BIT_OS_VAL_4[0]\);
    
    \REG40M.SEQCNTS_27_RNIP2OU[4]\ : MX2
      port map(A => \SEQCNTS_27[4]\, B => \SEQCNTS_28[4]\, S => 
        \INDEX_CNT[0]_net_1\, Y => N_4112);
    
    \REG40M.SEQCNTS_15_RNI0LAD[3]\ : MX2
      port map(A => \SEQCNTS_15[3]\, B => \SEQCNTS_16[3]\, S => 
        \INDEX_CNT_0[0]_net_1\, Y => N_4091);
    
    \REG40M.SEQCNTS_1_RNINQ9K[3]\ : MX2
      port map(A => \SEQCNTS_1[3]\, B => \SEQCNTS_2[3]\, S => 
        \INDEX_CNT_1[0]_net_1\, Y => N_4001);
    
    \BEST_SEQCNT[1]\ : DFN1E1C0
      port map(D => \N_BEST_SEQCNT[1]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_8, E => N_5724, Q => 
        \BEST_SEQCNT[1]_net_1\);
    
    \BEST_BIT_OS_VAL_RNO_10[2]\ : MX2
      port map(A => N_3920, B => \BIT_OS_VAL_29[2]\, S => 
        \INDEX_CNT[3]_net_1\, Y => N_3924);
    
    \MAX_CNT_RNIRTK22[5]\ : OR2A
      port map(A => \MAX_CNT[5]_net_1\, B => N_385, Y => N_388);
    
    \REG40M.SEQCNTS_5_RNIQF5U[0]\ : MX2
      port map(A => \SEQCNTS_5[0]\, B => \SEQCNTS_6[0]\, S => 
        \INDEX_CNT_2[0]_net_1\, Y => N_4013);
    
    \BEST_BIT_OS_VAL_RNO_28[2]\ : MX2
      port map(A => \BIT_OS_VAL_23[2]\, B => \BIT_OS_VAL_24[2]\, 
        S => \INDEX_CNT_2[0]_net_1\, Y => N_3976);
    
    \REG40M.BIT_OS_CNT_0_RNII9K8[4]\ : OR2A
      port map(A => \BIT_OS_CNT_0[4]\, B => N_377, Y => N_383);
    
    \RECD_SER_WORD_RNO_5[7]\ : NOR3C
      port map(A => n_recd_ser_word165_2, B => 
        n_recd_ser_word166_0, C => \ARB_BYTE[9]_net_1\, Y => 
        \ARB_BYTE_m_4[9]\);
    
    \REG40M.BIT_OS_VAL_1_RNI15HO[3]\ : MX2
      port map(A => \BIT_OS_VAL_1[3]\, B => \BIT_OS_VAL_17[3]\, S
         => \CLKPHASE_0[4]_net_1\, Y => N_3630);
    
    \BEST_BIT_OS_VAL_RNO[1]\ : NOR2A
      port map(A => \N_BEST_BIT_OS_VAL_3[1]\, B => 
        \DES_SM[8]_net_1\, Y => \N_BEST_BIT_OS_VAL[1]\);
    
    \REG40M.SEQCNTS_20_RNI1TMJ[2]\ : MX2
      port map(A => \SEQCNTS_19[2]\, B => \SEQCNTS_20[2]\, S => 
        \INDEX_CNT_4[0]_net_1\, Y => N_4105);
    
    \INDEX_CNT_0_RNIEU7A1[3]\ : MX2
      port map(A => N_4119, B => N_4124, S => 
        \INDEX_CNT_0[3]_net_1\, Y => N_4129);
    
    \REG40M.BIT_OS_CNT_6_RNIDCTO[2]\ : OR3C
      port map(A => \BIT_OS_CNT_6[1]\, B => \BIT_OS_CNT_6[2]\, C
         => \BIT_OS_CNT_6[0]\, Y => N_430);
    
    \RECD_SER_WORD_RNO_5[2]\ : NOR3C
      port map(A => n_recd_ser_word165_2, B => 
        n_recd_ser_word166_0, C => \ARB_BYTE[4]_net_1\, Y => 
        \ARB_BYTE_m_1[4]\);
    
    \BEST_BIT_OS_VAL_RNO_5[1]\ : MX2
      port map(A => N_3943, B => N_3955, S => 
        \INDEX_CNT_0[2]_net_1\, Y => N_3959);
    
    \DES_SM_0_RNI4V77I1[8]\ : NOR2A
      port map(A => I_12, B => \DES_SM_0[8]_net_1\, Y => 
        \N_SEQCNTS_1_0[4]\);
    
    \CLKPHASE_1_RNIB4P92[2]\ : MX2
      port map(A => N_3772, B => N_3787, S => 
        \CLKPHASE_1[2]_net_1\, Y => N_3792);
    
    \BEST_BIT_OS_VAL_RNO_14[2]\ : MX2
      port map(A => N_3976, B => N_3980, S => 
        \INDEX_CNT_2[3]_net_1\, Y => N_3984);
    
    \BEST_BIT_OS_VAL_RNO_4[2]\ : MX2
      port map(A => N_3916, B => N_3924, S => 
        \INDEX_CNT_0[2]_net_1\, Y => N_3928);
    
    \CLKPHASE_RNIPVP75[1]\ : MX2
      port map(A => N_3829, B => N_3864, S => \CLKPHASE[1]_net_1\, 
        Y => N_3869);
    
    \BEST_BIT_OS_VAL_RNO_26[1]\ : MX2
      port map(A => \BIT_OS_VAL_19[1]\, B => \BIT_OS_VAL_20[1]\, 
        S => \INDEX_CNT_1[0]_net_1\, Y => N_3963);
    
    \REG40M.BIT_OS_VAL_16_RNO[0]\ : MX2
      port map(A => \BIT_OS_VAL_16[0]\, B => N_5666_0, S => 
        \un36_n_bit_os_val[15]\, Y => N_255);
    
    \REG40M.BIT_OS_VAL_7_RNI2L9J[0]\ : MX2
      port map(A => \BIT_OS_VAL_7[0]\, B => \BIT_OS_VAL_23[0]\, S
         => \CLKPHASE_4[4]_net_1\, Y => N_3603);
    
    \RECD_SER_WORD_RNO[0]\ : OR3
      port map(A => \N_RECD_SER_WORD_iv_1[0]\, B => 
        \N_RECD_SER_WORD_iv_0[0]\, C => \N_RECD_SER_WORD_iv_5[0]\, 
        Y => \N_RECD_SER_WORD[0]\);
    
    \ARB_BYTE_RNIAIJU_0[2]\ : NOR3B
      port map(A => \ARB_BYTE[5]_net_1\, B => N_772, C => 
        \ARB_BYTE[2]_net_1\, Y => BIT_OS_CNT_6lde_0_a3_0);
    
    \REG40M.BIT_OS_VAL_16_RNO[2]\ : MX2
      port map(A => \BIT_OS_VAL_16[2]\, B => N_781_0, S => 
        \un36_n_bit_os_val[15]\, Y => N_189);
    
    \MAX_CNT_RNI3HOD2[6]\ : OR2A
      port map(A => \MAX_CNT[6]_net_1\, B => N_388, Y => N_405);
    
    \MAX_CNT_RNIEQDC1[3]\ : OR2A
      port map(A => \MAX_CNT[3]_net_1\, B => N_370, Y => N_375);
    
    \BEST_BIT_OS_VAL_RNO_0[1]\ : MX2
      port map(A => N_3931, B => N_3991, S => 
        \INDEX_CNT[1]_net_1\, Y => \N_BEST_BIT_OS_VAL_3[1]\);
    
    \Q[10]\ : DFN1C0
      port map(D => \ADJ_Q[10]_net_1\, CLK => CCC_160M_FXD, CLR
         => P_MASTER_POR_B_c_23, Q => \Q[10]_net_1\);
    
    \BEST_BIT_OS_VAL_RNO_4[3]\ : MX2
      port map(A => N_3917, B => N_3925, S => 
        \INDEX_CNT_0[2]_net_1\, Y => N_3929);
    
    \REG40M.BIT_OS_CNT_7_RNO[5]\ : XA1B
      port map(A => BIT_OS_CNT_7_c4, B => \BIT_OS_CNT_7[5]\, C
         => N_4530_2, Y => BIT_OS_CNT_7_n5);
    
    \REG40M.BIT_OS_CNT_2_RNIG7H72[1]\ : OR2
      port map(A => N_BIT_OS_VAL_3110, B => N_BIT_OS_VAL_3114, Y
         => N_445);
    
    \ARB_BYTE_RNI5P9F[1]\ : NOR2A
      port map(A => \ARB_BYTE[4]_net_1\, B => \ARB_BYTE[1]_net_1\, 
        Y => N_776);
    
    \BIT_OS_SEL_1[0]\ : DFN1C0
      port map(D => \BEST_BIT_OS_VAL[0]_net_1\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_27_0, Q => 
        \BIT_OS_SEL_1[0]_net_1\);
    
    \CLKPHASE_RNIP0JI_1[3]\ : OR2A
      port map(A => N_5072_2, B => N_5672, Y => N_5673);
    
    \WAITCNT_RNIEK3P[3]\ : OR2A
      port map(A => \WAITCNT[3]_net_1\, B => N_5773, Y => N_5774);
    
    \REG40M.SEQCNTS_29_RNIV2G41[0]\ : MX2
      port map(A => N_4048, B => \SEQCNTS_29[0]\, S => 
        \INDEX_CNT_2[3]_net_1\, Y => N_4053);
    
    \CLKPHASE_0_RNIN4P33[2]\ : MX2
      port map(A => N_3607, B => N_3619, S => 
        \CLKPHASE_0[2]_net_1\, Y => N_3623);
    
    \REG40M.SEQCNTS_29_RNI59G41[2]\ : MX2
      port map(A => N_4050, B => \SEQCNTS_29[2]\, S => 
        \INDEX_CNT_2[3]_net_1\, Y => N_4055);
    
    \REG40M.BIT_OS_VAL_8_RNI1I6I[0]\ : MX2
      port map(A => \BIT_OS_VAL_8[0]\, B => \BIT_OS_VAL_24[0]\, S
         => \CLKPHASE_1[4]_net_1\, Y => N_3663);
    
    \REG40M.BIT_OS_VAL_2_RNO[2]\ : MX2
      port map(A => N_781, B => \BIT_OS_VAL_2[2]\, S => N_5678, Y
         => N_5653);
    
    \DES_SM_RNO[2]\ : OA1C
      port map(A => \DES_SM_ns_0_i_0_a3_0_1[6]\, B => N_5787, C
         => N_142, Y => N_36);
    
    ADJ_SER_IN_F_0DEL_RNO : MX2
      port map(A => TFC_IN_F, B => ELK0_IN_F, S => DCB_SALT_SEL_c, 
        Y => SER_RX_IN_F);
    
    \DES_SM_0_RNI89UCU2[8]\ : OR3
      port map(A => N_759, B => N_717_0, C => 
        \CLKPHASE_RNIPQFPE1[0]_net_1\, Y => 
        un1_DES_SM_1034_i_o2_2);
    
    \SYNC_SM.N_TUNE_CLKPHASE_2_0_0_ADD_5x5_slow_I1_CO1\ : AO13
      port map(A => I0_un1_CO1, B => \BEST_CLKPHASE[1]_net_1\, C
         => \BEST_SEQCNT[2]_net_1\, Y => N86);
    
    \INDEX_CNT_RNIDMREG[1]\ : MX2
      port map(A => N_4066, B => N_4141, S => 
        \INDEX_CNT[1]_net_1\, Y => \un6_n_best_seqcnt[3]\);
    
    \REG40M.BIT_OS_CNT_4[3]\ : DFN1E1C0
      port map(D => N_45, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_9, E => BIT_OS_CNT_4e, Q => 
        \BIT_OS_CNT_4[3]\);
    
    \REG40M.BIT_OS_CNT_0_RNISOE3[8]\ : OR2
      port map(A => \BIT_OS_CNT_0[4]\, B => \BIT_OS_CNT_0[8]\, Y
         => N_BIT_OS_VAL_312lto8_0_o3_1);
    
    \REG40M.BIT_OS_VAL_15_RNO[2]\ : MX2
      port map(A => \BIT_OS_VAL_15[2]\, B => N_781, S => 
        \un36_n_bit_os_val[16]\, Y => N_191);
    
    \REG40M.BIT_OS_CNT_2[0]\ : DFN1E1C0
      port map(D => N_5610, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_5, E => BIT_OS_CNT_2e, Q => 
        \BIT_OS_CNT_2[0]\);
    
    \INDEX_CNT_RNILFBG2[3]\ : MX2
      port map(A => N_4072, B => N_4077, S => 
        \INDEX_CNT[3]_net_1\, Y => N_4082);
    
    \CLKPHASE_RNIP0JI_0[2]\ : NOR3A
      port map(A => N_211, B => \CLKPHASE[2]_net_1\, C => 
        \CLKPHASE[1]_net_1\, Y => \un36_n_bit_os_val[7]\);
    
    \CLKPHASE_1_RNI845U[3]\ : MX2
      port map(A => N_3775, B => N_3780, S => 
        \CLKPHASE_1[3]_net_1\, Y => N_3785);
    
    \REG40M.BIT_OS_VAL_3_RNI5P911[1]\ : MX2
      port map(A => \BIT_OS_VAL_3[1]\, B => \BIT_OS_VAL_19[1]\, S
         => \CLKPHASE_4[4]_net_1\, Y => N_3612);
    
    \BIT_OS_SEL_2[0]\ : DFN1C0
      port map(D => \BEST_BIT_OS_VAL[0]_net_1\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_27_0, Q => BIT_OS_SEL_2(0));
    
    \REG40M.BIT_OS_VAL_26_RNO[0]\ : MX2
      port map(A => \BIT_OS_VAL_26[0]\, B => N_5666, S => 
        \un36_n_bit_os_val[5]\, Y => N_225);
    
    \CLKPHASE_RNIP0JI[1]\ : OR3A
      port map(A => \CLKPHASE[1]_net_1\, B => N_5663, C => N_5668, 
        Y => N_5675);
    
    \REG40M.SEQCNTS_25[3]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[3]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_10, E => N_296, Q => \SEQCNTS_25[3]\);
    
    \REG40M.BIT_OS_VAL_2_RNO[1]\ : MX2A
      port map(A => N_206, B => \BIT_OS_VAL_2[1]\, S => N_5678, Y
         => N_5660);
    
    \REG40M.SEQCNTS_3[2]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[2]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_11, E => N_340, Q => \SEQCNTS_3[2]\);
    
    \CLKPHASE_2_RNI6IEB1[3]\ : MX2
      port map(A => N_3700, B => N_3704, S => 
        \CLKPHASE_2[3]_net_1\, Y => N_3708);
    
    \CLKPHASE_1_RNI9H5K1[3]\ : MX2
      port map(A => N_3689, B => N_3693, S => 
        \CLKPHASE_1[3]_net_1\, Y => N_3697);
    
    \CLKPHASE_1[3]\ : DFN1C0
      port map(D => \TUNE_CLKPHASE_RNILF0P2[3]_net_1\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_24_0, Q => 
        \CLKPHASE_1[3]_net_1\);
    
    \CLKPHASE_0_RNITQ401[3]\ : MX2
      port map(A => N_3852, B => N_3857, S => 
        \CLKPHASE_0[3]_net_1\, Y => N_3862);
    
    \REG40M.BIT_OS_VAL_26_RNO[2]\ : MX2
      port map(A => \BIT_OS_VAL_26[2]\, B => N_781_0, S => 
        \un36_n_bit_os_val[5]\, Y => N_169);
    
    \REG40M.BIT_OS_VAL_19_RNO[2]\ : MX2
      port map(A => \BIT_OS_VAL_19[2]\, B => N_781, S => 
        \un36_n_bit_os_val[12]\, Y => N_183);
    
    \REG40M.BIT_OS_CNT_4_RNO[2]\ : NOR3A
      port map(A => N_429, B => N_505, C => N_4530_0, Y => N_47);
    
    \REG40M.BIT_OS_VAL_7[0]\ : DFN1E1C0
      port map(D => N_279, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_3, E => \DES_SM_0[6]_net_1\, Q => 
        \BIT_OS_VAL_7[0]\);
    
    \RECD_SER_WORD_RNO_2[2]\ : OR3
      port map(A => \ARB_BYTE_m_1[4]\, B => \ARB_BYTE_m_1[2]\, C
         => \N_RECD_SER_WORD_iv_3[2]\, Y => 
        \N_RECD_SER_WORD_iv_5[2]\);
    
    \CLKPHASE_0_RNI7QOR[3]\ : MX2
      port map(A => N_3726, B => N_3731, S => 
        \CLKPHASE_0[3]_net_1\, Y => N_3736);
    
    \CLKPHASE_0_RNIV0GK5[1]\ : MX2
      port map(A => N_3685, B => N_3713, S => 
        \CLKPHASE_0[1]_net_1\, Y => N_3717);
    
    \REG40M.BIT_OS_VAL_12_RNO[3]\ : MX2
      port map(A => \BIT_OS_VAL_12[3]\, B => N_209, S => 
        \un36_n_bit_os_val[19]\, Y => \N_BIT_OS_VAL_12_18[3]\);
    
    \CLKPHASE_RNIP0JI_8[0]\ : NOR2A
      port map(A => N_214, B => N_5663, Y => 
        \un36_n_bit_os_val[24]\);
    
    un1_CLKPHASE_I_26 : NOR2B
      port map(A => \DWACT_ADD_CI_0_g_array_1[0]\, B => 
        \DWACT_ADD_CI_0_pog_array_1[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_2[0]\);
    
    \REG40M.SEQCNTS_17[4]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[4]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_7, E => N_312, Q => \SEQCNTS_17[4]\);
    
    \MAX_CNT_RNI4OHI[8]\ : NOR2A
      port map(A => \DES_SM[7]_net_1\, B => \MAX_CNT[8]_net_1\, Y
         => DES_SM_tr5_0_a3_1);
    
    \CLKPHASE_0_RNIT8FH4[1]\ : MX2
      port map(A => N_3754, B => N_3789, S => 
        \CLKPHASE_0[1]_net_1\, Y => N_3794);
    
    \BEST_BIT_OS_VAL_RNO_14[0]\ : MX2
      port map(A => N_3974, B => N_3978, S => 
        \INDEX_CNT_2[3]_net_1\, Y => N_3982);
    
    \REG40M.BIT_OS_VAL_10_RNIDMPM[0]\ : MX2
      port map(A => \BIT_OS_VAL_10[0]\, B => \BIT_OS_VAL_26[0]\, 
        S => \CLKPHASE_2[4]_net_1\, Y => N_3691);
    
    \BIT_OS_SEL_2[2]\ : DFN1C0
      port map(D => \BEST_BIT_OS_VAL[2]_net_1\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_27_1, Q => BIT_OS_SEL_2(2));
    
    \REG40M.SEQCNTS_29[4]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[4]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_16_0, E => N_288, Q => \SEQCNTS_29[4]\);
    
    \REG40M.SEQCNTS_28_RNIKDCT[2]\ : MX2
      port map(A => \SEQCNTS_12[2]\, B => \SEQCNTS_28[2]\, S => 
        \CLKPHASE_3[4]_net_1\, Y => N_3820);
    
    \RECD_SER_WORD[6]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[6]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_30, Q => \RECD_SER_WORD[6]_net_1\);
    
    ADJ_SER_IN_F_1DEL : DFN1C0
      port map(D => \ADJ_SER_IN_F_0DEL\, CLK => CCC_160M_ADJ, CLR
         => P_MASTER_POR_B_c_32, Q => \ADJ_SER_IN_F_1DEL\);
    
    \WAITCNT_RNO[5]\ : XA1C
      port map(A => \WAITCNT[5]_net_1\, B => N_5775, C => N_4539, 
        Y => N_34);
    
    \REG40M.BIT_OS_CNT_0_RNI6VS6[3]\ : OR2A
      port map(A => \BIT_OS_CNT_0[3]\, B => N_372, Y => N_377);
    
    \MAX_CNT_RNI9AA11[2]\ : OR3C
      port map(A => \MAX_CNT[0]_net_1\, B => \MAX_CNT[1]_net_1\, 
        C => \MAX_CNT[2]_net_1\, Y => N_370);
    
    \REG40M.SEQCNTS_13_RNITF7C[2]\ : MX2
      port map(A => \SEQCNTS_13[2]\, B => \SEQCNTS_14[2]\, S => 
        \INDEX_CNT_3[0]_net_1\, Y => N_4020);
    
    \CLKPHASE_RNIGVA33[2]\ : MX2
      port map(A => N_3696, B => N_3708, S => \CLKPHASE[2]_net_1\, 
        Y => N_3712);
    
    \REG40M.SEQCNTS_5_RNISH5U[1]\ : MX2
      port map(A => \SEQCNTS_5[1]\, B => \SEQCNTS_6[1]\, S => 
        \INDEX_CNT_2[0]_net_1\, Y => N_4014);
    
    \REG40M.BIT_OS_VAL_21[2]\ : DFN1E1C0
      port map(D => N_179, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_14, E => \DES_SM_2[6]_net_1\, Q => 
        \BIT_OS_VAL_21[2]\);
    
    \BEST_BIT_OS_VAL_RNO_25[2]\ : MX2
      port map(A => \BIT_OS_VAL_15[2]\, B => \BIT_OS_VAL_16[2]\, 
        S => \INDEX_CNT_2[0]_net_1\, Y => N_3952);
    
    \CLKPHASE_RNIINDF1[3]\ : MX2
      port map(A => N_3833, B => N_3838, S => \CLKPHASE[3]_net_1\, 
        Y => N_3843);
    
    \BEST_BIT_OS_VAL_RNO_4[1]\ : MX2
      port map(A => N_3915, B => N_3923, S => 
        \INDEX_CNT_0[2]_net_1\, Y => N_3927);
    
    un3_n_index_cnt_I_11 : NOR2B
      port map(A => \INDEX_CNT[3]_net_1\, B => 
        \DWACT_FINC_E_0[0]\, Y => N_2_0);
    
    \ARB_BYTE_RNI82M33_1[1]\ : AO1
      port map(A => BIT_OS_CNT_6lde_0_a3_1, B => 
        BIT_OS_CNT_6lde_0_a3_0, C => N_4530_1, Y => BIT_OS_CNT_6e);
    
    \REG40M.SEQCNTS_27[2]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[2]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_13, E => N_292, Q => \SEQCNTS_27[2]\);
    
    \REG40M.BIT_OS_VAL_29_RNI82FE[3]\ : MX2
      port map(A => \BIT_OS_VAL_13[3]\, B => \BIT_OS_VAL_29[3]\, 
        S => \CLKPHASE[4]_net_1\, Y => N_3646);
    
    \REG40M.BIT_OS_CNT_0_RNI00B4B[1]\ : NOR2A
      port map(A => N_BIT_OS_VAL_14_18_3_0_a2_1, B => N_781_0, Y
         => N_209_0);
    
    \CLKPHASE_RNIM41A5[1]\ : MX2
      port map(A => N_3832, B => N_3867, S => \CLKPHASE[1]_net_1\, 
        Y => N_3872);
    
    \REG40M.BIT_OS_CNT_4_RNI5I7C[8]\ : OR2
      port map(A => \BIT_OS_CNT_4[8]\, B => \BIT_OS_CNT_4[5]\, Y
         => N_BIT_OS_VAL_3118lto8_0_o3_1);
    
    \CLKPHASE_RNO[0]\ : OA1B
      port map(A => N_5780, B => \TUNE_CLKPHASE[0]_net_1\, C => 
        N_5797, Y => \CLKPHASE_RNO[0]_net_1\);
    
    \REG40M.SEQCNTS_1[3]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[3]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_8, E => N_344, Q => \SEQCNTS_1[3]\);
    
    \REG40M.BIT_OS_CNT_0_RNO_0[8]\ : OR2A
      port map(A => \BIT_OS_CNT_0[7]\, B => N_404, Y => N_435);
    
    \REG40M.BIT_OS_CNT_5[6]\ : DFN1E1C0
      port map(D => N_5626, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_11, E => BIT_OS_CNT_5e, Q => 
        \BIT_OS_CNT_5[6]\);
    
    \REG40M.BIT_OS_VAL_17_RNO[0]\ : MX2
      port map(A => \BIT_OS_VAL_17[0]\, B => N_5666, S => 
        \un36_n_bit_os_val[14]\, Y => N_252);
    
    \CLKPHASE_0_RNIPM401[3]\ : MX2
      port map(A => N_3851, B => N_3856, S => 
        \CLKPHASE_0[3]_net_1\, Y => N_3861);
    
    \BEST_SEQCNT[2]\ : DFN1E1C0
      port map(D => \N_BEST_SEQCNT[2]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_8, E => N_5724, Q => 
        \BEST_SEQCNT[2]_net_1\);
    
    \CLKPHASE_RNIAB7UH7[2]\ : AO1
      port map(A => \un36_n_bit_os_val[23]\, B => N_782_0, C => 
        N_717_0, Y => N_330);
    
    \REG40M.SEQCNTS_30[0]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[0]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_7, E => N_286, Q => \SEQCNTS_30[0]\);
    
    \ARB_WRD_40M_FIXED[13]\ : DFN1C0
      port map(D => \Q[13]_net_1\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_28, Q => \ARB_WRD_40M_FIXED[13]_net_1\);
    
    \REG40M.SEQCNTS_27_RNIF23Q[1]\ : MX2
      port map(A => \SEQCNTS_11[1]\, B => \SEQCNTS_27[1]\, S => 
        \CLKPHASE_2[4]_net_1\, Y => N_3744);
    
    \REG40M.SEQCNTS_13_RNIPKFE[4]\ : MX2
      port map(A => \SEQCNTS_13[4]\, B => \SEQCNTS_29[4]\, S => 
        \CLKPHASE_2[4]_net_1\, Y => N_3782);
    
    \REG40M.BIT_OS_VAL_25_RNO[2]\ : MX2
      port map(A => \BIT_OS_VAL_25[2]\, B => N_781, S => 
        \un36_n_bit_os_val[6]\, Y => N_171);
    
    \MAX_CNT[8]\ : DFN1E0C0
      port map(D => N_89, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_16, E => N_558, Q => \MAX_CNT[8]_net_1\);
    
    \REG40M.BIT_OS_VAL_10[2]\ : DFN1E1C0
      port map(D => N_199, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_6, E => \DES_SM_1[6]_net_1\, Q => 
        \BIT_OS_VAL_10[2]\);
    
    \BEST_BIT_OS_VAL_RNO_12[3]\ : MX2
      port map(A => N_3949, B => N_3953, S => 
        \INDEX_CNT_0[3]_net_1\, Y => N_3957);
    
    \REG40M.SEQCNTS_16[1]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[1]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_5, E => N_314, Q => \SEQCNTS_16[1]\);
    
    \REG40M.BIT_OS_CNT_7[6]\ : DFN1E1C0
      port map(D => BIT_OS_CNT_7_n6, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_14, E => BIT_OS_CNT_7e, Q => 
        \BIT_OS_CNT_7[6]\);
    
    \CLKPHASE_RNIPQFPE1[0]\ : NOR3B
      port map(A => N_762, B => N_1151_tz, C => 
        \un107_bit_os_val[2]\, Y => \CLKPHASE_RNIPQFPE1[0]_net_1\);
    
    \REG40M.SEQCNTS_26_RNIF23Q[1]\ : MX2
      port map(A => \SEQCNTS_10[1]\, B => \SEQCNTS_26[1]\, S => 
        \CLKPHASE_4[4]_net_1\, Y => N_3839);
    
    \MAX_CNT_RNO[3]\ : XA1C
      port map(A => \MAX_CNT[3]_net_1\, B => N_370, C => 
        un1_DES_SM_19, Y => N_5637);
    
    \ARB_BYTE_RNI8GJU[0]\ : NOR3C
      port map(A => \ARB_BYTE[3]_net_1\, B => \ARB_BYTE[0]_net_1\, 
        C => N_776, Y => BIT_OS_CNT_1lde_0_a3_1);
    
    \REG40M.BIT_OS_VAL_29_RNO[2]\ : MX2
      port map(A => \BIT_OS_VAL_29[2]\, B => N_781_0, S => 
        \un36_n_bit_os_val[2]\, Y => N_163);
    
    \REG40M.BIT_OS_CNT_6[6]\ : DFN1E1C0
      port map(D => N_75, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_12, E => BIT_OS_CNT_6e, Q => 
        \BIT_OS_CNT_6[6]\);
    
    \REG40M.BIT_OS_CNT_3[3]\ : DFN1E1C0
      port map(D => BIT_OS_CNT_3_n3, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_7, E => BIT_OS_CNT_3e, Q => 
        \BIT_OS_CNT_3[3]\);
    
    \WAITCNT[11]\ : DFN1E0C0
      port map(D => N_5812, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_21, E => N_5790, Q => 
        \WAITCNT[11]_net_1\);
    
    \BEST_BIT_OS_VAL_RNO_19[0]\ : MX2
      port map(A => \BIT_OS_VAL_17[0]\, B => \BIT_OS_VAL_18[0]\, 
        S => \INDEX_CNT_3[0]_net_1\, Y => N_3906);
    
    \CLKPHASE_RNITRDKE1[0]\ : NOR3A
      port map(A => un1_DES_SM_1034_i_a2_4_2, B => 
        \un107_bit_os_val[0]\, C => \un107_bit_os_val[2]\, Y => 
        N_759);
    
    \REG40M.BIT_OS_VAL_9_RNO[1]\ : MX2B
      port map(A => \BIT_OS_VAL_9[1]\, B => N_206, S => 
        \un36_n_bit_os_val[22]\, Y => \N_BIT_OS_VAL_9_18[1]\);
    
    \REG40M.BIT_OS_VAL_22_RNO[3]\ : MX2
      port map(A => \BIT_OS_VAL_22[3]\, B => N_209_0, S => 
        \un36_n_bit_os_val[9]\, Y => \N_BIT_OS_VAL_22_18[3]\);
    
    \CLKPHASE_1_RNII5VI2[2]\ : MX2
      port map(A => N_3808, B => N_3823, S => 
        \CLKPHASE_1[2]_net_1\, Y => N_3828);
    
    \REG40M.SEQCNTS_5[3]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[3]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_15, E => N_336, Q => \SEQCNTS_5[3]\);
    
    \DES_SM_RNO_1[7]\ : AO1B
      port map(A => DES_SM_tr2_i_a3_6, B => DES_SM_tr2_i_a3_5, C
         => \DES_SM[7]_net_1\, Y => N_54);
    
    \REG40M.BIT_OS_CNT_7[5]\ : DFN1E1C0
      port map(D => BIT_OS_CNT_7_n5, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_14, E => BIT_OS_CNT_7e, Q => 
        \BIT_OS_CNT_7[5]\);
    
    \REG40M.BIT_OS_CNT_6[4]\ : DFN1E1C0
      port map(D => N_79, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_12, E => BIT_OS_CNT_6e, Q => 
        \BIT_OS_CNT_6[4]\);
    
    \DES_SM[6]\ : DFN1C0
      port map(D => N_MAX_CNT_0_sqmuxa, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_27, Q => \DES_SM[6]_net_1\);
    
    \REG40M.SEQCNTS_22[0]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[0]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_5, E => N_302, Q => \SEQCNTS_22[0]\);
    
    \REG40M.BIT_OS_CNT_7_RNI2KJ51[3]\ : NOR2B
      port map(A => BIT_OS_CNT_7_c2, B => \BIT_OS_CNT_7[3]\, Y
         => BIT_OS_CNT_7_c3);
    
    \REG40M.SEQCNTS_8[2]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[2]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_19, E => N_330, Q => \SEQCNTS_8[2]\);
    
    \REG40M.BIT_OS_VAL_31_RNO[2]\ : MX2
      port map(A => \BIT_OS_VAL_31[2]\, B => N_781_0, S => 
        \un36_n_bit_os_val[0]\, Y => N_159);
    
    un1_CLKPHASE_I_18 : XOR2
      port map(A => \CLKPHASE[1]_net_1\, B => 
        \DWACT_ADD_CI_0_TMP[0]\, Y => I_18);
    
    \REG40M.SEQCNTS_8[1]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[1]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_19, E => N_330, Q => \SEQCNTS_8[1]\);
    
    \REG40M.SEQCNTS_12[2]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[2]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_21, E => N_322, Q => \SEQCNTS_12[2]\);
    
    \REG40M.BIT_OS_VAL_17[1]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_17_18[1]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_18, E => \DES_SM_3[6]_net_1\, Q
         => \BIT_OS_VAL_17[1]\);
    
    \REG40M.SEQCNTS_20_RNI1HAG[3]\ : MX2
      port map(A => \SEQCNTS_4[3]\, B => \SEQCNTS_20[3]\, S => 
        \CLKPHASE_5[4]_net_1\, Y => N_3816);
    
    \CLKPHASE_1_RNIDL5K1[3]\ : MX2
      port map(A => N_3690, B => N_3694, S => 
        \CLKPHASE_1[3]_net_1\, Y => N_3698);
    
    \CLKPHASE_0_RNIU0V31[3]\ : MX2
      port map(A => N_3671, B => N_3675, S => 
        \CLKPHASE_0[3]_net_1\, Y => N_3679);
    
    un1_N_CCC_RESET_EN_0_sqmuxa_0_0_a3 : AND2
      port map(A => n_best_clkphase14, B => 
        un1_N_CCC_RESET_EN_0_sqmuxa_0_0_a3_0, Y => N_128);
    
    \REG40M.BIT_OS_VAL_2_RNO[0]\ : MX2
      port map(A => N_5666_0, B => \BIT_OS_VAL_2[0]\, S => N_5678, 
        Y => \N_BIT_OS_VAL_2_18[0]\);
    
    \RECD_SER_WORD_RNO_0[0]\ : AO1
      port map(A => n_recd_ser_word170, B => \ARB_BYTE[6]_net_1\, 
        C => \ARB_BYTE_m[7]\, Y => \N_RECD_SER_WORD_iv_1[0]\);
    
    \DES_SM[8]\ : DFN1P0
      port map(D => \DES_SM_ns[0]\, CLK => CLK_40M_GL, PRE => 
        P_MASTER_POR_B_c_27, Q => \DES_SM[8]_net_1\);
    
    \CLKPHASE_2_RNISS521[3]\ : MX2
      port map(A => N_3798, B => N_3803, S => 
        \CLKPHASE_2[3]_net_1\, Y => N_3808);
    
    \REG40M.SEQCNTS_26_RNIJ63Q[3]\ : MX2
      port map(A => \SEQCNTS_10[3]\, B => \SEQCNTS_26[3]\, S => 
        \CLKPHASE_4[4]_net_1\, Y => N_3841);
    
    \REG40M.BIT_OS_VAL_27_RNO[0]\ : MX2
      port map(A => \BIT_OS_VAL_27[0]\, B => N_5666_0, S => 
        \un36_n_bit_os_val[4]\, Y => N_222);
    
    \REG40M.BIT_OS_VAL_30_RNIHRSP[2]\ : MX2
      port map(A => \BIT_OS_VAL_14[2]\, B => \BIT_OS_VAL_30[2]\, 
        S => \CLKPHASE_3[4]_net_1\, Y => N_3705);
    
    \WAITCNT_RNI5OHC[1]\ : OR2B
      port map(A => \WAITCNT[1]_net_1\, B => \WAITCNT[0]_net_1\, 
        Y => N_5772);
    
    \BEST_CLKPHASE_RNO[0]\ : NOR2
      port map(A => \INDEX_CNT[0]_net_1\, B => 
        \DES_SM_1[8]_net_1\, Y => \N_BEST_CLKPHASE[0]\);
    
    \SYNC_SM.N_TUNE_CLKPHASE_2_0_0_ADD_5x5_slow_I0_un1_CO1\ : 
        OR2A
      port map(A => \BEST_SEQCNT[1]_net_1\, B => 
        \BEST_CLKPHASE[0]_net_1\, Y => I0_un1_CO1);
    
    \REG40M.BIT_OS_CNT_1_RNINO3E[4]\ : OR2A
      port map(A => \BIT_OS_CNT_1[4]\, B => N_380, Y => N_381);
    
    \CLKPHASE_RNI9VD7_0[2]\ : NOR2B
      port map(A => \CLKPHASE[1]_net_1\, B => \CLKPHASE[2]_net_1\, 
        Y => N_5072_2);
    
    \RECD_SER_WORD_RNO_6[4]\ : OA1
      port map(A => \BIT_OS_SEL[3]_net_1\, B => 
        n_recd_ser_word164, C => \ARB_BYTE[4]_net_1\, Y => 
        \ARB_BYTE_m_3[4]\);
    
    \BEST_SEQCNT_RNO[3]\ : NOR2A
      port map(A => \un6_n_best_seqcnt[3]\, B => 
        \DES_SM[8]_net_1\, Y => \N_BEST_SEQCNT[3]\);
    
    \Q[1]\ : DFN1C0
      port map(D => \ADJ_Q[1]_net_1\, CLK => CCC_160M_FXD, CLR
         => P_MASTER_POR_B_c_34, Q => \Q[1]_net_1\);
    
    \INDEX_CNT_RNIIM2N4[2]\ : MX2
      port map(A => N_4079, B => N_4094, S => 
        \INDEX_CNT[2]_net_1\, Y => N_4099);
    
    \DES_SM_1_RNIPHVL2[8]\ : NOR3B
      port map(A => N_5730, B => I_7_0, C => \DES_SM_1[8]_net_1\, 
        Y => \N_INDEX_CNT[2]\);
    
    \BEST_CLKPHASE[3]\ : DFN1E1C0
      port map(D => \N_BEST_CLKPHASE[3]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_10, E => un1_N_CCC_RESET_EN_0_sqmuxa, 
        Q => \BEST_CLKPHASE[3]_net_1\);
    
    \ARB_WRD_40M_FIXED[5]\ : DFN1C0
      port map(D => \Q[5]_net_1\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_26, Q => \ARB_WRD_40M_FIXED[5]_net_1\);
    
    \CLKPHASE_RNIMRDF1[3]\ : MX2
      port map(A => N_3834, B => N_3839, S => \CLKPHASE[3]_net_1\, 
        Y => N_3844);
    
    \BEST_BIT_OS_VAL_RNO_1[1]\ : MX2
      port map(A => N_3903, B => N_3927, S => 
        \INDEX_CNT[4]_net_1\, Y => N_3931);
    
    \REG40M.SEQCNTS_21[2]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[2]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_3, E => N_304, Q => \SEQCNTS_21[2]\);
    
    \INDEX_CNT_RNIHRHU3[2]\ : MX2
      port map(A => N_4012, B => N_4027, S => 
        \INDEX_CNT[2]_net_1\, Y => N_4032);
    
    \BIT_OS_SEL_RNIQPQF[3]\ : NOR2
      port map(A => \BIT_OS_SEL[3]_net_1\, B => 
        \BIT_OS_SEL[1]_net_1\, Y => n_recd_ser_word168_2);
    
    \REG40M.BIT_OS_CNT_2[7]\ : DFN1E1C0
      port map(D => BIT_OS_CNT_2_n7, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_5, E => BIT_OS_CNT_2e, Q => 
        \BIT_OS_CNT_2[7]\);
    
    \REG40M.SEQCNTS_15_RNICQS9[1]\ : MX2
      port map(A => \SEQCNTS_31[1]\, B => \SEQCNTS_15[1]\, S => 
        \CLKPHASE_0[4]_net_1\, Y => N_3724);
    
    \REG40M.BIT_OS_VAL_3_RNI8UC21[2]\ : MX2
      port map(A => \BIT_OS_VAL_3[2]\, B => \BIT_OS_VAL_19[2]\, S
         => \CLKPHASE_5[4]_net_1\, Y => N_3613);
    
    \DES_SM_RNI74OM_1[7]\ : NOR3B
      port map(A => \ARB_BYTE[7]_net_1\, B => \DES_SM[7]_net_1\, 
        C => \ARB_BYTE[6]_net_1\, Y => N_559_1);
    
    \REG40M.BIT_OS_VAL_14[0]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_14_18[0]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_13, E => \DES_SM_2[6]_net_1\, Q
         => \BIT_OS_VAL_14[0]\);
    
    \REG40M.BIT_OS_VAL_6_RNO[1]\ : MX2A
      port map(A => N_206_0, B => \BIT_OS_VAL_6[1]\, S => N_5677, 
        Y => N_5657);
    
    \DES_SM_RNI652GA[0]\ : AO1
      port map(A => un1_DES_SM_471_i_0_0_a3_0_0, B => N_5859, C
         => un1_DES_SM_471_i_0_0_0_1, Y => N_4539);
    
    \CLKPHASE_1_RNI405U[3]\ : MX2
      port map(A => N_3774, B => N_3779, S => 
        \CLKPHASE_1[3]_net_1\, Y => N_3784);
    
    \BEST_BIT_OS_VAL_RNO_20[1]\ : MX2
      port map(A => \BIT_OS_VAL_25[1]\, B => \BIT_OS_VAL_26[1]\, 
        S => \INDEX_CNT_3[0]_net_1\, Y => N_3911);
    
    \WAITCNT_RNO[2]\ : XA1C
      port map(A => \WAITCNT[2]_net_1\, B => N_5772, C => N_4539, 
        Y => N_41);
    
    \REG40M.SEQCNTS_13_RNIHCFE[0]\ : MX2
      port map(A => \SEQCNTS_13[0]\, B => \SEQCNTS_29[0]\, S => 
        \CLKPHASE_2[4]_net_1\, Y => N_3778);
    
    \REG40M.SEQCNTS_24_RNIA80O[4]\ : MX2
      port map(A => \SEQCNTS_8[4]\, B => \SEQCNTS_24[4]\, S => 
        \CLKPHASE_4[4]_net_1\, Y => N_3807);
    
    \REG40M.BIT_OS_CNT_4_RNIG8KA3[4]\ : OR2
      port map(A => N_BIT_OS_VAL_3118, B => N_BIT_OS_VAL_3122, Y
         => N_437);
    
    \CLKPHASE_RNIU3EF1[3]\ : MX2
      port map(A => N_3836, B => N_3841, S => \CLKPHASE[3]_net_1\, 
        Y => N_3846);
    
    \CLKPHASE_0_RNISN8K5[1]\ : MX2
      port map(A => N_3623, B => N_3651, S => 
        \CLKPHASE_0[1]_net_1\, Y => N_3655);
    
    \BEST_CLKPHASE[2]\ : DFN1E1C0
      port map(D => \N_BEST_CLKPHASE[2]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_10, E => un1_N_CCC_RESET_EN_0_sqmuxa, 
        Q => \BEST_CLKPHASE[2]_net_1\);
    
    \REG40M.BIT_OS_VAL_0_RNO[2]\ : MX2
      port map(A => N_781, B => \BIT_OS_VAL_0[2]\, S => N_5679, Y
         => N_5655);
    
    un3_n_index_cnt_I_5 : XOR2
      port map(A => \INDEX_CNT[0]_net_1\, B => 
        \INDEX_CNT[1]_net_1\, Y => I_5_0);
    
    \REG40M.SEQCNTS_4[4]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[4]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_13, E => N_338, Q => \SEQCNTS_4[4]\);
    
    \REG40M.BIT_OS_VAL_11[1]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_11_18[1]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_8, E => \DES_SM_1[6]_net_1\, Q
         => \BIT_OS_VAL_11[1]\);
    
    \CLKPHASE_RNI80B0A[0]\ : MX2
      port map(A => N_3796, B => N_3871, S => \CLKPHASE[0]_net_1\, 
        Y => \un39_n_seqcnts[3]\);
    
    un1_N_CCC_RESET_EN_0_sqmuxa_0_0 : OR2
      port map(A => N_5784_i, B => N_128, Y => 
        un1_N_CCC_RESET_EN_0_sqmuxa);
    
    \REG40M.SEQCNTS_16[0]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[0]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_5, E => N_314, Q => \SEQCNTS_16[0]\);
    
    \REG40M.SEQCNTS_11_RNIS8U81[3]\ : MX2
      port map(A => \SEQCNTS_11[3]\, B => \SEQCNTS_12[3]\, S => 
        \INDEX_CNT_4[0]_net_1\, Y => N_4076);
    
    \RECD_SER_WORD_RNI82R61[1]\ : NOR3B
      port map(A => \RECD_SER_WORD[1]_net_1\, B => 
        \RECD_SER_WORD[2]_net_1\, C => \ELK_RX_SER_WORD_0[4]\, Y
         => ELK0_SYNC_DET_1_1);
    
    \REG40M.SEQCNTS_23[3]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[3]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_6, E => N_300, Q => \SEQCNTS_23[3]\);
    
    \INDEX_CNT_1[3]\ : DFN1E0C0
      port map(D => \N_INDEX_CNT[3]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_17_0, E => N_5149, Q => 
        \INDEX_CNT_1[3]_net_1\);
    
    \ADJ_Q[0]\ : DFN1C0
      port map(D => \ADJ_SER_IN_R_1DEL\, CLK => CCC_160M_ADJ, CLR
         => P_MASTER_POR_B_c_34_0, Q => \ADJ_Q[0]_net_1\);
    
    \BEST_BIT_OS_VAL_RNO_2[2]\ : MX2
      port map(A => N_3960, B => N_3988, S => 
        \INDEX_CNT[4]_net_1\, Y => N_3992);
    
    \REG40M.SEQCNTS_1[1]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[1]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_8, E => N_344, Q => \SEQCNTS_1[1]\);
    
    \REG40M.BIT_OS_CNT_6_RNIK8F22[7]\ : OR3A
      port map(A => N_365, B => N_BIT_OS_VAL_3126lto8_0_o3_0, C
         => N_354, Y => N_BIT_OS_VAL_3126);
    
    \REG40M.BIT_OS_CNT_1[5]\ : DFN1E1C0
      port map(D => N_131, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_4, E => BIT_OS_CNT_1e, Q => 
        \BIT_OS_CNT_1[5]\);
    
    \BEST_BIT_OS_VAL_RNO_8[1]\ : MX2
      port map(A => N_3891, B => N_3895, S => 
        \INDEX_CNT_1[3]_net_1\, Y => N_3899);
    
    \BEST_BIT_OS_VAL[3]\ : DFN1E1C0
      port map(D => \N_BEST_BIT_OS_VAL[3]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_14, E => 
        un1_N_CCC_RESET_EN_0_sqmuxa, Q => 
        \BEST_BIT_OS_VAL[3]_net_1\);
    
    \BEST_BIT_OS_VAL_RNO_7[3]\ : MX2
      port map(A => N_3881, B => N_3885, S => 
        \INDEX_CNT_0[3]_net_1\, Y => N_3889);
    
    \RECD_SER_WORD_RNO_0[5]\ : AO1
      port map(A => \ARB_BYTE[11]_net_1\, B => n_recd_ser_word170, 
        C => \ARB_BYTE_m[12]\, Y => \N_RECD_SER_WORD_iv_1[5]\);
    
    \INDEX_CNT_RNITNR6G[1]\ : MX2
      port map(A => N_4064, B => N_4139, S => 
        \INDEX_CNT[1]_net_1\, Y => \un6_n_best_seqcnt[1]\);
    
    \BIT_OS_SEL_5[0]\ : DFN1C0
      port map(D => \BEST_BIT_OS_VAL[0]_net_1\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_27_0, Q => BIT_OS_SEL_5(0));
    
    \INDEX_CNT_4[0]\ : DFN1E0C0
      port map(D => \N_INDEX_CNT[0]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_16_0, E => N_5149, Q => 
        \INDEX_CNT_4[0]_net_1\);
    
    \DES_SM_RNITN4L[2]\ : AO16
      port map(A => \WAITCNT[0]_net_1\, B => \DES_SM[2]_net_1\, C
         => \DES_SM[3]_net_1\, Y => N_123);
    
    \REG40M.BIT_OS_VAL_18[1]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_18_18[1]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_19, E => \DES_SM_4[6]_net_1\, Q
         => \BIT_OS_VAL_18[1]\);
    
    \REG40M.SEQCNTS_7[1]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[1]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_17_0, E => N_332, Q => \SEQCNTS_7[1]\);
    
    \CLKPHASE_RNIP0JI_5[0]\ : NOR2B
      port map(A => N_214, B => N_215, Y => 
        \un36_n_bit_os_val[0]\);
    
    \CLKPHASE_1_RNIH5I72[2]\ : MX2
      port map(A => N_3769, B => N_3784, S => 
        \CLKPHASE_1[2]_net_1\, Y => N_3789);
    
    \SYNC_SM.N_TUNE_CLKPHASE_2_0_0_ADD_5x5_slow_I3_CO1\ : AO13
      port map(A => I2_un1_CO1, B => \BEST_CLKPHASE[3]_net_1\, C
         => \BEST_SEQCNT[4]_net_1\, Y => N90);
    
    \DES_SM_RNI1EH11[0]\ : MX2B
      port map(A => \DES_SM[0]_net_1\, B => CCC_RX_CLK_LOCK, S
         => N_5783, Y => un1_DES_SM_471_i_0_0_a3_0_0);
    
    \BIT_OS_SEL_1_RNII4DE1_0[0]\ : NOR3B
      port map(A => \BIT_OS_SEL_1[2]_net_1\, B => 
        n_recd_ser_word168_2, C => \BIT_OS_SEL_1[0]_net_1\, Y => 
        n_recd_ser_word168);
    
    \ADJ_Q[4]\ : DFN1C0
      port map(D => \ADJ_Q[2]_net_1\, CLK => CCC_160M_ADJ, CLR
         => P_MASTER_POR_B_c_34_0, Q => \ADJ_Q[4]_net_1\);
    
    \REG40M.SEQCNTS_18_RNI3QJH[2]\ : MX2
      port map(A => \SEQCNTS_2[2]\, B => \SEQCNTS_18[2]\, S => 
        \CLKPHASE_4[4]_net_1\, Y => N_3835);
    
    \REG40M.BIT_OS_CNT_0_RNO[3]\ : XA1C
      port map(A => \BIT_OS_CNT_0[3]\, B => N_372, C => N_4530_2, 
        Y => N_117);
    
    \REG40M.SEQCNTS_26_RNID03Q[0]\ : MX2
      port map(A => \SEQCNTS_10[0]\, B => \SEQCNTS_26[0]\, S => 
        \CLKPHASE_4[4]_net_1\, Y => N_3838);
    
    \REG40M.SEQCNTS_19_RNIUIGG[0]\ : MX2
      port map(A => \SEQCNTS_3[0]\, B => \SEQCNTS_19[0]\, S => 
        \CLKPHASE_1[4]_net_1\, Y => N_3738);
    
    \DES_SM_RNIDEA0K[8]\ : NOR2A
      port map(A => I_5, B => \DES_SM[8]_net_1\, Y => 
        \N_SEQCNTS_1[1]\);
    
    \CLKPHASE_2_RNIK1FE1[3]\ : MX2
      port map(A => N_3627, B => N_3631, S => 
        \CLKPHASE_2[3]_net_1\, Y => N_3635);
    
    \BEST_BIT_OS_VAL_RNO_25[1]\ : MX2
      port map(A => \BIT_OS_VAL_15[1]\, B => \BIT_OS_VAL_16[1]\, 
        S => \INDEX_CNT_2[0]_net_1\, Y => N_3951);
    
    \DES_SM[4]\ : DFN1C0
      port map(D => \DES_SM_RNO[4]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_27, Q => \DES_SM[4]_net_1\);
    
    \CLKPHASE_1_RNIBEK8H7_0[2]\ : AO1
      port map(A => \un36_n_bit_os_val[5]\, B => N_782, C => 
        N_717, Y => N_294);
    
    \RECD_SER_WORD_RNILBNR[0]\ : NOR3A
      port map(A => \RECD_SER_WORD[3]_net_1\, B => 
        \RECD_SER_WORD[4]_net_1\, C => \RECD_SER_WORD[0]_net_1\, 
        Y => TFC_SYNC_DET_1_2);
    
    \RECD_SER_WORD_RNO[5]\ : OR3
      port map(A => \N_RECD_SER_WORD_iv_1[5]\, B => 
        \N_RECD_SER_WORD_iv_0[5]\, C => \N_RECD_SER_WORD_iv_5[5]\, 
        Y => \N_RECD_SER_WORD[5]\);
    
    \REG40M.BIT_OS_VAL_20[2]\ : DFN1E1C0
      port map(D => N_181, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_13, E => \DES_SM_2[6]_net_1\, Q => 
        \BIT_OS_VAL_20[2]\);
    
    \RECD_SER_WORD_RNIJJBK[6]\ : NOR2B
      port map(A => \RECD_SER_WORD[6]_net_1\, B => DCB_SALT_SEL_c, 
        Y => \ELK_RX_SER_WORD_0[6]\);
    
    \RECD_SER_WORD_RNO_7[3]\ : AO1
      port map(A => n_recd_ser_word165, B => \ARB_BYTE[4]_net_1\, 
        C => \ARB_BYTE_m_2[6]\, Y => \N_RECD_SER_WORD_iv_3[3]\);
    
    \BEST_BIT_OS_VAL_RNO_11[1]\ : MX2
      port map(A => N_3935, B => N_3939, S => 
        \INDEX_CNT_0[3]_net_1\, Y => N_3943);
    
    \REG40M.SEQCNTS_27_RNIHQNU[0]\ : MX2
      port map(A => \SEQCNTS_27[0]\, B => \SEQCNTS_28[0]\, S => 
        \INDEX_CNT[0]_net_1\, Y => N_4108);
    
    \REG40M.BIT_OS_VAL_2_RNI2CQR[2]\ : MX2
      port map(A => \BIT_OS_VAL_2[2]\, B => \BIT_OS_VAL_18[2]\, S
         => \CLKPHASE_1[4]_net_1\, Y => N_3689);
    
    \CLKPHASE_RNIP0JI_2[2]\ : NOR3
      port map(A => \CLKPHASE[2]_net_1\, B => \CLKPHASE[1]_net_1\, 
        C => N_5672, Y => \un36_n_bit_os_val[23]\);
    
    \REG40M.SEQCNTS_21[4]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[4]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_3, E => N_304, Q => \SEQCNTS_21[4]\);
    
    \CLKPHASE_1_RNI6E2A1[3]\ : MX2
      port map(A => N_3762, B => N_3767, S => 
        \CLKPHASE_1[3]_net_1\, Y => N_3772);
    
    \REG40M.SEQCNTS_30[1]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[1]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_7, E => N_286, Q => \SEQCNTS_30[1]\);
    
    \REG40M.SEQCNTS_20_RNITCAG[1]\ : MX2
      port map(A => \SEQCNTS_4[1]\, B => \SEQCNTS_20[1]\, S => 
        \CLKPHASE_5[4]_net_1\, Y => N_3814);
    
    \REG40M.SEQCNTS_18_RNI1OJH[1]\ : MX2
      port map(A => \SEQCNTS_2[1]\, B => \SEQCNTS_18[1]\, S => 
        \CLKPHASE_4[4]_net_1\, Y => N_3834);
    
    \INDEX_CNT_1_RNILK2O1[3]\ : MX2
      port map(A => N_4036, B => N_4041, S => 
        \INDEX_CNT_1[3]_net_1\, Y => N_4046);
    
    \DES_SM_0_RNIII0V[8]\ : OR2
      port map(A => \DES_SM_0[8]_net_1\, B => \DES_SM_0[6]_net_1\, 
        Y => N_4530_2);
    
    \BEST_BIT_OS_VAL_RNO_10[3]\ : MX2
      port map(A => N_3921, B => \BIT_OS_VAL_29[3]\, S => 
        \INDEX_CNT[3]_net_1\, Y => N_3925);
    
    \INDEX_CNT_1_RNIFI3J1[3]\ : OR3B
      port map(A => \INDEX_CNT_1[3]_net_1\, B => 
        \INDEX_CNT_2[0]_net_1\, C => DES_SM_tr8_i_o2_1, Y => 
        N_5730);
    
    \DES_SM_RNI5E9L1[0]\ : NOR3A
      port map(A => I_21, B => \DES_SM_1[8]_net_1\, C => 
        \DES_SM[0]_net_1\, Y => N_5795);
    
    \CLKPHASE_RNICU2EH7[1]\ : AO1
      port map(A => \un36_n_bit_os_val[14]\, B => N_782, C => 
        N_717, Y => N_312);
    
    \CLKPHASE[3]\ : DFN1C0
      port map(D => \TUNE_CLKPHASE_RNILF0P2[3]_net_1\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_24_0, Q => 
        \CLKPHASE[3]_net_1\);
    
    \ARB_BYTE_RNIEV161[2]\ : NOR3B
      port map(A => \ARB_BYTE[2]_net_1\, B => N_559_1, C => 
        \ARB_BYTE[5]_net_1\, Y => BIT_OS_CNT_0lde_0_a3_1);
    
    \DES_SM_1[8]\ : DFN1P0
      port map(D => \DES_SM_ns[0]\, CLK => CLK_40M_GL, PRE => 
        P_MASTER_POR_B_c_27_1, Q => \DES_SM_1[8]_net_1\);
    
    \REG40M.BIT_OS_VAL_27[1]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_27_18[1]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_2, E => \DES_SM_0[6]_net_1\, Q
         => \BIT_OS_VAL_27[1]\);
    
    \WAITCNT_RNI1T1L3[1]\ : NOR3C
      port map(A => un1_DES_SM_471_i_0_a2_0_0_a2_8, B => 
        un1_DES_SM_471_i_0_a2_0_0_a2_7, C => 
        un1_DES_SM_471_i_0_a2_0_0_a2_9, Y => N_116);
    
    \REG40M.SEQCNTS_31_RNIFN4I[2]\ : NOR2A
      port map(A => \SEQCNTS_31[2]\, B => \INDEX_CNT[0]_net_1\, Y
         => N_4125);
    
    \REG40M.BIT_OS_CNT_5_RNICGMP1[1]\ : OR3
      port map(A => N_760, B => N_BIT_OS_VAL_3122lto8_0_o3_1, C
         => N_BIT_OS_VAL_3122lto8_0_o3_2, Y => N_BIT_OS_VAL_3122);
    
    \CLKPHASE_RNIB5DBB[0]\ : MX2
      port map(A => N_3657, B => N_3717, S => \CLKPHASE[0]_net_1\, 
        Y => \un107_bit_os_val[2]\);
    
    \REG40M.SEQCNTS_20[2]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[2]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_2, E => N_306, Q => \SEQCNTS_20[2]\);
    
    \REG40M.BIT_OS_VAL_9_RNI8R9J[3]\ : MX2
      port map(A => \BIT_OS_VAL_9[3]\, B => \BIT_OS_VAL_25[3]\, S
         => \CLKPHASE_0[4]_net_1\, Y => N_3634);
    
    \CLKPHASE_0_RNIJ91G2[2]\ : MX2
      port map(A => N_3847, B => N_3862, S => 
        \CLKPHASE_0[2]_net_1\, Y => N_3867);
    
    \INDEX_CNT_2_RNIR9AR1[3]\ : MX2
      port map(A => N_4086, B => N_4091, S => 
        \INDEX_CNT_2[3]_net_1\, Y => N_4096);
    
    \BEST_BIT_OS_VAL_RNO_15[0]\ : MX2
      port map(A => \BIT_OS_VAL_1[0]\, B => \BIT_OS_VAL_2[0]\, S
         => \INDEX_CNT_0[0]_net_1\, Y => N_3878);
    
    \REG40M.BIT_OS_CNT_1_RNO[2]\ : NOR3A
      port map(A => N_428, B => N_555, C => N_4530_0, Y => N_137);
    
    \REG40M.SEQCNTS_8[0]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[0]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_19, E => N_330, Q => \SEQCNTS_8[0]\);
    
    \REG40M.BIT_OS_CNT_7[1]\ : DFN1E1C0
      port map(D => BIT_OS_CNT_7_n1, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_14, E => BIT_OS_CNT_7e, Q => 
        \BIT_OS_CNT_7[1]\);
    
    \REG40M.SEQCNTS_3_RNIQBVR[1]\ : MX2
      port map(A => \SEQCNTS_3[1]\, B => \SEQCNTS_4[1]\, S => 
        \INDEX_CNT_4[0]_net_1\, Y => N_4069);
    
    \RECD_SER_WORD_RNIGGBK_0[3]\ : NOR2A
      port map(A => \RECD_SER_WORD[3]_net_1\, B => DCB_SALT_SEL_c, 
        Y => TFC_RX_SER_WORD(3));
    
    \REG40M.SEQCNTS_17_RNI360L[1]\ : MX2
      port map(A => \SEQCNTS_17[1]\, B => \SEQCNTS_18[1]\, S => 
        \INDEX_CNT_3[0]_net_1\, Y => N_4034);
    
    \REG40M.SEQCNTS_25[1]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[1]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_10, E => N_296, Q => \SEQCNTS_25[1]\);
    
    \REG40M.BIT_OS_CNT_7[0]\ : DFN1E1C0
      port map(D => N_5615, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_14, E => BIT_OS_CNT_7e, Q => 
        \BIT_OS_CNT_7[0]\);
    
    \REG40M.BIT_OS_VAL_5_RNO[3]\ : MX2
      port map(A => \BIT_OS_VAL_5[3]\, B => N_209_0, S => 
        \un36_n_bit_os_val[26]\, Y => \N_BIT_OS_VAL_5_18[3]\);
    
    \REG40M.SEQCNTS_25[2]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[2]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_10, E => N_296, Q => \SEQCNTS_25[2]\);
    
    \INDEX_CNT_0[3]\ : DFN1E0C0
      port map(D => \N_INDEX_CNT[3]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_17_0, E => N_5149, Q => 
        \INDEX_CNT_0[3]_net_1\);
    
    \REG40M.SEQCNTS_16_RNI3FH7[0]\ : NOR2B
      port map(A => \SEQCNTS_16[0]\, B => \CLKPHASE[4]_net_1\, Y
         => N_3798);
    
    \CLKPHASE_1_RNI9TH72[2]\ : MX2
      port map(A => N_3768, B => N_3783, S => 
        \CLKPHASE_1[2]_net_1\, Y => N_3788);
    
    \BEST_SEQCNT[4]\ : DFN1E1C0
      port map(D => \N_BEST_SEQCNT[4]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_9, E => N_5724, Q => 
        \BEST_SEQCNT[4]_net_1\);
    
    \RECD_SER_WORD[1]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[1]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_29, Q => \RECD_SER_WORD[1]_net_1\);
    
    \BIT_OS_SEL_RNIONQF[0]\ : NOR2B
      port map(A => \BIT_OS_SEL[0]_net_1\, B => 
        \BIT_OS_SEL[2]_net_1\, Y => n_recd_ser_word169_0);
    
    \REG40M.BIT_OS_VAL_24[0]\ : DFN1E1C0
      port map(D => N_231, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_18, E => \DES_SM_4[6]_net_1\, Q => 
        \BIT_OS_VAL_24[0]\);
    
    \WAITCNT_RNI12QU1[9]\ : OR2A
      port map(A => \WAITCNT[9]_net_1\, B => N_5779, Y => N_5781);
    
    \CLKPHASE_2[3]\ : DFN1C0
      port map(D => \TUNE_CLKPHASE_RNILF0P2[3]_net_1\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_24_0, Q => 
        \CLKPHASE_2[3]_net_1\);
    
    \CLKPHASE_2_RNIG81I1[3]\ : MX2
      port map(A => N_3601, B => N_3605, S => 
        \CLKPHASE_2[3]_net_1\, Y => N_3609);
    
    \CLKPHASE_0_RNIADV31[3]\ : MX2
      port map(A => N_3674, B => N_3678, S => 
        \CLKPHASE_0[3]_net_1\, Y => N_3682);
    
    \REG40M.BIT_OS_VAL_3[2]\ : DFN1E1C0
      port map(D => N_5652, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_19, E => \DES_SM_4[6]_net_1\, Q => 
        \BIT_OS_VAL_3[2]\);
    
    \REG40M.BIT_OS_CNT_5_RNIBL141[4]\ : OR2A
      port map(A => \BIT_OS_CNT_5[4]\, B => N_376, Y => N_384);
    
    \DES_SM_RNO_2[7]\ : MX2
      port map(A => \DES_SM[3]_net_1\, B => \DES_SM[2]_net_1\, S
         => \WAITCNT[0]_net_1\, Y => N_70);
    
    \REG40M.BIT_OS_VAL_27_RNII59C[0]\ : MX2
      port map(A => \BIT_OS_VAL_11[0]\, B => \BIT_OS_VAL_27[0]\, 
        S => \CLKPHASE_5[4]_net_1\, Y => N_3615);
    
    \REG40M.BIT_OS_VAL_13_RNO[1]\ : MX2B
      port map(A => \BIT_OS_VAL_13[1]\, B => N_206, S => 
        \un36_n_bit_os_val[18]\, Y => \N_BIT_OS_VAL_13_18[1]\);
    
    \REG40M.BIT_OS_VAL_21[1]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_21_18[1]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_14, E => \DES_SM_2[6]_net_1\, Q
         => \BIT_OS_VAL_21[1]\);
    
    \CLKPHASE_1_RNI965C1[3]\ : MX2
      port map(A => N_3740, B => N_3745, S => 
        \CLKPHASE_1[3]_net_1\, Y => N_3750);
    
    \REG40M.SEQCNTS_5[4]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[4]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_15, E => N_336, Q => \SEQCNTS_5[4]\);
    
    \INDEX_CNT_RNI4CEH8[4]\ : MX2
      port map(A => N_4101, B => N_4136, S => 
        \INDEX_CNT[4]_net_1\, Y => N_4141);
    
    \CLKPHASE_1_RNI1N2K2[2]\ : MX2
      port map(A => N_3810, B => N_3825, S => 
        \CLKPHASE_1[2]_net_1\, Y => N_3830);
    
    \REG40M.BIT_OS_VAL_28_RNIJ009[2]\ : MX2
      port map(A => \BIT_OS_VAL_12[2]\, B => \BIT_OS_VAL_28[2]\, 
        S => \CLKPHASE_0[4]_net_1\, Y => N_3677);
    
    \BEST_BIT_OS_VAL_RNO_6[1]\ : MX2
      port map(A => N_3971, B => N_3983, S => 
        \INDEX_CNT[2]_net_1\, Y => N_3987);
    
    \INDEX_CNT_RNI93BG2[3]\ : MX2
      port map(A => N_4069, B => N_4074, S => 
        \INDEX_CNT[3]_net_1\, Y => N_4079);
    
    \BEST_BIT_OS_VAL_RNO_12[2]\ : MX2
      port map(A => N_3948, B => N_3952, S => 
        \INDEX_CNT_0[3]_net_1\, Y => N_3956);
    
    \REG40M.BIT_OS_CNT_3_RNO[1]\ : XA1B
      port map(A => \BIT_OS_CNT_3[1]\, B => \BIT_OS_CNT_3[0]\, C
         => N_4530_1, Y => BIT_OS_CNT_3_n1);
    
    \BEST_BIT_OS_VAL_RNO_8[2]\ : MX2
      port map(A => N_3892, B => N_3896, S => 
        \INDEX_CNT_1[3]_net_1\, Y => N_3900);
    
    \REG40M.BIT_OS_VAL_10_RNIFOPM[1]\ : MX2
      port map(A => \BIT_OS_VAL_10[1]\, B => \BIT_OS_VAL_26[1]\, 
        S => \CLKPHASE_2[4]_net_1\, Y => N_3692);
    
    \RECD_SER_WORD_RNO_7[0]\ : AO1
      port map(A => \ARB_BYTE[1]_net_1\, B => n_recd_ser_word165, 
        C => \ARB_BYTE_m[3]\, Y => \N_RECD_SER_WORD_iv_3[0]\);
    
    \BEST_BIT_OS_VAL_RNO_0[2]\ : MX2
      port map(A => N_3932, B => N_3992, S => 
        \INDEX_CNT[1]_net_1\, Y => \N_BEST_BIT_OS_VAL_3[2]\);
    
    \REG40M.BIT_OS_CNT_0_RNO[6]\ : XA1C
      port map(A => \BIT_OS_CNT_0[6]\, B => N_390, C => N_4530_2, 
        Y => N_111);
    
    \ARB_BYTE_RNIEV161_1[2]\ : NOR3B
      port map(A => \ARB_BYTE[2]_net_1\, B => N_560_2, C => 
        \ARB_BYTE[5]_net_1\, Y => BIT_OS_CNT_1lde_0_a3_2);
    
    \REG40M.BIT_OS_VAL_28[1]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_28_18[1]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_2, E => \DES_SM_0[6]_net_1\, Q
         => \BIT_OS_VAL_28[1]\);
    
    \RECD_SER_WORD_RNO[7]\ : OR3
      port map(A => \N_RECD_SER_WORD_iv_1[7]\, B => 
        \N_RECD_SER_WORD_iv_0[7]\, C => \N_RECD_SER_WORD_iv_5[7]\, 
        Y => \N_RECD_SER_WORD[7]\);
    
    \REG40M.SEQCNTS_21_RNIP97G[1]\ : MX2
      port map(A => \SEQCNTS_21[1]\, B => \SEQCNTS_22[1]\, S => 
        \INDEX_CNT_3[0]_net_1\, Y => N_4049);
    
    \CLKPHASE_RNI83F1A[0]\ : MX2
      port map(A => N_3797, B => N_3872, S => \CLKPHASE[0]_net_1\, 
        Y => \un39_n_seqcnts[4]\);
    
    \SYNC_SM.N_TUNE_CLKPHASE_2_0_0_ADD_5x5_slow_I2_un1_CO1\ : 
        AO13
      port map(A => N86, B => \BEST_CLKPHASE[2]_net_1\, C => 
        \BEST_SEQCNT[3]_net_1\, Y => I2_un1_CO1);
    
    \REG40M.SEQCNTS_13[4]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[4]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_1, E => N_320, Q => \SEQCNTS_13[4]\);
    
    \REG40M.BIT_OS_VAL_5[0]\ : DFN1E1C0
      port map(D => N_282, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_1, E => \DES_SM_0[6]_net_1\, Q => 
        \BIT_OS_VAL_5[0]\);
    
    \ARB_BYTE[13]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[13]_net_1\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_32_0, Q => 
        \ARB_BYTE[13]_net_1\);
    
    \BEST_BIT_OS_VAL_RNO_1[3]\ : MX2
      port map(A => N_3905, B => N_3929, S => 
        \INDEX_CNT[4]_net_1\, Y => N_3933);
    
    \CLKPHASE_RNI8NA33[2]\ : MX2
      port map(A => N_3695, B => N_3707, S => \CLKPHASE[2]_net_1\, 
        Y => N_3711);
    
    \WAITCNT_RNO[10]\ : XA1C
      port map(A => \WAITCNT[10]_net_1\, B => N_5781, C => N_4539, 
        Y => N_5811);
    
    \REG40M.BIT_OS_CNT_6_RNO[8]\ : XA1C
      port map(A => \BIT_OS_CNT_6[8]\, B => N_419, C => N_4530_2, 
        Y => N_5632);
    
    \CLKPHASE_RNIP0JI_1[2]\ : NOR3A
      port map(A => N_212, B => \CLKPHASE[2]_net_1\, C => 
        \CLKPHASE[1]_net_1\, Y => \un36_n_bit_os_val[15]\);
    
    \REG40M.BIT_OS_VAL_5_RNO[2]\ : MX2
      port map(A => \BIT_OS_VAL_5[2]\, B => N_781, S => 
        \un36_n_bit_os_val[26]\, Y => N_207);
    
    \REG40M.BIT_OS_VAL_27_RNIM99C[2]\ : MX2
      port map(A => \BIT_OS_VAL_11[2]\, B => \BIT_OS_VAL_27[2]\, 
        S => \CLKPHASE_5[4]_net_1\, Y => N_3617);
    
    \REG40M.BIT_OS_CNT_6_RNO_0[3]\ : NOR2A
      port map(A => N_430, B => \BIT_OS_CNT_6[3]\, Y => N_524);
    
    \REG40M.BIT_OS_CNT_3_RNO[5]\ : XA1B
      port map(A => BIT_OS_CNT_3_c4, B => \BIT_OS_CNT_3[5]\, C
         => N_4530_1, Y => BIT_OS_CNT_3_n5);
    
    \REG40M.BIT_OS_CNT_2_RNO_0[8]\ : NOR2B
      port map(A => \BIT_OS_CNT_2[7]\, B => BIT_OS_CNT_2_c6, Y
         => BIT_OS_CNT_2_260_0);
    
    \MAX_CNT_RNO[6]\ : XA1C
      port map(A => \MAX_CNT[6]_net_1\, B => N_388, C => 
        un1_DES_SM_19, Y => N_5634);
    
    \CLKPHASE_2_RNIO5FE1[3]\ : MX2
      port map(A => N_3628, B => N_3632, S => 
        \CLKPHASE_2[3]_net_1\, Y => N_3636);
    
    un1_CLKPHASE_I_22 : XOR2
      port map(A => \CLKPHASE[2]_net_1\, B => 
        \DWACT_ADD_CI_0_g_array_1[0]\, Y => I_22);
    
    \REG40M.BIT_OS_CNT_6_RNO[5]\ : NOR3A
      port map(A => N_387, B => BIT_OS_CNT_6_n5_i_0, C => 
        N_4530_1, Y => N_77);
    
    \INDEX_CNT_RNIHBBG2[3]\ : MX2
      port map(A => N_4071, B => N_4076, S => 
        \INDEX_CNT[3]_net_1\, Y => N_4081);
    
    \REG40M.BIT_OS_VAL_31[0]\ : DFN1E1C0
      port map(D => N_210, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_20, E => \DES_SM_4[6]_net_1\, Q => 
        \BIT_OS_VAL_31[0]\);
    
    \DES_SM_RNI74OM_0[7]\ : NOR3B
      port map(A => \DES_SM[7]_net_1\, B => \ARB_BYTE[6]_net_1\, 
        C => \ARB_BYTE[7]_net_1\, Y => N_562_3);
    
    \REG40M.SEQCNTS_5_RNI0M5U[3]\ : MX2
      port map(A => \SEQCNTS_5[3]\, B => \SEQCNTS_6[3]\, S => 
        \INDEX_CNT_2[0]_net_1\, Y => N_4016);
    
    \CLKPHASE_0_RNI966J5[1]\ : MX2
      port map(A => N_3625, B => N_3653, S => 
        \CLKPHASE_0[1]_net_1\, Y => N_3657);
    
    \REG40M.BIT_OS_CNT_3_RNISV481[2]\ : OR3
      port map(A => N_BIT_OS_VAL_3114lt8, B => 
        N_BIT_OS_VAL_3114lto8_1, C => N_BIT_OS_VAL_3114lto8_2, Y
         => N_BIT_OS_VAL_3114);
    
    \DES_SM_RNI5G18[7]\ : NOR2
      port map(A => \DES_SM[7]_net_1\, B => \DES_SM_1[8]_net_1\, 
        Y => N_558);
    
    \RECD_SER_WORD_RNO_6[1]\ : OA1
      port map(A => \BIT_OS_SEL[3]_net_1\, B => 
        n_recd_ser_word164, C => \ARB_BYTE[1]_net_1\, Y => 
        \ARB_BYTE_m_0[1]\);
    
    \REG40M.SEQCNTS_30_RNIPBVA[0]\ : MX2
      port map(A => \SEQCNTS_14[0]\, B => \SEQCNTS_30[0]\, S => 
        \CLKPHASE[4]_net_1\, Y => N_3853);
    
    \REG40M.BIT_OS_CNT_4[5]\ : DFN1E1C0
      port map(D => N_5622, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_9, E => BIT_OS_CNT_4e, Q => 
        \BIT_OS_CNT_4[5]\);
    
    \RECD_SER_WORD_RNICS6E1[1]\ : NOR3C
      port map(A => \RECD_SER_WORD[1]_net_1\, B => 
        \RECD_SER_WORD[2]_net_1\, C => TFC_SYNC_DET_1_2, Y => 
        TFC_SYNC_DET_1_4);
    
    \REG40M.SEQCNTS_13_RNIJEFE[1]\ : MX2
      port map(A => \SEQCNTS_13[1]\, B => \SEQCNTS_29[1]\, S => 
        \CLKPHASE_2[4]_net_1\, Y => N_3779);
    
    \REG40M.BIT_OS_VAL_23_RNO[1]\ : MX2B
      port map(A => \BIT_OS_VAL_23[1]\, B => N_206, S => 
        \un36_n_bit_os_val[8]\, Y => \N_BIT_OS_VAL_23_18[1]\);
    
    \INDEX_CNT_0_RNI3DKU1[3]\ : MX2
      port map(A => N_3999, B => N_4004, S => 
        \INDEX_CNT_0[3]_net_1\, Y => N_4009);
    
    \BIT_OS_SEL_RNINMQF[1]\ : NOR2B
      port map(A => \BIT_OS_SEL[0]_net_1\, B => 
        \BIT_OS_SEL[1]_net_1\, Y => n_recd_ser_word167_1);
    
    \DES_SM_RNIK5SE[8]\ : OR2
      port map(A => \DES_SM[8]_net_1\, B => \DES_SM[6]_net_1\, Y
         => N_4530);
    
    \REG40M.BIT_OS_VAL_14_RNO[3]\ : MX2
      port map(A => N_209, B => \BIT_OS_VAL_14[3]\, S => N_5673, 
        Y => \N_BIT_OS_VAL_14_18[3]\);
    
    \REG40M.BIT_OS_CNT_3_RNO[0]\ : NOR2
      port map(A => \BIT_OS_CNT_3[0]\, B => N_4530, Y => N_5619);
    
    \BEST_BIT_OS_VAL_RNO_23[3]\ : MX2
      port map(A => \BIT_OS_VAL_11[3]\, B => \BIT_OS_VAL_12[3]\, 
        S => \INDEX_CNT_1[0]_net_1\, Y => N_3941);
    
    \BEST_BIT_OS_VAL_RNO_18[0]\ : MX2
      port map(A => \BIT_OS_VAL_13[0]\, B => \BIT_OS_VAL_14[0]\, 
        S => \INDEX_CNT_2[0]_net_1\, Y => N_3894);
    
    \WAITCNT_RNIJOAR3[7]\ : NOR3B
      port map(A => \WAITCNT[7]_net_1\, B => 
        \DES_SM_ns_0_0_0_a2_4[0]\, C => N_5777, Y => N_5859);
    
    \BIT_OS_SEL[3]\ : DFN1C0
      port map(D => \BEST_BIT_OS_VAL[3]_net_1\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_27_1, Q => \BIT_OS_SEL[3]_net_1\);
    
    \INDEX_CNT_2_RNIJ1AR1[3]\ : MX2
      port map(A => N_4084, B => N_4089, S => 
        \INDEX_CNT_2[3]_net_1\, Y => N_4094);
    
    \ARB_BYTE[14]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[14]_net_1\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_33, Q => 
        \ARB_BYTE[14]_net_1\);
    
    \REG40M.BIT_OS_CNT_4_RNICVO86[4]\ : AO1A
      port map(A => N_BIT_OS_VAL_3118, B => N_82, C => 
        N_BIT_OS_VAL_3122, Y => N_84);
    
    \REG40M.BIT_OS_VAL_1[0]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_1_18[0]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_17, E => \DES_SM_3[6]_net_1\, Q
         => \BIT_OS_VAL_1[0]\);
    
    \CLKPHASE_RNIP0JI[2]\ : OR3
      port map(A => \CLKPHASE[2]_net_1\, B => N_80, C => 
        \CLKPHASE[1]_net_1\, Y => N_5679);
    
    \CLKPHASE_RNICT4B[0]\ : NOR2B
      port map(A => N_5072_2, B => \CLKPHASE[0]_net_1\, Y => 
        N_214);
    
    \BEST_BIT_OS_VAL_RNO_8[3]\ : MX2
      port map(A => N_3893, B => N_3897, S => 
        \INDEX_CNT_1[3]_net_1\, Y => N_3901);
    
    \CLKPHASE_2_RNIVV521[3]\ : MX2
      port map(A => N_3799, B => N_3804, S => 
        \CLKPHASE_2[3]_net_1\, Y => N_3809);
    
    \WAITCNT_RNIPLQI[2]\ : OR2A
      port map(A => \WAITCNT[2]_net_1\, B => N_5772, Y => N_5773);
    
    \REG40M.BIT_OS_CNT_5[5]\ : DFN1E1C0
      port map(D => N_5627, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_11, E => BIT_OS_CNT_5e, Q => 
        \BIT_OS_CNT_5[5]\);
    
    \INDEX_CNT_RNIQU2N4[2]\ : MX2
      port map(A => N_4080, B => N_4095, S => 
        \INDEX_CNT[2]_net_1\, Y => N_4100);
    
    \RECD_SER_WORD[3]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[3]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_29, Q => \RECD_SER_WORD[3]_net_1\);
    
    CONFIG_ONCE_TRIG_RNO_0 : NOR2A
      port map(A => \DES_SM_i_0[5]\, B => \DES_SM[1]_net_1\, Y
         => N_CONFIG_ONCE_TRIG_i_a3_0);
    
    \ARB_WRD_40M_FIXED[11]\ : DFN1C0
      port map(D => \Q[11]_net_1\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_28, Q => \ARB_WRD_40M_FIXED[11]_net_1\);
    
    \REG40M.BIT_OS_VAL_2[3]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_2_18[3]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_18, E => \DES_SM_4[6]_net_1\, Q
         => \BIT_OS_VAL_2[3]\);
    
    \CLKPHASE_1_RNIBEK8H7[2]\ : AO1
      port map(A => \un36_n_bit_os_val[13]\, B => N_782, C => 
        N_717, Y => N_310);
    
    \BEST_BIT_OS_VAL_RNO_29[2]\ : MX2
      port map(A => \BIT_OS_VAL_31[2]\, B => \BIT_OS_VAL_0[2]\, S
         => \INDEX_CNT_3[0]_net_1\, Y => N_3980);
    
    \REG40M.BIT_OS_CNT_7_RNIVNPI[0]\ : NOR2B
      port map(A => \BIT_OS_CNT_7[0]\, B => \BIT_OS_CNT_7[1]\, Y
         => BIT_OS_CNT_7_c1);
    
    \ARB_BYTE[7]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[7]_net_1\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_27, Q => 
        \ARB_BYTE[7]_net_1\);
    
    \REG40M.BIT_OS_VAL_20_RNIU0HQ[2]\ : MX2
      port map(A => \BIT_OS_VAL_4[2]\, B => \BIT_OS_VAL_20[2]\, S
         => \CLKPHASE_2[4]_net_1\, Y => N_3673);
    
    \BEST_BIT_OS_VAL_RNO_15[3]\ : MX2
      port map(A => \BIT_OS_VAL_1[3]\, B => \BIT_OS_VAL_2[3]\, S
         => \INDEX_CNT_0[0]_net_1\, Y => N_3881);
    
    \MAX_CNT[3]\ : DFN1E0C0
      port map(D => N_5637, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_16, E => N_558, Q => \MAX_CNT[3]_net_1\);
    
    \CLKPHASE_RNIAB7UH7[1]\ : AO1A
      port map(A => N_5675, B => N_782_0, C => N_717_0, Y => 
        N_340);
    
    \REG40M.BIT_OS_VAL_7[3]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_7_18[3]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_3, E => \DES_SM_1[6]_net_1\, Q
         => \BIT_OS_VAL_7[3]\);
    
    \REG40M.SEQCNTS_10_RNIARH31[1]\ : MX2
      port map(A => \SEQCNTS_9[1]\, B => \SEQCNTS_10[1]\, S => 
        \INDEX_CNT_1[0]_net_1\, Y => N_4004);
    
    \Q[12]\ : DFN1C0
      port map(D => \ADJ_Q[12]_net_1\, CLK => CCC_160M_FXD, CLR
         => P_MASTER_POR_B_c_23, Q => \Q[12]_net_1\);
    
    \BEST_BIT_OS_VAL_RNO_8[0]\ : MX2
      port map(A => N_3890, B => N_3894, S => 
        \INDEX_CNT_1[3]_net_1\, Y => N_3898);
    
    \RECD_SER_WORD_RNO_3[3]\ : NOR3C
      port map(A => n_recd_ser_word167_1, B => 
        n_recd_ser_word171_0, C => \ARB_BYTE[10]_net_1\, Y => 
        \ARB_BYTE_m[10]\);
    
    \BEST_BIT_OS_VAL_RNO_21[3]\ : MX2
      port map(A => \BIT_OS_VAL_21[3]\, B => \BIT_OS_VAL_22[3]\, 
        S => \INDEX_CNT[0]_net_1\, Y => N_3921);
    
    \ARB_BYTE_RNIAIJU_1[2]\ : NOR3A
      port map(A => N_772, B => \ARB_BYTE[5]_net_1\, C => 
        \ARB_BYTE[2]_net_1\, Y => BIT_OS_CNT_5lde_0_a3_1);
    
    \REG40M.BIT_OS_VAL_5_RNO[0]\ : MX2
      port map(A => \BIT_OS_VAL_5[0]\, B => N_5666, S => 
        \un36_n_bit_os_val[26]\, Y => N_282);
    
    \REG40M.BIT_OS_VAL_15[2]\ : DFN1E1C0
      port map(D => N_191, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_15, E => \DES_SM_2[6]_net_1\, Q => 
        \BIT_OS_VAL_15[2]\);
    
    \CLKPHASE_RNIG15B[0]\ : OR2
      port map(A => N_5663, B => \CLKPHASE[0]_net_1\, Y => N_80);
    
    \ARB_WRD_40M_FIXED[12]\ : DFN1C0
      port map(D => \Q[12]_net_1\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_28, Q => \ARB_WRD_40M_FIXED[12]_net_1\);
    
    \ARB_WRD_40M_FIXED[6]\ : DFN1C0
      port map(D => \Q[6]_net_1\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_26, Q => \ARB_WRD_40M_FIXED[6]_net_1\);
    
    \CLKPHASE_1[2]\ : DFN1C0
      port map(D => \TUNE_CLKPHASE_RNIDA643[2]_net_1\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_24_0, Q => 
        \CLKPHASE_1[2]_net_1\);
    
    \BEST_BIT_OS_VAL_RNO_6[0]\ : MX2
      port map(A => N_3970, B => N_3982, S => 
        \INDEX_CNT[2]_net_1\, Y => N_3986);
    
    ADJ_SER_IN_R_0DEL_RNO : MX2
      port map(A => TFC_IN_R, B => ELK0_IN_R, S => DCB_SALT_SEL_c, 
        Y => SER_RX_IN_R);
    
    \CLKPHASE_1_RNI9EF92[2]\ : MX2
      port map(A => N_3736, B => N_3751, S => 
        \CLKPHASE_1[2]_net_1\, Y => N_3756);
    
    \REG40M.SEQCNTS_24[1]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[1]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_8, E => N_298, Q => \SEQCNTS_24[1]\);
    
    \REG40M.SEQCNTS_10[0]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[0]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_18, E => N_326, Q => \SEQCNTS_10[0]\);
    
    \REG40M.SEQCNTS_17_RNI140L[0]\ : MX2
      port map(A => \SEQCNTS_17[0]\, B => \SEQCNTS_18[0]\, S => 
        \INDEX_CNT_3[0]_net_1\, Y => N_4033);
    
    \REG40M.BIT_OS_VAL_11_RNO[3]\ : MX2
      port map(A => \BIT_OS_VAL_11[3]\, B => N_209_0, S => 
        \un36_n_bit_os_val[20]\, Y => \N_BIT_OS_VAL_11_18[3]\);
    
    \BEST_BIT_OS_VAL_RNO_27[0]\ : MX2
      port map(A => \BIT_OS_VAL_27[0]\, B => \BIT_OS_VAL_28[0]\, 
        S => \INDEX_CNT_1[0]_net_1\, Y => N_3966);
    
    \DES_SM_RNII3SE[4]\ : NOR2
      port map(A => \DES_SM[4]_net_1\, B => \DES_SM[8]_net_1\, Y
         => N_5149);
    
    \BEST_BIT_OS_VAL_RNO_3[0]\ : MX2
      port map(A => N_3886, B => N_3898, S => 
        \INDEX_CNT_0[2]_net_1\, Y => N_3902);
    
    \REG40M.BIT_OS_CNT_5_RNIOHKL[8]\ : OR3
      port map(A => \BIT_OS_CNT_5[4]\, B => \BIT_OS_CNT_5[5]\, C
         => \BIT_OS_CNT_5[8]\, Y => N_BIT_OS_VAL_3122lto8_0_o3_2);
    
    \RECD_SER_WORD_RNO_8[3]\ : NOR3C
      port map(A => n_recd_ser_word165_2, B => 
        n_recd_ser_word167_1, C => \ARB_BYTE[6]_net_1\, Y => 
        \ARB_BYTE_m_2[6]\);
    
    \ARB_BYTE[12]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[12]_net_1\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_32_0, Q => 
        \ARB_BYTE[12]_net_1\);
    
    \REG40M.BIT_OS_CNT_0_RNI0EVB3[1]\ : NOR2A
      port map(A => N_BIT_OS_VAL_14_18_3_0_a2_0, B => N_445, Y
         => N_BIT_OS_VAL_14_18_3_0_a2_1);
    
    \BEST_BIT_OS_VAL_RNO_27[2]\ : MX2
      port map(A => \BIT_OS_VAL_27[2]\, B => \BIT_OS_VAL_28[2]\, 
        S => \INDEX_CNT_1[0]_net_1\, Y => N_3968);
    
    \REG40M.SEQCNTS_15_RNIESS9[2]\ : MX2
      port map(A => \SEQCNTS_31[2]\, B => \SEQCNTS_15[2]\, S => 
        \CLKPHASE_0[4]_net_1\, Y => N_3725);
    
    \REG40M.BIT_OS_VAL_14[3]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_14_18[3]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_13, E => \DES_SM_2[6]_net_1\, Q
         => \BIT_OS_VAL_14[3]\);
    
    \CLKPHASE_RNI8DDI1[3]\ : MX2
      port map(A => N_3614, B => N_3618, S => \CLKPHASE[3]_net_1\, 
        Y => N_3622);
    
    \CLKPHASE_1_RNIP06B1[3]\ : MX2
      port map(A => N_3661, B => N_3665, S => 
        \CLKPHASE_1[3]_net_1\, Y => N_3669);
    
    \REG40M.BIT_OS_VAL_24_RNO[3]\ : MX2
      port map(A => \BIT_OS_VAL_24[3]\, B => N_209, S => 
        \un36_n_bit_os_val[7]\, Y => \N_BIT_OS_VAL_24_18[3]\);
    
    \CLKPHASE_0_RNILI401[3]\ : MX2
      port map(A => N_3850, B => N_3855, S => 
        \CLKPHASE_0[3]_net_1\, Y => N_3860);
    
    \INDEX_CNT_RNI5AVH7[4]\ : MX2
      port map(A => N_4030, B => N_4060, S => 
        \INDEX_CNT[4]_net_1\, Y => N_4065);
    
    \REG40M.BIT_OS_VAL_6_RNO[3]\ : MX2
      port map(A => N_209, B => \BIT_OS_VAL_6[3]\, S => N_5677, Y
         => \N_BIT_OS_VAL_6_18[3]\);
    
    \DES_SM_RNIL3LTN[6]\ : NOR3B
      port map(A => un1_DES_SM_1034_i_a2_4_0, B => 
        \un107_bit_os_val[1]\, C => \un107_bit_os_val[3]\, Y => 
        un1_DES_SM_1034_i_a2_4_2);
    
    \ARB_WRD_40M_FIXED[7]\ : DFN1C0
      port map(D => \Q[7]_net_1\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_26, Q => \ARB_WRD_40M_FIXED[7]_net_1\);
    
    \TUNE_CLKPHASE_RNILF0P2[3]\ : AO1A
      port map(A => N_5780, B => \TUNE_CLKPHASE[3]_net_1\, C => 
        N_5795, Y => \TUNE_CLKPHASE_RNILF0P2[3]_net_1\);
    
    \RECD_SER_WORD_RNIVOFI[5]\ : NOR2
      port map(A => \RECD_SER_WORD[5]_net_1\, B => 
        \RECD_SER_WORD[6]_net_1\, Y => TFC_SYNC_DET_1_1);
    
    \REG40M.BIT_OS_CNT_4_RNI66IU[4]\ : OR2A
      port map(A => \BIT_OS_CNT_4[4]\, B => N_379, Y => N_382);
    
    ADJ_SER_IN_R_0DEL : DFN1C0
      port map(D => SER_RX_IN_R, CLK => CCC_160M_ADJ, CLR => 
        P_MASTER_POR_B_c_26, Q => \ADJ_SER_IN_R_0DEL\);
    
    \INDEX_CNT_RNIKPVH7[4]\ : MX2
      port map(A => N_4031, B => N_4061, S => 
        \INDEX_CNT[4]_net_1\, Y => N_4066);
    
    \ARB_WRD_40M_FIXED[2]\ : DFN1C0
      port map(D => \Q[2]_net_1\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_26, Q => \ARB_WRD_40M_FIXED[2]_net_1\);
    
    \REG40M.BIT_OS_CNT_6_RNIGFTO[3]\ : OR3C
      port map(A => \BIT_OS_CNT_6[1]\, B => \BIT_OS_CNT_6[2]\, C
         => \BIT_OS_CNT_6[3]\, Y => N_365);
    
    \REG40M.BIT_OS_CNT_2[2]\ : DFN1E1C0
      port map(D => BIT_OS_CNT_2_n2, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_5, E => BIT_OS_CNT_2e, Q => 
        \BIT_OS_CNT_2[2]\);
    
    \RECD_SER_WORD_RNO_7[1]\ : AO1
      port map(A => \ARB_BYTE[2]_net_1\, B => n_recd_ser_word165, 
        C => \ARB_BYTE_m_0[4]\, Y => \N_RECD_SER_WORD_iv_3[1]\);
    
    \DES_SM_RNO_1[4]\ : NOR2A
      port map(A => \DES_SM[6]_net_1\, B => \CLKPHASE[0]_net_1\, 
        Y => DES_SM_tr7_0);
    
    \REG40M.SEQCNTS_21_RNIT84E[2]\ : MX2
      port map(A => \SEQCNTS_5[2]\, B => \SEQCNTS_21[2]\, S => 
        \CLKPHASE_1[4]_net_1\, Y => N_3775);
    
    \BEST_BIT_OS_VAL_RNO_20[2]\ : MX2
      port map(A => \BIT_OS_VAL_25[2]\, B => \BIT_OS_VAL_26[2]\, 
        S => \INDEX_CNT_3[0]_net_1\, Y => N_3912);
    
    \REG40M.SEQCNTS_24[4]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[4]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_8, E => N_298, Q => \SEQCNTS_24[4]\);
    
    \REG40M.SEQCNTS_28[3]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[3]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_15, E => N_290, Q => \SEQCNTS_28[3]\);
    
    \REG40M.BIT_OS_VAL_10[0]\ : DFN1E1C0
      port map(D => N_270, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_6, E => \DES_SM_1[6]_net_1\, Q => 
        \BIT_OS_VAL_10[0]\);
    
    \REG40M.BIT_OS_VAL_3[1]\ : DFN1E1C0
      port map(D => N_5659, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_19, E => \DES_SM_4[6]_net_1\, Q => 
        \BIT_OS_VAL_3[1]\);
    
    \REG40M.BIT_OS_CNT_7_RNI9KDO1[5]\ : NOR2B
      port map(A => BIT_OS_CNT_7_c4, B => \BIT_OS_CNT_7[5]\, Y
         => BIT_OS_CNT_7_c5);
    
    \DES_SM_RNID9Q61[6]\ : NOR2B
      port map(A => \DES_SM[6]_net_1\, B => N_BIT_OS_VAL_3110, Y
         => un1_DES_SM_1034_i_a2_4_0);
    
    \REG40M.SEQCNTS_21_RNIP44E[0]\ : MX2
      port map(A => \SEQCNTS_5[0]\, B => \SEQCNTS_21[0]\, S => 
        \CLKPHASE_1[4]_net_1\, Y => N_3773);
    
    \REG40M.SEQCNTS_31_RNIEM4I[1]\ : NOR2A
      port map(A => \SEQCNTS_31[1]\, B => \INDEX_CNT[0]_net_1\, Y
         => N_4124);
    
    \RECD_SER_WORD_RNO[2]\ : OR3
      port map(A => \N_RECD_SER_WORD_iv_1[2]\, B => 
        \N_RECD_SER_WORD_iv_0[2]\, C => \N_RECD_SER_WORD_iv_5[2]\, 
        Y => \N_RECD_SER_WORD[2]\);
    
    \CLKPHASE_0_RNI3MOR[3]\ : MX2
      port map(A => N_3725, B => N_3730, S => 
        \CLKPHASE_0[3]_net_1\, Y => N_3735);
    
    \REG40M.BIT_OS_VAL_19[3]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_19_18[3]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_20, E => \DES_SM[6]_net_1\, Q => 
        \BIT_OS_VAL_19[3]\);
    
    \BEST_BIT_OS_VAL_RNO_2[3]\ : MX2
      port map(A => N_3961, B => N_3989, S => 
        \INDEX_CNT[4]_net_1\, Y => N_3993);
    
    \REG40M.BIT_OS_VAL_6_RNO[0]\ : MX2
      port map(A => N_5666_0, B => \BIT_OS_VAL_6[0]\, S => N_5677, 
        Y => \N_BIT_OS_VAL_6_18[0]\);
    
    \INDEX_CNT_RNI5VAG2[3]\ : MX2
      port map(A => N_4068, B => N_4073, S => 
        \INDEX_CNT[3]_net_1\, Y => N_4078);
    
    \BIT_OS_SEL_1[1]\ : DFN1C0
      port map(D => \BEST_BIT_OS_VAL[1]_net_1\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_27_0, Q => 
        \BIT_OS_SEL_1[1]_net_1\);
    
    \REG40M.SEQCNTS_21_RNITD7G[3]\ : MX2
      port map(A => \SEQCNTS_21[3]\, B => \SEQCNTS_22[3]\, S => 
        \INDEX_CNT_3[0]_net_1\, Y => N_4051);
    
    \BIT_OS_SEL_3[1]\ : DFN1C0
      port map(D => \BEST_BIT_OS_VAL[1]_net_1\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_27_0, Q => BIT_OS_SEL_3(1));
    
    \BEST_BIT_OS_VAL_RNO_24[2]\ : MX2
      port map(A => \BIT_OS_VAL_7[2]\, B => \BIT_OS_VAL_8[2]\, S
         => \INDEX_CNT_2[0]_net_1\, Y => N_3948);
    
    \REG40M.BIT_OS_CNT_6[3]\ : DFN1E1C0
      port map(D => N_81, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_12, E => BIT_OS_CNT_6e, Q => 
        \BIT_OS_CNT_6[3]\);
    
    \REG40M.BIT_OS_CNT_6[5]\ : DFN1E1C0
      port map(D => N_77, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_12, E => BIT_OS_CNT_6e, Q => 
        \BIT_OS_CNT_6[5]\);
    
    \REG40M.BIT_OS_VAL_13[0]\ : DFN1E1C0
      port map(D => N_261, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_12, E => \DES_SM_2[6]_net_1\, Q => 
        \BIT_OS_VAL_13[0]\);
    
    \REG40M.BIT_OS_CNT_0_RNIA565[5]\ : OR3
      port map(A => \BIT_OS_CNT_0[5]\, B => \BIT_OS_CNT_0[6]\, C
         => \BIT_OS_CNT_0[7]\, Y => N_BIT_OS_VAL_312lto8_0_o3_2);
    
    \DES_SM_RNID8OB[8]\ : NOR2A
      port map(A => \DES_SM[8]_net_1\, B => OP_MODE_c_0, Y => 
        N_140);
    
    \CLKPHASE_RNI36QUE[0]\ : MX2
      port map(A => N_BIT_OS_VAL_3114, B => N_BIT_OS_VAL_3130, S
         => \un107_bit_os_val[2]\, Y => N_427);
    
    \REG40M.SEQCNTS_23_RNI0IDH[2]\ : MX2
      port map(A => \SEQCNTS_7[2]\, B => \SEQCNTS_23[2]\, S => 
        \CLKPHASE_0[4]_net_1\, Y => N_3730);
    
    \REG40M.BIT_OS_CNT_0[7]\ : DFN1E1C0
      port map(D => N_5639, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_3, E => BIT_OS_CNT_0e, Q => 
        \BIT_OS_CNT_0[7]\);
    
    \SYNC_SM.N_TUNE_CLKPHASE_2_0_0_ADD_5x5_slow_I2_S\ : XNOR3
      port map(A => \BEST_SEQCNT[3]_net_1\, B => 
        \BEST_CLKPHASE[2]_net_1\, C => N86, Y => 
        \N_TUNE_CLKPHASE_2[2]\);
    
    \REG40M.BIT_OS_VAL_6_RNO[2]\ : MX2
      port map(A => N_781_0, B => \BIT_OS_VAL_6[2]\, S => N_5677, 
        Y => N_5650);
    
    \REG40M.BIT_OS_VAL_30_RNIJTSP[3]\ : MX2
      port map(A => \BIT_OS_VAL_14[3]\, B => \BIT_OS_VAL_30[3]\, 
        S => \CLKPHASE_3[4]_net_1\, Y => N_3706);
    
    \REG40M.BIT_OS_VAL_21_RNO[3]\ : MX2
      port map(A => \BIT_OS_VAL_21[3]\, B => N_209, S => 
        \un36_n_bit_os_val[10]\, Y => \N_BIT_OS_VAL_21_18[3]\);
    
    \INDEX_CNT_RNITPS63[2]\ : MX2
      port map(A => N_4043, B => N_4053, S => 
        \INDEX_CNT[2]_net_1\, Y => N_4058);
    
    \REG40M.BIT_OS_VAL_16_RNO[3]\ : MX2
      port map(A => \BIT_OS_VAL_16[3]\, B => N_209_0, S => 
        \un36_n_bit_os_val[15]\, Y => \N_BIT_OS_VAL_16_18[3]\);
    
    \WAITCNT_RNO[13]\ : XA1C
      port map(A => \WAITCNT[13]_net_1\, B => N_5787, C => N_4539, 
        Y => WAITCNT_n13);
    
    \REG40M.SEQCNTS_31[2]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[2]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_10, E => N_284, Q => \SEQCNTS_31[2]\);
    
    \REG40M.SEQCNTS_27_RNID03Q[0]\ : MX2
      port map(A => \SEQCNTS_11[0]\, B => \SEQCNTS_27[0]\, S => 
        \CLKPHASE_2[4]_net_1\, Y => N_3743);
    
    \REG40M.SEQCNTS_25[4]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[4]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_10, E => N_296, Q => \SEQCNTS_25[4]\);
    
    \REG40M.SEQCNTS_23_RNI4MDH[4]\ : MX2
      port map(A => \SEQCNTS_7[4]\, B => \SEQCNTS_23[4]\, S => 
        \CLKPHASE_0[4]_net_1\, Y => N_3732);
    
    \REG40M.SEQCNTS_22_RNI3RMK[2]\ : MX2
      port map(A => \SEQCNTS_6[2]\, B => \SEQCNTS_22[2]\, S => 
        \CLKPHASE_5[4]_net_1\, Y => N_3850);
    
    \RECD_SER_WORD_RNO_2[5]\ : OR3
      port map(A => \ARB_BYTE_m_4[7]\, B => \ARB_BYTE_m_4[5]\, C
         => \N_RECD_SER_WORD_iv_3[5]\, Y => 
        \N_RECD_SER_WORD_iv_5[5]\);
    
    \REG40M.BIT_OS_VAL_31_RNO[0]\ : MX2
      port map(A => \BIT_OS_VAL_31[0]\, B => N_5666_0, S => 
        \un36_n_bit_os_val[0]\, Y => N_210);
    
    \DES_SM_RNIIU5J5[0]\ : AO1
      port map(A => un1_DES_SM_471_i_0_0_0_a3_0, B => N_116, C
         => un1_DES_SM_471_i_0_0_0_0, Y => 
        un1_DES_SM_471_i_0_0_0_1);
    
    \BIT_OS_SEL_1_RNI4GRD1[0]\ : NOR3
      port map(A => \BIT_OS_SEL_1[1]_net_1\, B => 
        \BIT_OS_SEL_1[0]_net_1\, C => \BIT_OS_SEL_1[2]_net_1\, Y
         => n_recd_ser_word164);
    
    \REG40M.SEQCNTS_25_RNI993P[3]\ : MX2
      port map(A => \SEQCNTS_9[3]\, B => \SEQCNTS_25[3]\, S => 
        \CLKPHASE_3[4]_net_1\, Y => N_3766);
    
    \DES_SM_RNICU2EH7_5[8]\ : AO1
      port map(A => \un36_n_bit_os_val[3]\, B => N_782, C => 
        N_717, Y => N_290);
    
    \BIT_OS_SEL_1_RNII4DE1[1]\ : NOR3C
      port map(A => \BIT_OS_SEL_1[2]_net_1\, B => 
        \BIT_OS_SEL_1[1]_net_1\, C => n_recd_ser_word170_0, Y => 
        n_recd_ser_word170);
    
    \RECD_SER_WORD_RNO_0[4]\ : AO1
      port map(A => \ARB_BYTE[10]_net_1\, B => n_recd_ser_word170, 
        C => \ARB_BYTE_m[11]\, Y => \N_RECD_SER_WORD_iv_1[4]\);
    
    \SYNC_SM.N_TUNE_CLKPHASE_2_0_0_ADD_5x5_slow_I4_Y\ : XNOR2
      port map(A => N90, B => \BEST_CLKPHASE[4]_net_1\, Y => N_1);
    
    \REG40M.BIT_OS_CNT_5[3]\ : DFN1E1C0
      port map(D => N_5629, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_11, E => BIT_OS_CNT_5e, Q => 
        \BIT_OS_CNT_5[3]\);
    
    \INDEX_CNT_0_RNIHOTE3[2]\ : MX2
      port map(A => N_4117, B => N_4132, S => 
        \INDEX_CNT_0[2]_net_1\, Y => N_4137);
    
    \CLKPHASE[0]\ : DFN1C0
      port map(D => \CLKPHASE_RNO[0]_net_1\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_24, Q => \CLKPHASE[0]_net_1\);
    
    \REG40M.BIT_OS_CNT_3_RNO_0[8]\ : NOR2B
      port map(A => \BIT_OS_CNT_3[7]\, B => BIT_OS_CNT_3_c6, Y
         => BIT_OS_CNT_3_432_0);
    
    \REG40M.SEQCNTS_29_RNI8CG41[3]\ : MX2
      port map(A => N_4051, B => \SEQCNTS_29[3]\, S => 
        \INDEX_CNT_2[3]_net_1\, Y => N_4056);
    
    \INDEX_CNT_RNI6DDH8[4]\ : MX2
      port map(A => N_4099, B => N_4134, S => 
        \INDEX_CNT[4]_net_1\, Y => N_4139);
    
    \REG40M.BIT_OS_CNT_7[2]\ : DFN1E1C0
      port map(D => BIT_OS_CNT_7_n2, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_14, E => BIT_OS_CNT_7e, Q => 
        \BIT_OS_CNT_7[2]\);
    
    \REG40M.SEQCNTS_31_RNIHP4I[4]\ : NOR2A
      port map(A => \SEQCNTS_31[4]\, B => \INDEX_CNT[0]_net_1\, Y
         => N_4127);
    
    \INDEX_CNT_RNI1BHU3[2]\ : MX2
      port map(A => N_4010, B => N_4025, S => 
        \INDEX_CNT[2]_net_1\, Y => N_4030);
    
    \REG40M.SEQCNTS_7_RNILL051[4]\ : MX2
      port map(A => \SEQCNTS_7[4]\, B => \SEQCNTS_8[4]\, S => 
        \INDEX_CNT[0]_net_1\, Y => N_4087);
    
    \REG40M.SEQCNTS_28[2]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[2]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_15, E => N_290, Q => \SEQCNTS_28[2]\);
    
    \REG40M.SEQCNTS_20[3]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[3]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_2, E => N_306, Q => \SEQCNTS_20[3]\);
    
    \REG40M.BIT_OS_VAL_10[3]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_10_18[3]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_6, E => \DES_SM_1[6]_net_1\, Q
         => \BIT_OS_VAL_10[3]\);
    
    ADJ_SER_IN_R_1DEL : DFN1C0
      port map(D => \ADJ_SER_IN_R_0DEL\, CLK => CCC_160M_ADJ, CLR
         => P_MASTER_POR_B_c_27_1, Q => \ADJ_SER_IN_R_1DEL\);
    
    \REG40M.SEQCNTS_21_RNIVF7G[4]\ : MX2
      port map(A => \SEQCNTS_21[4]\, B => \SEQCNTS_22[4]\, S => 
        \INDEX_CNT_3[0]_net_1\, Y => N_4052);
    
    \CLKPHASE_RNIVNJCG7_0[0]\ : OR3
      port map(A => un1_DES_SM_1034_i_o2_1, B => N_754, C => 
        un1_DES_SM_1034_i_o2_2, Y => N_782);
    
    \CLKPHASE_RNIP0JI_4[0]\ : NOR2A
      port map(A => N_212, B => N_90, Y => 
        \un36_n_bit_os_val[11]\);
    
    \REG40M.SEQCNTS_26[3]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[3]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_12, E => N_294, Q => \SEQCNTS_26[3]\);
    
    \RECD_SER_WORD_RNO_7[2]\ : AO1
      port map(A => \ARB_BYTE[3]_net_1\, B => n_recd_ser_word165, 
        C => \ARB_BYTE_m_1[5]\, Y => \N_RECD_SER_WORD_iv_3[2]\);
    
    \ARB_BYTE_RNI82M33[0]\ : AO1
      port map(A => BIT_OS_CNT_1lde_0_a3_2, B => 
        BIT_OS_CNT_1lde_0_a3_1, C => N_4530_0, Y => BIT_OS_CNT_1e);
    
    \REG40M.SEQCNTS_3[1]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[1]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_11, E => N_340, Q => \SEQCNTS_3[1]\);
    
    \REG40M.BIT_OS_CNT_3_RNI3C1A[6]\ : OR2
      port map(A => \BIT_OS_CNT_3[7]\, B => \BIT_OS_CNT_3[6]\, Y
         => N_BIT_OS_VAL_3114lto8_1);
    
    \DES_SM[3]\ : DFN1C0
      port map(D => \DES_SM_RNO[3]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_27, Q => \DES_SM[3]_net_1\);
    
    \REG40M.BIT_OS_CNT_6_RNO[0]\ : NOR2
      port map(A => \BIT_OS_CNT_6[0]\, B => N_4530, Y => N_527);
    
    \REG40M.BIT_OS_CNT_4_RNO[1]\ : XA1B
      port map(A => \BIT_OS_CNT_4[0]\, B => \BIT_OS_CNT_4[1]\, C
         => N_4530_0, Y => N_5624);
    
    \REG40M.BIT_OS_VAL_28_RNIFSV8[0]\ : MX2
      port map(A => \BIT_OS_VAL_12[0]\, B => \BIT_OS_VAL_28[0]\, 
        S => \CLKPHASE_0[4]_net_1\, Y => N_3675);
    
    \REG40M.SEQCNTS_9[3]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[3]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_20, E => N_328, Q => \SEQCNTS_9[3]\);
    
    \CLKPHASE_RNIP0JI[0]\ : NOR3B
      port map(A => \CLKPHASE[0]_net_1\, B => N_215, C => N_90, Y
         => \un36_n_bit_os_val[2]\);
    
    \RECD_SER_WORD_RNO_5[4]\ : NOR3C
      port map(A => n_recd_ser_word165_2, B => 
        n_recd_ser_word166_0, C => \ARB_BYTE[6]_net_1\, Y => 
        \ARB_BYTE_m_3[6]\);
    
    \ADJ_Q[6]\ : DFN1C0
      port map(D => \ADJ_Q[4]_net_1\, CLK => CCC_160M_ADJ, CLR
         => P_MASTER_POR_B_c_34_0, Q => \ADJ_Q[6]_net_1\);
    
    \REG40M.BIT_OS_CNT_7_RNO[2]\ : XA1B
      port map(A => BIT_OS_CNT_7_c1, B => \BIT_OS_CNT_7[2]\, C
         => N_4530_2, Y => BIT_OS_CNT_7_n2);
    
    \BEST_BIT_OS_VAL_RNO[0]\ : NOR2A
      port map(A => \N_BEST_BIT_OS_VAL_3[0]\, B => 
        \DES_SM[8]_net_1\, Y => \N_BEST_BIT_OS_VAL[0]\);
    
    \REG40M.BIT_OS_VAL_25[2]\ : DFN1E1C0
      port map(D => N_171, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_20, E => \DES_SM[6]_net_1\, Q => 
        \BIT_OS_VAL_25[2]\);
    
    \RECD_SER_WORD_RNO_8[5]\ : NOR3C
      port map(A => n_recd_ser_word165_2, B => 
        n_recd_ser_word167_1, C => \ARB_BYTE[8]_net_1\, Y => 
        \ARB_BYTE_m_3[8]\);
    
    \REG40M.BIT_OS_VAL_26_RNO[3]\ : MX2
      port map(A => \BIT_OS_VAL_26[3]\, B => N_209, S => 
        \un36_n_bit_os_val[5]\, Y => \N_BIT_OS_VAL_26_18[3]\);
    
    \CLKPHASE_0_RNIQL1G2[2]\ : MX2
      port map(A => N_3636, B => N_3648, S => 
        \CLKPHASE_0[2]_net_1\, Y => N_3652);
    
    \REG40M.SEQCNTS_10_RNI8PH31[0]\ : MX2
      port map(A => \SEQCNTS_9[0]\, B => \SEQCNTS_10[0]\, S => 
        \INDEX_CNT_1[0]_net_1\, Y => N_4003);
    
    \RECD_SER_WORD_RNO_8[2]\ : NOR3C
      port map(A => n_recd_ser_word165_2, B => 
        n_recd_ser_word167_1, C => \ARB_BYTE[5]_net_1\, Y => 
        \ARB_BYTE_m_1[5]\);
    
    \REG40M.SEQCNTS_24_RNI200O[0]\ : MX2
      port map(A => \SEQCNTS_8[0]\, B => \SEQCNTS_24[0]\, S => 
        \CLKPHASE_4[4]_net_1\, Y => N_3803);
    
    \REG40M.SEQCNTS_23[2]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[2]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_6, E => N_300, Q => \SEQCNTS_23[2]\);
    
    \RECD_SER_WORD_RNO_0[2]\ : AO1
      port map(A => \ARB_BYTE[8]_net_1\, B => n_recd_ser_word170, 
        C => \ARB_BYTE_m[9]\, Y => \N_RECD_SER_WORD_iv_1[2]\);
    
    \RECD_SER_WORD_RNO_1[1]\ : AO1
      port map(A => n_recd_ser_word168, B => \ARB_BYTE[5]_net_1\, 
        C => \ARB_BYTE_m_0[6]\, Y => \N_RECD_SER_WORD_iv_0[1]\);
    
    \BEST_BIT_OS_VAL_RNO_24[0]\ : MX2
      port map(A => \BIT_OS_VAL_7[0]\, B => \BIT_OS_VAL_8[0]\, S
         => \INDEX_CNT_2[0]_net_1\, Y => N_3946);
    
    \REG40M.BIT_OS_CNT_5[7]\ : DFN1E1C0
      port map(D => N_5625, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_11, E => BIT_OS_CNT_5e, Q => 
        \BIT_OS_CNT_5[7]\);
    
    \REG40M.BIT_OS_CNT_3[4]\ : DFN1E1C0
      port map(D => BIT_OS_CNT_3_n4, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_7, E => BIT_OS_CNT_3e, Q => 
        \BIT_OS_CNT_3[4]\);
    
    \RECD_SER_WORD_RNO_5[0]\ : NOR3C
      port map(A => n_recd_ser_word165_2, B => 
        n_recd_ser_word166_0, C => \ARB_BYTE[2]_net_1\, Y => 
        \ARB_BYTE_m[2]\);
    
    \CLKPHASE_0[2]\ : DFN1C0
      port map(D => \TUNE_CLKPHASE_RNIDA643[2]_net_1\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_24_0, Q => 
        \CLKPHASE_0[2]_net_1\);
    
    \REG40M.BIT_OS_VAL_31[2]\ : DFN1E1C0
      port map(D => N_159, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_20, E => \DES_SM_4[6]_net_1\, Q => 
        \BIT_OS_VAL_31[2]\);
    
    \REG40M.BIT_OS_CNT_4_RNIL8BI[4]\ : OR3
      port map(A => \BIT_OS_CNT_4[4]\, B => \BIT_OS_CNT_4[6]\, C
         => \BIT_OS_CNT_4[7]\, Y => N_BIT_OS_VAL_3118lto8_0_o3_2);
    
    \BEST_SEQCNT_RNO[4]\ : NOR2A
      port map(A => \un6_n_best_seqcnt[4]\, B => 
        \DES_SM[8]_net_1\, Y => \N_BEST_SEQCNT[4]\);
    
    \ARB_BYTE[6]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[6]_net_1\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_27, Q => 
        \ARB_BYTE[6]_net_1\);
    
    \RECD_SER_WORD_RNO_4[0]\ : NOR3C
      port map(A => n_recd_ser_word168_2, B => 
        n_recd_ser_word169_0, C => \ARB_BYTE[5]_net_1\, Y => 
        \ARB_BYTE_m[5]\);
    
    \REG40M.SEQCNTS_25_RNI333P[0]\ : MX2
      port map(A => \SEQCNTS_9[0]\, B => \SEQCNTS_25[0]\, S => 
        \CLKPHASE_3[4]_net_1\, Y => N_3763);
    
    \BEST_BIT_OS_VAL_RNO_10[0]\ : MX2
      port map(A => N_3918, B => \BIT_OS_VAL_29[0]\, S => 
        \INDEX_CNT[3]_net_1\, Y => N_3922);
    
    \BEST_BIT_OS_VAL_RNO_12[1]\ : MX2
      port map(A => N_3947, B => N_3951, S => 
        \INDEX_CNT_0[3]_net_1\, Y => N_3955);
    
    \REG40M.BIT_OS_VAL_8_RNO[1]\ : MX2B
      port map(A => \BIT_OS_VAL_8[1]\, B => N_206_0, S => 
        \un36_n_bit_os_val[23]\, Y => \N_BIT_OS_VAL_8_18[1]\);
    
    \REG40M.BIT_OS_CNT_7_RNO_0[8]\ : NOR2B
      port map(A => \BIT_OS_CNT_7[7]\, B => BIT_OS_CNT_7_c6, Y
         => BIT_OS_CNT_7_360_0);
    
    \RECD_SER_WORD[0]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[0]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_29, Q => \RECD_SER_WORD[0]_net_1\);
    
    \REG40M.SEQCNTS_16_RNI4GH7[1]\ : NOR2B
      port map(A => \SEQCNTS_16[1]\, B => \CLKPHASE[4]_net_1\, Y
         => N_3799);
    
    \REG40M.BIT_OS_VAL_24[3]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_24_18[3]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_18, E => \DES_SM_4[6]_net_1\, Q
         => \BIT_OS_VAL_24[3]\);
    
    \WAITCNT[7]\ : DFN1E0C0
      port map(D => N_5719, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_9, E => N_5790, Q => \WAITCNT[7]_net_1\);
    
    un1_CLKPHASE_I_23 : NOR2B
      port map(A => \DWACT_ADD_CI_0_TMP[0]\, B => 
        \CLKPHASE[1]_net_1\, Y => \DWACT_ADD_CI_0_g_array_1[0]\);
    
    \CLKPHASE_RNICU2EH7[0]\ : AO1
      port map(A => \un36_n_bit_os_val[10]\, B => N_782, C => 
        N_717, Y => N_304);
    
    \REG40M.SEQCNTS_31[4]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[4]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_10, E => N_284, Q => \SEQCNTS_31[4]\);
    
    \REG40M.BIT_OS_VAL_15_RNO[3]\ : MX2
      port map(A => \BIT_OS_VAL_15[3]\, B => N_209_0, S => 
        \un36_n_bit_os_val[16]\, Y => \N_BIT_OS_VAL_15_18[3]\);
    
    \Q[0]\ : DFN1C0
      port map(D => \ADJ_Q[0]_net_1\, CLK => CCC_160M_FXD, CLR
         => P_MASTER_POR_B_c_34, Q => \Q[0]_net_1\);
    
    \REG40M.SEQCNTS_14[0]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[0]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_2, E => N_318, Q => \SEQCNTS_14[0]\);
    
    \REG40M.BIT_OS_VAL_2_RNIU7QR[0]\ : MX2
      port map(A => \BIT_OS_VAL_2[0]\, B => \BIT_OS_VAL_18[0]\, S
         => \CLKPHASE_1[4]_net_1\, Y => N_3687);
    
    \REG40M.BIT_OS_CNT_5_RNO[5]\ : XA1C
      port map(A => \BIT_OS_CNT_5[5]\, B => N_384, C => N_4530, Y
         => N_5627);
    
    \REG40M.BIT_OS_CNT_1[4]\ : DFN1E1C0
      port map(D => N_133, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_4, E => BIT_OS_CNT_1e, Q => 
        \BIT_OS_CNT_1[4]\);
    
    \BEST_BIT_OS_VAL_RNO_19[3]\ : MX2
      port map(A => \BIT_OS_VAL_17[3]\, B => \BIT_OS_VAL_18[3]\, 
        S => \INDEX_CNT_3[0]_net_1\, Y => N_3909);
    
    \REG40M.SEQCNTS_7[4]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[4]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_18, E => N_332, Q => \SEQCNTS_7[4]\);
    
    \REG40M.SEQCNTS_19_RNI2NGG[2]\ : MX2
      port map(A => \SEQCNTS_3[2]\, B => \SEQCNTS_19[2]\, S => 
        \CLKPHASE_1[4]_net_1\, Y => N_3740);
    
    \BIT_OS_SEL_7[2]\ : DFN1C0
      port map(D => \BEST_BIT_OS_VAL[2]_net_1\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_27_0, Q => BIT_OS_SEL_7_0);
    
    \REG40M.SEQCNTS_16_RNI5HH7[2]\ : NOR2B
      port map(A => \SEQCNTS_16[2]\, B => \CLKPHASE[4]_net_1\, Y
         => N_3800);
    
    \REG40M.BIT_OS_CNT_2_RNIBPGN[5]\ : NOR2B
      port map(A => BIT_OS_CNT_2_c4, B => \BIT_OS_CNT_2[5]\, Y
         => BIT_OS_CNT_2_c5);
    
    \REG40M.SEQCNTS_10[1]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[1]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_18, E => N_326, Q => \SEQCNTS_10[1]\);
    
    \REG40M.BIT_OS_VAL_12[3]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_12_18[3]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_10, E => \DES_SM_2[6]_net_1\, Q
         => \BIT_OS_VAL_12[3]\);
    
    \REG40M.BIT_OS_VAL_5_RNIVB0G[0]\ : MX2
      port map(A => \BIT_OS_VAL_5[0]\, B => \BIT_OS_VAL_21[0]\, S
         => \CLKPHASE_5[4]_net_1\, Y => N_3639);
    
    \REG40M.BIT_OS_CNT_0_RNIG6E41[1]\ : NOR2
      port map(A => N_BIT_OS_VAL_312, B => N_BIT_OS_VAL_316, Y
         => N_BIT_OS_VAL_14_18_3_0_a2_0);
    
    \INDEX_CNT[3]\ : DFN1E0C0
      port map(D => \N_INDEX_CNT[3]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_17, E => N_5149, Q => 
        \INDEX_CNT[3]_net_1\);
    
    \DES_SM_RNI95TM[0]\ : NOR3
      port map(A => \DES_SM_1[8]_net_1\, B => \DES_SM[0]_net_1\, 
        C => N_5783, Y => N_5790);
    
    \CLKPHASE_0_RNI2STU[3]\ : MX2
      port map(A => N_3642, B => N_3646, S => 
        \CLKPHASE_0[3]_net_1\, Y => N_3650);
    
    \REG40M.SEQCNTS_1[2]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[2]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_8, E => N_344, Q => \SEQCNTS_1[2]\);
    
    \REG40M.BIT_OS_VAL_20[0]\ : DFN1E1C0
      port map(D => N_243, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_13, E => \DES_SM_2[6]_net_1\, Q => 
        \BIT_OS_VAL_20[0]\);
    
    \REG40M.BIT_OS_VAL_6_RNI0BTE[1]\ : MX2
      port map(A => \BIT_OS_VAL_6[1]\, B => \BIT_OS_VAL_22[1]\, S
         => \CLKPHASE_2[4]_net_1\, Y => N_3700);
    
    \DES_SM[5]\ : DFN1P0
      port map(D => \DES_SM_RNO[5]_net_1\, CLK => CLK_40M_GL, PRE
         => P_MASTER_POR_B_c_27, Q => \DES_SM_i_0[5]\);
    
    \RECD_SER_WORD_RNO_3[7]\ : NOR3C
      port map(A => n_recd_ser_word167_1, B => 
        n_recd_ser_word171_0, C => \ARB_BYTE[14]_net_1\, Y => 
        \ARB_BYTE_m[14]\);
    
    \CLKPHASE_2_RNIEQEB1[3]\ : MX2
      port map(A => N_3702, B => N_3706, S => 
        \CLKPHASE_2[3]_net_1\, Y => N_3710);
    
    \REG40M.BIT_OS_VAL_29[3]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_29_18[3]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_4, E => \DES_SM_1[6]_net_1\, Q
         => \BIT_OS_VAL_29[3]\);
    
    \REG40M.BIT_OS_VAL_30_RNO[0]\ : MX2
      port map(A => \BIT_OS_VAL_30[0]\, B => N_5666_0, S => 
        \un36_n_bit_os_val[1]\, Y => N_213);
    
    \RECD_SER_WORD_RNIB4H14[1]\ : NOR3C
      port map(A => ELK0_SYNC_DET_1_2, B => ELK0_SYNC_DET_1_1, C
         => ELK0_SYNC_DET_1_3, Y => ELK0_SYNC_DET_1);
    
    \BEST_BIT_OS_VAL_RNO_22[3]\ : MX2
      port map(A => \BIT_OS_VAL_3[3]\, B => \BIT_OS_VAL_4[3]\, S
         => \INDEX_CNT_0[0]_net_1\, Y => N_3937);
    
    \REG40M.SEQCNTS_20_RNIRAAG[0]\ : MX2
      port map(A => \SEQCNTS_4[0]\, B => \SEQCNTS_20[0]\, S => 
        \CLKPHASE_5[4]_net_1\, Y => N_3813);
    
    \REG40M.BIT_OS_VAL_1_RNIT0HO[1]\ : MX2
      port map(A => \BIT_OS_VAL_1[1]\, B => \BIT_OS_VAL_17[1]\, S
         => \CLKPHASE_0[4]_net_1\, Y => N_3628);
    
    \DES_SM_RNO_1[3]\ : NOR2A
      port map(A => \DES_SM_i_0[5]\, B => \DES_SM[3]_net_1\, Y
         => N_5813);
    
    \REG40M.SEQCNTS_30[2]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[2]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_7, E => N_286, Q => \SEQCNTS_30[2]\);
    
    \BEST_BIT_OS_VAL_RNO_29[0]\ : MX2
      port map(A => \BIT_OS_VAL_31[0]\, B => \BIT_OS_VAL_0[0]\, S
         => \INDEX_CNT_3[0]_net_1\, Y => N_3978);
    
    \ARB_BYTE[2]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[2]_net_1\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_27, Q => 
        \ARB_BYTE[2]_net_1\);
    
    \REG40M.BIT_OS_VAL_23[0]\ : DFN1E1C0
      port map(D => N_234, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_17_0, E => \DES_SM_3[6]_net_1\, Q => 
        \BIT_OS_VAL_23[0]\);
    
    \REG40M.SEQCNTS_19[2]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[2]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_11, E => N_308, Q => \SEQCNTS_19[2]\);
    
    \REG40M.BIT_OS_CNT_7_RNO[7]\ : XA1B
      port map(A => BIT_OS_CNT_7_c6, B => \BIT_OS_CNT_7[7]\, C
         => N_4530_2, Y => BIT_OS_CNT_7_n7);
    
    \REG40M.BIT_OS_CNT_7_RNIGL6S[2]\ : NOR2B
      port map(A => BIT_OS_CNT_7_c1, B => \BIT_OS_CNT_7[2]\, Y
         => BIT_OS_CNT_7_c2);
    
    \REG40M.SEQCNTS_20[4]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[4]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_2, E => N_306, Q => \SEQCNTS_20[4]\);
    
    \BEST_BIT_OS_VAL_RNO_13[2]\ : MX2
      port map(A => N_3964, B => N_3968, S => 
        \INDEX_CNT_1[3]_net_1\, Y => N_3972);
    
    \CLKPHASE_1_RNIHMF92[2]\ : MX2
      port map(A => N_3737, B => N_3752, S => 
        \CLKPHASE_1[2]_net_1\, Y => N_3757);
    
    \BEST_BIT_OS_VAL_RNO_11[2]\ : MX2
      port map(A => N_3936, B => N_3940, S => 
        \INDEX_CNT_0[3]_net_1\, Y => N_3944);
    
    \REG40M.BIT_OS_VAL_9[2]\ : DFN1E1C0
      port map(D => N_201, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_6, E => \DES_SM_1[6]_net_1\, Q => 
        \BIT_OS_VAL_9[2]\);
    
    \ARB_BYTE_RNICT161_0[1]\ : NOR3B
      port map(A => \ARB_BYTE[1]_net_1\, B => N_559_1, C => 
        \ARB_BYTE[4]_net_1\, Y => BIT_OS_CNT_6lde_0_a3_1);
    
    \REG40M.SEQCNTS_23_RNISDDH[0]\ : MX2
      port map(A => \SEQCNTS_7[0]\, B => \SEQCNTS_23[0]\, S => 
        \CLKPHASE_0[4]_net_1\, Y => N_3728);
    
    \REG40M.BIT_OS_CNT_4_RNI0IBO7_0[4]\ : OR2
      port map(A => N_360, B => N_437, Y => N_781_0);
    
    \REG40M.BIT_OS_VAL_14[2]\ : DFN1E1C0
      port map(D => N_5649, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_13, E => \DES_SM_2[6]_net_1\, Q => 
        \BIT_OS_VAL_14[2]\);
    
    \BIT_OS_SEL[0]\ : DFN1C0
      port map(D => \BEST_BIT_OS_VAL[0]_net_1\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_27_1, Q => \BIT_OS_SEL[0]_net_1\);
    
    \CLKPHASE_1_RNI2PL82[2]\ : MX2
      port map(A => N_3771, B => N_3786, S => 
        \CLKPHASE_1[2]_net_1\, Y => N_3791);
    
    \CLKPHASE_RNID3E7_0[3]\ : NOR2B
      port map(A => \CLKPHASE[3]_net_1\, B => \CLKPHASE[4]_net_1\, 
        Y => N_215);
    
    \REG40M.BIT_OS_VAL_25_RNO[3]\ : MX2
      port map(A => \BIT_OS_VAL_25[3]\, B => N_209, S => 
        \un36_n_bit_os_val[6]\, Y => \N_BIT_OS_VAL_25_18[3]\);
    
    \CLKPHASE_RNIP0JI_0[0]\ : NOR3B
      port map(A => \CLKPHASE[0]_net_1\, B => N_5711, C => N_90, 
        Y => \un36_n_bit_os_val[18]\);
    
    \RECD_SER_WORD_RNO_2[7]\ : OR3
      port map(A => \ARB_BYTE_m_4[9]\, B => \ARB_BYTE_m_6[7]\, C
         => \N_RECD_SER_WORD_iv_3[7]\, Y => 
        \N_RECD_SER_WORD_iv_5[7]\);
    
    \WAITCNT[4]\ : DFN1E0C0
      port map(D => N_37, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_9, E => N_5790, Q => \WAITCNT[4]_net_1\);
    
    un41_n_seqcnts_I_12 : XOR2
      port map(A => N_2, B => \un39_n_seqcnts[4]\, Y => I_12);
    
    \REG40M.SEQCNTS_27_RNIJSNU[1]\ : MX2
      port map(A => \SEQCNTS_27[1]\, B => \SEQCNTS_28[1]\, S => 
        \INDEX_CNT[0]_net_1\, Y => N_4109);
    
    \REG40M.BIT_OS_CNT_1_RNO[6]\ : NOR3A
      port map(A => N_403, B => N_551, C => N_4530_1, Y => N_129);
    
    \INDEX_CNT_RNO[4]\ : NOR3B
      port map(A => N_5730, B => I_12_0, C => \DES_SM_1[8]_net_1\, 
        Y => \N_INDEX_CNT[4]\);
    
    \REG40M.BIT_OS_CNT_2_RNO[3]\ : XA1B
      port map(A => BIT_OS_CNT_2_c2, B => \BIT_OS_CNT_2[3]\, C
         => N_4530_0, Y => BIT_OS_CNT_2_n3);
    
    \REG40M.BIT_OS_VAL_6_RNI4FTE[3]\ : MX2
      port map(A => \BIT_OS_VAL_6[3]\, B => \BIT_OS_VAL_22[3]\, S
         => \CLKPHASE_2[4]_net_1\, Y => N_3702);
    
    \DES_SM_RNO[1]\ : NOR2A
      port map(A => \DES_SM[4]_net_1\, B => N_5730, Y => 
        \DES_SM_RNO[1]_net_1\);
    
    \CLKPHASE_1_RNIOG4D_0[2]\ : NOR3B
      port map(A => \CLKPHASE_0[1]_net_1\, B => N_212, C => 
        \CLKPHASE_1[2]_net_1\, Y => \un36_n_bit_os_val[13]\);
    
    \BEST_SEQCNT_RNO[1]\ : NOR2A
      port map(A => \un6_n_best_seqcnt[1]\, B => 
        \DES_SM_1[8]_net_1\, Y => \N_BEST_SEQCNT[1]\);
    
    \CLKPHASE_RNIOK8M2[2]\ : MX2
      port map(A => N_3811, B => N_3826, S => \CLKPHASE[2]_net_1\, 
        Y => N_3831);
    
    \WAITCNT_RNIJMUB1[6]\ : OR2A
      port map(A => \WAITCNT[6]_net_1\, B => N_5776, Y => N_5777);
    
    \REG40M.SEQCNTS_21_RNIVA4E[3]\ : MX2
      port map(A => \SEQCNTS_5[3]\, B => \SEQCNTS_21[3]\, S => 
        \CLKPHASE_1[4]_net_1\, Y => N_3776);
    
    \REG40M.BIT_OS_VAL_15_RNIFT2S[0]\ : MX2
      port map(A => \BIT_OS_VAL_31[0]\, B => \BIT_OS_VAL_15[0]\, 
        S => \CLKPHASE_3[4]_net_1\, Y => N_3599);
    
    \REG40M.BIT_OS_VAL_8[0]\ : DFN1E1C0
      port map(D => N_276, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_5, E => \DES_SM_1[6]_net_1\, Q => 
        \BIT_OS_VAL_8[0]\);
    
    \REG40M.BIT_OS_VAL_17_RNO[2]\ : MX2
      port map(A => \BIT_OS_VAL_17[2]\, B => N_781, S => 
        \un36_n_bit_os_val[14]\, Y => N_187);
    
    \REG40M.BIT_OS_CNT_3_RNO[2]\ : NOR2A
      port map(A => BIT_OS_CNT_3_n2_tz, B => N_4530, Y => 
        BIT_OS_CNT_3_n2);
    
    \MAX_CNT_RNILVO81[6]\ : NOR3A
      port map(A => DES_SM_tr5_0_a3_1, B => \MAX_CNT[6]_net_1\, C
         => \MAX_CNT[7]_net_1\, Y => DES_SM_tr5_0_a3_3);
    
    \DES_SM_RNICU2EH7_2[8]\ : AO1
      port map(A => \un36_n_bit_os_val[8]\, B => N_782, C => 
        N_717, Y => N_300);
    
    \CLKPHASE_RNIP0JI_0[1]\ : NOR3A
      port map(A => N_215, B => \CLKPHASE[1]_net_1\, C => N_5668, 
        Y => \un36_n_bit_os_val[6]\);
    
    \RECD_SER_WORD_RNO_3[0]\ : NOR3C
      port map(A => n_recd_ser_word167_1, B => 
        n_recd_ser_word171_0, C => \ARB_BYTE[7]_net_1\, Y => 
        \ARB_BYTE_m[7]\);
    
    \REG40M.BIT_OS_VAL_20[3]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_20_18[3]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_13, E => \DES_SM_2[6]_net_1\, Q
         => \BIT_OS_VAL_20[3]\);
    
    \Q[11]\ : DFN1C0
      port map(D => \ADJ_Q[11]_net_1\, CLK => CCC_160M_FXD, CLR
         => P_MASTER_POR_B_c_23, Q => \Q[11]_net_1\);
    
    \REG40M.BIT_OS_CNT_2_RNO[7]\ : XA1B
      port map(A => BIT_OS_CNT_2_c6, B => \BIT_OS_CNT_2[7]\, C
         => N_4530_0, Y => BIT_OS_CNT_2_n7);
    
    \DES_SM_0_RNIAB7UH7_1[8]\ : AO1A
      port map(A => N_5674, B => N_782_0, C => N_717_0, Y => 
        N_338);
    
    \REG40M.BIT_OS_VAL_8_RNI7O6I[3]\ : MX2
      port map(A => \BIT_OS_VAL_8[3]\, B => \BIT_OS_VAL_24[3]\, S
         => \CLKPHASE_1[4]_net_1\, Y => N_3666);
    
    \REG40M.BIT_OS_VAL_6_RNI2DTE[2]\ : MX2
      port map(A => \BIT_OS_VAL_6[2]\, B => \BIT_OS_VAL_22[2]\, S
         => \CLKPHASE_2[4]_net_1\, Y => N_3701);
    
    \DES_SM_RNI82M33[7]\ : AO1
      port map(A => BIT_OS_CNT_3lde_0_a3_3, B => N_562_3, C => 
        N_4530_1, Y => BIT_OS_CNT_3e);
    
    \REG40M.SEQCNTS_1_RNILO9K[2]\ : MX2
      port map(A => \SEQCNTS_1[2]\, B => \SEQCNTS_2[2]\, S => 
        \INDEX_CNT_1[0]_net_1\, Y => N_4000);
    
    \REG40M.SEQCNTS_25_RNI033Q[0]\ : MX2
      port map(A => \SEQCNTS_25[0]\, B => \SEQCNTS_26[0]\, S => 
        \INDEX_CNT_4[0]_net_1\, Y => N_4038);
    
    \INDEX_CNT_RNI390I7[4]\ : MX2
      port map(A => N_4032, B => N_4062, S => 
        \INDEX_CNT[4]_net_1\, Y => N_4067);
    
    \DES_SM_RNIBSRE[2]\ : OR2
      port map(A => \DES_SM[2]_net_1\, B => \DES_SM[3]_net_1\, Y
         => N_5783);
    
    \RECD_SER_WORD_RNO[6]\ : OR3
      port map(A => \N_RECD_SER_WORD_iv_1[6]\, B => 
        \N_RECD_SER_WORD_iv_0[6]\, C => \N_RECD_SER_WORD_iv_5[6]\, 
        Y => \N_RECD_SER_WORD[6]\);
    
    \INDEX_CNT_1_RNI8KNV1[3]\ : MX2
      port map(A => N_4000, B => N_4005, S => 
        \INDEX_CNT_1[3]_net_1\, Y => N_4010);
    
    \REG40M.SEQCNTS_9[4]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[4]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_20, E => N_328, Q => \SEQCNTS_9[4]\);
    
    \REG40M.SEQCNTS_20_RNIVQMJ[1]\ : MX2
      port map(A => \SEQCNTS_19[1]\, B => \SEQCNTS_20[1]\, S => 
        \INDEX_CNT_4[0]_net_1\, Y => N_4104);
    
    \REG40M.BIT_OS_VAL_15[0]\ : DFN1E1C0
      port map(D => N_258, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_15, E => \DES_SM_2[6]_net_1\, Q => 
        \BIT_OS_VAL_15[0]\);
    
    \REG40M.SEQCNTS_27_RNIH43Q[2]\ : MX2
      port map(A => \SEQCNTS_11[2]\, B => \SEQCNTS_27[2]\, S => 
        \CLKPHASE_2[4]_net_1\, Y => N_3745);
    
    \REG40M.BIT_OS_CNT_1_RNIKMOJ[6]\ : OR3B
      port map(A => \BIT_OS_CNT_1[5]\, B => \BIT_OS_CNT_1[6]\, C
         => N_381, Y => N_403);
    
    \REG40M.BIT_OS_VAL_7[2]\ : DFN1E1C0
      port map(D => N_205, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_3, E => \DES_SM_0[6]_net_1\, Q => 
        \BIT_OS_VAL_7[2]\);
    
    \CLKPHASE_RNIP60T9[0]\ : MX2
      port map(A => N_3794, B => N_3869, S => \CLKPHASE[0]_net_1\, 
        Y => \un39_n_seqcnts[1]\);
    
    \REG40M.BIT_OS_VAL_19[0]\ : DFN1E1C0
      port map(D => N_246, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_20, E => \DES_SM[6]_net_1\, Q => 
        \BIT_OS_VAL_19[0]\);
    
    \REG40M.BIT_OS_CNT_2_RNIENLF[3]\ : NOR2B
      port map(A => BIT_OS_CNT_2_c2, B => \BIT_OS_CNT_2[3]\, Y
         => BIT_OS_CNT_2_c3);
    
    \CLKPHASE_RNIP3SR9[0]\ : MX2
      port map(A => N_3793, B => N_3868, S => \CLKPHASE[0]_net_1\, 
        Y => \un39_n_seqcnts[0]\);
    
    \CLKPHASE_RNIP0JI[3]\ : NOR2B
      port map(A => N_211, B => N_5072_2, Y => 
        \un36_n_bit_os_val[1]\);
    
    \REG40M.BIT_OS_VAL_13[3]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_13_18[3]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_12, E => \DES_SM_2[6]_net_1\, Q
         => \BIT_OS_VAL_13[3]\);
    
    \INDEX_CNT_0_RNIU5HT1[3]\ : MX2
      port map(A => N_3998, B => N_4003, S => 
        \INDEX_CNT_0[3]_net_1\, Y => N_4008);
    
    \REG40M.BIT_OS_VAL_30_RNO[2]\ : MX2
      port map(A => \BIT_OS_VAL_30[2]\, B => N_781_0, S => 
        \un36_n_bit_os_val[1]\, Y => N_161);
    
    \REG40M.BIT_OS_CNT_3_RNO_0[2]\ : AX1C
      port map(A => \BIT_OS_CNT_3[1]\, B => \BIT_OS_CNT_3[0]\, C
         => \BIT_OS_CNT_3[2]\, Y => BIT_OS_CNT_3_n2_tz);
    
    \REG40M.BIT_OS_VAL_2[2]\ : DFN1E1C0
      port map(D => N_5653, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_18, E => \DES_SM_4[6]_net_1\, Q => 
        \BIT_OS_VAL_2[2]\);
    
    \WAITCNT_RNIFE3H1[9]\ : NOR3C
      port map(A => \WAITCNT[9]_net_1\, B => \WAITCNT[10]_net_1\, 
        C => un1_DES_SM_471_i_0_a2_0_0_a2_6, Y => 
        un1_DES_SM_471_i_0_a2_0_0_a2_9);
    
    \SYNC_SM.n_best_clkphase14_0_I_9\ : AO1C
      port map(A => \BEST_SEQCNT[3]_net_1\, B => 
        \un6_n_best_seqcnt[3]\, C => N_5, Y => N_10);
    
    \REG40M.BIT_OS_VAL_13_RNO[2]\ : MX2
      port map(A => \BIT_OS_VAL_13[2]\, B => N_781, S => 
        \un36_n_bit_os_val[18]\, Y => N_193);
    
    \REG40M.BIT_OS_CNT_5_RNIA3KL[2]\ : OR2A
      port map(A => \BIT_OS_CNT_5[2]\, B => N_367, Y => N_373);
    
    \BEST_BIT_OS_VAL[2]\ : DFN1E1C0
      port map(D => \N_BEST_BIT_OS_VAL[2]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_14, E => 
        un1_N_CCC_RESET_EN_0_sqmuxa, Q => 
        \BEST_BIT_OS_VAL[2]_net_1\);
    
    \REG40M.BIT_OS_VAL_7_RNO[3]\ : MX2
      port map(A => \BIT_OS_VAL_7[3]\, B => N_209, S => 
        \un36_n_bit_os_val[24]\, Y => \N_BIT_OS_VAL_7_18[3]\);
    
    \BEST_SEQCNT_RNO[0]\ : NOR2A
      port map(A => \un6_n_best_seqcnt[0]\, B => 
        \DES_SM_1[8]_net_1\, Y => \N_BEST_SEQCNT[0]\);
    
    \REG40M.SEQCNTS_29[1]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[1]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_16_0, E => N_288, Q => \SEQCNTS_29[1]\);
    
    \REG40M.SEQCNTS_28[0]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[0]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_15, E => N_290, Q => \SEQCNTS_28[0]\);
    
    \REG40M.BIT_OS_CNT_7_RNILJ0F1[4]\ : NOR2B
      port map(A => BIT_OS_CNT_7_c3, B => \BIT_OS_CNT_7[4]\, Y
         => BIT_OS_CNT_7_c4);
    
    \CLKPHASE_0_RNIVHOR[3]\ : MX2
      port map(A => N_3724, B => N_3729, S => 
        \CLKPHASE_0[3]_net_1\, Y => N_3734);
    
    \CLKPHASE_1_RNIQF2K2[2]\ : MX2
      port map(A => N_3809, B => N_3824, S => 
        \CLKPHASE_1[2]_net_1\, Y => N_3829);
    
    \REG40M.BIT_OS_VAL_27_RNO[2]\ : MX2
      port map(A => \BIT_OS_VAL_27[2]\, B => N_781_0, S => 
        \un36_n_bit_os_val[4]\, Y => N_167);
    
    \REG40M.BIT_OS_VAL_0_RNIUVDN[2]\ : MX2
      port map(A => \BIT_OS_VAL_0[2]\, B => \BIT_OS_VAL_16[2]\, S
         => \CLKPHASE_1[4]_net_1\, Y => N_3661);
    
    \REG40M.SEQCNTS_3_RNI0IVR[4]\ : MX2
      port map(A => \SEQCNTS_3[4]\, B => \SEQCNTS_4[4]\, S => 
        \INDEX_CNT_4[0]_net_1\, Y => N_4072);
    
    \REG40M.BIT_OS_VAL_15_RNIHV2S[1]\ : MX2
      port map(A => \BIT_OS_VAL_31[1]\, B => \BIT_OS_VAL_15[1]\, 
        S => \CLKPHASE_3[4]_net_1\, Y => N_3600);
    
    \REG40M.SEQCNTS_15[3]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[3]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_4, E => N_316, Q => \SEQCNTS_15[3]\);
    
    \RECD_SER_WORD_RNO_0[6]\ : AO1
      port map(A => \ARB_BYTE[12]_net_1\, B => n_recd_ser_word170, 
        C => \ARB_BYTE_m[13]\, Y => \N_RECD_SER_WORD_iv_1[6]\);
    
    \SYNC_SM.n_best_clkphase14_0_I_8\ : OR2A
      port map(A => \BEST_SEQCNT[4]_net_1\, B => 
        \un6_n_best_seqcnt[4]\, Y => N_9);
    
    \REG40M.BIT_OS_CNT_2_RNO[2]\ : XA1B
      port map(A => BIT_OS_CNT_2_c1, B => \BIT_OS_CNT_2[2]\, C
         => N_4530_0, Y => BIT_OS_CNT_2_n2);
    
    \DES_SM_0_RNIAB7UH7_4[8]\ : AO1
      port map(A => \un36_n_bit_os_val[20]\, B => N_782_0, C => 
        N_717_0, Y => N_324);
    
    \TUNE_CLKPHASE[3]\ : DFN1E1C0
      port map(D => \N_TUNE_CLKPHASE_2[3]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_13, E => \DES_SM[1]_net_1\, Q => 
        \TUNE_CLKPHASE[3]_net_1\);
    
    \REG40M.SEQCNTS_9[1]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[1]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_20, E => N_328, Q => \SEQCNTS_9[1]\);
    
    \REG40M.BIT_OS_VAL_22[3]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_22_18[3]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_15, E => \DES_SM_3[6]_net_1\, Q
         => \BIT_OS_VAL_22[3]\);
    
    \ARB_BYTE_RNI82M33[1]\ : AO1
      port map(A => BIT_OS_CNT_4lde_0_a3_1, B => N_561_3, C => 
        N_4530_0, Y => BIT_OS_CNT_4e);
    
    \REG40M.BIT_OS_VAL_30[2]\ : DFN1E1C0
      port map(D => N_161, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_18, E => \DES_SM_4[6]_net_1\, Q => 
        \BIT_OS_VAL_30[2]\);
    
    \REG40M.BIT_OS_CNT_5_RNO[1]\ : XA1B
      port map(A => \BIT_OS_CNT_5[0]\, B => \BIT_OS_CNT_5[1]\, C
         => N_4530, Y => N_5631);
    
    \REG40M.SEQCNTS_28_RNIG9CT[0]\ : MX2
      port map(A => \SEQCNTS_12[0]\, B => \SEQCNTS_28[0]\, S => 
        \CLKPHASE_3[4]_net_1\, Y => N_3818);
    
    un3_n_index_cnt_I_8 : AND3
      port map(A => \INDEX_CNT_0[0]_net_1\, B => 
        \INDEX_CNT[1]_net_1\, C => \INDEX_CNT_0[2]_net_1\, Y => 
        N_3);
    
    \REG40M.BIT_OS_VAL_2[1]\ : DFN1E1C0
      port map(D => N_5660, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_18, E => \DES_SM_4[6]_net_1\, Q => 
        \BIT_OS_VAL_2[1]\);
    
    \REG40M.BIT_OS_VAL_15[3]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_15_18[3]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_15, E => \DES_SM_2[6]_net_1\, Q
         => \BIT_OS_VAL_15[3]\);
    
    \REG40M.SEQCNTS_2[2]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[2]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_10, E => N_342, Q => \SEQCNTS_2[2]\);
    
    \DES_SM_RNIL4O0P[6]\ : NOR3C
      port map(A => \un107_bit_os_val[1]\, B => N_BIT_OS_VAL_3126, 
        C => N_761, Y => un1_DES_SM_1034_i_a2_3_2);
    
    \CLKPHASE_1_RNI17V81[3]\ : MX2
      port map(A => N_3761, B => N_3766, S => 
        \CLKPHASE_1[3]_net_1\, Y => N_3771);
    
    \INDEX_CNT_0_RNIH18A1[3]\ : MX2
      port map(A => N_4120, B => N_4125, S => 
        \INDEX_CNT_0[3]_net_1\, Y => N_4130);
    
    \REG40M.BIT_OS_CNT_1_RNO[1]\ : XA1B
      port map(A => \BIT_OS_CNT_1[0]\, B => \BIT_OS_CNT_1[1]\, C
         => N_4530_0, Y => N_139);
    
    \CLKPHASE_1_RNIT46B1[3]\ : MX2
      port map(A => N_3662, B => N_3666, S => 
        \CLKPHASE_1[3]_net_1\, Y => N_3670);
    
    \RECD_SER_WORD_RNIHHBK[4]\ : NOR2B
      port map(A => \RECD_SER_WORD[4]_net_1\, B => DCB_SALT_SEL_c, 
        Y => \ELK_RX_SER_WORD_0[4]\);
    
    \DES_SM_RNI74OM[7]\ : NOR3C
      port map(A => \ARB_BYTE[7]_net_1\, B => \DES_SM[7]_net_1\, 
        C => \ARB_BYTE[6]_net_1\, Y => N_563_2);
    
    \REG40M.BIT_OS_VAL_30_RNO[3]\ : MX2
      port map(A => \BIT_OS_VAL_30[3]\, B => N_209_0, S => 
        \un36_n_bit_os_val[1]\, Y => \N_BIT_OS_VAL_30_18[3]\);
    
    \MAX_CNT_RNIABA11[3]\ : NOR3C
      port map(A => \MAX_CNT[1]_net_1\, B => \MAX_CNT[3]_net_1\, 
        C => \MAX_CNT[0]_net_1\, Y => DES_SM_tr2_i_a3_4);
    
    \REG40M.SEQCNTS_23_RNI2KDH[3]\ : MX2
      port map(A => \SEQCNTS_7[3]\, B => \SEQCNTS_23[3]\, S => 
        \CLKPHASE_0[4]_net_1\, Y => N_3731);
    
    \BEST_BIT_OS_VAL_RNO_21[1]\ : MX2
      port map(A => \BIT_OS_VAL_21[1]\, B => \BIT_OS_VAL_22[1]\, 
        S => \INDEX_CNT[0]_net_1\, Y => N_3919);
    
    \REG40M.SEQCNTS_24_RNI640O[2]\ : MX2
      port map(A => \SEQCNTS_8[2]\, B => \SEQCNTS_24[2]\, S => 
        \CLKPHASE_4[4]_net_1\, Y => N_3805);
    
    \REG40M.SEQCNTS_19[4]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[4]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_11, E => N_308, Q => \SEQCNTS_19[4]\);
    
    \REG40M.BIT_OS_VAL_4_RNO[2]\ : MX2
      port map(A => N_781_0, B => \BIT_OS_VAL_4[2]\, S => N_5674, 
        Y => N_5651);
    
    \REG40M.BIT_OS_VAL_15_RNO[1]\ : MX2B
      port map(A => \BIT_OS_VAL_15[1]\, B => N_206, S => 
        \un36_n_bit_os_val[16]\, Y => \N_BIT_OS_VAL_15_18[1]\);
    
    \BEST_BIT_OS_VAL_RNO_0[0]\ : MX2
      port map(A => N_3930, B => N_3990, S => 
        \INDEX_CNT[1]_net_1\, Y => \N_BEST_BIT_OS_VAL_3[0]\);
    
    \CLKPHASE_0[1]\ : DFN1C0
      port map(D => \TUNE_CLKPHASE_RNI79F03[1]_net_1\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_24_0, Q => 
        \CLKPHASE_0[1]_net_1\);
    
    \SYNC_SM.n_best_clkphase14_0_I_7\ : AO1C
      port map(A => \BEST_SEQCNT[2]_net_1\, B => 
        \un6_n_best_seqcnt[2]\, C => N_2_1, Y => N_8);
    
    \CLKPHASE_RNIRT9H1[3]\ : MX2
      port map(A => N_3611, B => N_3615, S => \CLKPHASE[3]_net_1\, 
        Y => N_3619);
    
    \REG40M.BIT_OS_VAL_30_RNO[1]\ : MX2B
      port map(A => \BIT_OS_VAL_30[1]\, B => N_206, S => 
        \un36_n_bit_os_val[1]\, Y => \N_BIT_OS_VAL_30_18[1]\);
    
    \REG40M.SEQCNTS_17[2]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[2]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_7, E => N_312, Q => \SEQCNTS_17[2]\);
    
    \RECD_SER_WORD_RNIEEBK_0[1]\ : NOR2A
      port map(A => \RECD_SER_WORD[1]_net_1\, B => DCB_SALT_SEL_c, 
        Y => TFC_RX_SER_WORD(1));
    
    \REG40M.BIT_OS_CNT_7_RNIU37S[8]\ : OR3
      port map(A => \BIT_OS_CNT_7[4]\, B => \BIT_OS_CNT_7[8]\, C
         => \BIT_OS_CNT_7[5]\, Y => N_BIT_OS_VAL_3130lto8_2);
    
    \REG40M.SEQCNTS_22[4]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[4]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_5, E => N_302, Q => \SEQCNTS_22[4]\);
    
    \RECD_SER_WORD_RNO_1[0]\ : AO1
      port map(A => n_recd_ser_word168, B => \ARB_BYTE[4]_net_1\, 
        C => \ARB_BYTE_m[5]\, Y => \N_RECD_SER_WORD_iv_0[0]\);
    
    \BEST_BIT_OS_VAL_RNO_20[3]\ : MX2
      port map(A => \BIT_OS_VAL_25[3]\, B => \BIT_OS_VAL_26[3]\, 
        S => \INDEX_CNT_3[0]_net_1\, Y => N_3913);
    
    \ADJ_Q[5]\ : DFN1C0
      port map(D => \ADJ_Q[3]_net_1\, CLK => CCC_160M_ADJ, CLR
         => P_MASTER_POR_B_c_34_0, Q => \ADJ_Q[5]_net_1\);
    
    \REG40M.SEQCNTS_3[3]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[3]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_11, E => N_340, Q => \SEQCNTS_3[3]\);
    
    \REG40M.SEQCNTS_7[0]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[0]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_17_0, E => N_332, Q => \SEQCNTS_7[0]\);
    
    \REG40M.SEQCNTS_25[0]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[0]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_10, E => N_296, Q => \SEQCNTS_25[0]\);
    
    \REG40M.BIT_OS_VAL_24[2]\ : DFN1E1C0
      port map(D => N_173, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_18, E => \DES_SM_4[6]_net_1\, Q => 
        \BIT_OS_VAL_24[2]\);
    
    \MAX_CNT[6]\ : DFN1E0C0
      port map(D => N_5634, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_16, E => N_558, Q => \MAX_CNT[6]_net_1\);
    
    \CLKPHASE_RNITJCBB[0]\ : MX2
      port map(A => N_3656, B => N_3716, S => \CLKPHASE[0]_net_1\, 
        Y => \un107_bit_os_val[1]\);
    
    \RECD_SER_WORD_RNIFFBK_0[2]\ : NOR2A
      port map(A => \RECD_SER_WORD[2]_net_1\, B => DCB_SALT_SEL_c, 
        Y => TFC_RX_SER_WORD(2));
    
    \REG40M.BIT_OS_CNT_0[4]\ : DFN1E1C0
      port map(D => N_5640, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_3, E => BIT_OS_CNT_0e, Q => 
        \BIT_OS_CNT_0[4]\);
    
    \BIT_OS_SEL_1[2]\ : DFN1C0
      port map(D => \BEST_BIT_OS_VAL[2]_net_1\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_27_1, Q => 
        \BIT_OS_SEL_1[2]_net_1\);
    
    \REG40M.BIT_OS_VAL_23_RNO[2]\ : MX2
      port map(A => \BIT_OS_VAL_23[2]\, B => N_781, S => 
        \un36_n_bit_os_val[8]\, Y => N_5641);
    
    \CLKPHASE_RNITIBBB[0]\ : MX2
      port map(A => N_3655, B => N_3715, S => \CLKPHASE[0]_net_1\, 
        Y => \un107_bit_os_val[0]\);
    
    \CLKPHASE_2_RNIC41I1[3]\ : MX2
      port map(A => N_3600, B => N_3604, S => 
        \CLKPHASE_2[3]_net_1\, Y => N_3608);
    
    \REG40M.BIT_OS_CNT_0_RNO[8]\ : XA1C
      port map(A => \BIT_OS_CNT_0[8]\, B => N_435, C => N_4530_2, 
        Y => N_107);
    
    \REG40M.SEQCNTS_23_RNISEAH[2]\ : MX2
      port map(A => \SEQCNTS_23[2]\, B => \SEQCNTS_24[2]\, S => 
        \INDEX_CNT_0[0]_net_1\, Y => N_4120);
    
    \DES_SM_RNIJSGE4[0]\ : AO1
      port map(A => N_5859, B => \DES_SM[0]_net_1\, C => N_140, Y
         => \DES_SM_ns[0]\);
    
    \CLKPHASE_RNIP0JI_7[0]\ : NOR2B
      port map(A => N_214, B => N_204, Y => 
        \un36_n_bit_os_val[8]\);
    
    \RECD_SER_WORD_RNIDDBK[0]\ : NOR2B
      port map(A => \RECD_SER_WORD[0]_net_1\, B => DCB_SALT_SEL_c, 
        Y => \ELK_RX_SER_WORD_0[0]\);
    
    \REG40M.BIT_OS_VAL_17_RNO[3]\ : MX2
      port map(A => \BIT_OS_VAL_17[3]\, B => N_209, S => 
        \un36_n_bit_os_val[14]\, Y => \N_BIT_OS_VAL_17_18[3]\);
    
    \REG40M.SEQCNTS_6[0]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[0]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_16, E => N_334, Q => \SEQCNTS_6[0]\);
    
    \REG40M.SEQCNTS_18_RNI5SJH[3]\ : MX2
      port map(A => \SEQCNTS_2[3]\, B => \SEQCNTS_18[3]\, S => 
        \CLKPHASE_4[4]_net_1\, Y => N_3836);
    
    \BEST_BIT_OS_VAL_RNO_25[0]\ : MX2
      port map(A => \BIT_OS_VAL_15[0]\, B => \BIT_OS_VAL_16[0]\, 
        S => \INDEX_CNT_2[0]_net_1\, Y => N_3950);
    
    \REG40M.BIT_OS_VAL_11_RNO[2]\ : MX2
      port map(A => \BIT_OS_VAL_11[2]\, B => N_781_0, S => 
        \un36_n_bit_os_val[20]\, Y => N_197);
    
    \SYNC_SM.N_TUNE_CLKPHASE_2_0_0_ADD_5x5_slow_I0_un1_S\ : XOR2
      port map(A => \BEST_CLKPHASE[0]_net_1\, B => 
        \BEST_SEQCNT[1]_net_1\, Y => I0_un1_S);
    
    \MAX_CNT_RNO[4]\ : XA1C
      port map(A => \MAX_CNT[4]_net_1\, B => N_375, C => 
        un1_DES_SM_19, Y => N_5636);
    
    \ADJ_Q[12]\ : DFN1C0
      port map(D => \ADJ_Q[10]_net_1\, CLK => CCC_160M_ADJ, CLR
         => P_MASTER_POR_B_c_26, Q => \ADJ_Q[12]_net_1\);
    
    \REG40M.SEQCNTS_7_RNIHH051[2]\ : MX2
      port map(A => \SEQCNTS_7[2]\, B => \SEQCNTS_8[2]\, S => 
        \INDEX_CNT[0]_net_1\, Y => N_4085);
    
    \REG40M.SEQCNTS_17_RNISCAE[0]\ : MX2
      port map(A => \SEQCNTS_1[0]\, B => \SEQCNTS_17[0]\, S => 
        \CLKPHASE_3[4]_net_1\, Y => N_3758);
    
    \REG40M.BIT_OS_CNT_1_RNO_0[6]\ : OA1C
      port map(A => \BIT_OS_CNT_1[5]\, B => N_381, C => 
        \BIT_OS_CNT_1[6]\, Y => N_551);
    
    \REG40M.BIT_OS_VAL_15_RNIJ13S[2]\ : MX2
      port map(A => \BIT_OS_VAL_31[2]\, B => \BIT_OS_VAL_15[2]\, 
        S => \CLKPHASE_3[4]_net_1\, Y => N_3601);
    
    \REG40M.BIT_OS_CNT_1[3]\ : DFN1E1C0
      port map(D => N_135, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_4, E => BIT_OS_CNT_1e, Q => 
        \BIT_OS_CNT_1[3]\);
    
    \REG40M.SEQCNTS_24[2]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[2]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_8, E => N_298, Q => \SEQCNTS_24[2]\);
    
    \REG40M.BIT_OS_VAL_4[3]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_4_18[3]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_21, E => \DES_SM[6]_net_1\, Q => 
        \BIT_OS_VAL_4[3]\);
    
    \REG40M.BIT_OS_CNT_6_RNIS8GMA_0[7]\ : AO1A
      port map(A => N_BIT_OS_VAL_3126, B => N_84, C => 
        N_BIT_OS_VAL_3130, Y => N_5666_0);
    
    \REG40M.BIT_OS_VAL_3[0]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_3_18[0]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_19, E => \DES_SM_4[6]_net_1\, Q
         => \BIT_OS_VAL_3[0]\);
    
    \DES_SM_RNICU2EH7_4[8]\ : AO1
      port map(A => \un36_n_bit_os_val[1]\, B => N_782, C => 
        N_717, Y => N_286);
    
    \REG40M.BIT_OS_CNT_4_RNO_0[3]\ : NOR2A
      port map(A => N_429, B => \BIT_OS_CNT_4[3]\, Y => N_504);
    
    \REG40M.SEQCNTS_12[0]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[0]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_21, E => N_322, Q => \SEQCNTS_12[0]\);
    
    \REG40M.BIT_OS_VAL_7_RNO[0]\ : MX2
      port map(A => \BIT_OS_VAL_7[0]\, B => N_5666, S => 
        \un36_n_bit_os_val[24]\, Y => N_279);
    
    \Q[13]\ : DFN1C0
      port map(D => \ADJ_Q[13]_net_1\, CLK => CCC_160M_FXD, CLR
         => P_MASTER_POR_B_c_23, Q => \Q[13]_net_1\);
    
    \REG40M.BIT_OS_VAL_25_RNO[1]\ : MX2B
      port map(A => \BIT_OS_VAL_25[1]\, B => N_206_0, S => 
        \un36_n_bit_os_val[6]\, Y => \N_BIT_OS_VAL_25_18[1]\);
    
    \REG40M.SEQCNTS_8[3]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[3]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_19, E => N_330, Q => \SEQCNTS_8[3]\);
    
    \INDEX_CNT_3[0]\ : DFN1E0C0
      port map(D => \N_INDEX_CNT[0]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_16_0, E => N_5149, Q => 
        \INDEX_CNT_3[0]_net_1\);
    
    \REG40M.BIT_OS_CNT_7_RNO[0]\ : NOR2
      port map(A => \BIT_OS_CNT_7[0]\, B => N_4530, Y => N_5615);
    
    \INDEX_CNT_RNIJI083[2]\ : MX2
      port map(A => N_4046, B => N_4056, S => 
        \INDEX_CNT[2]_net_1\, Y => N_4061);
    
    \CLKPHASE_0_RNIRG0G2[2]\ : MX2
      port map(A => N_3844, B => N_3859, S => 
        \CLKPHASE_0[2]_net_1\, Y => N_3864);
    
    \REG40M.BIT_OS_VAL_5[2]\ : DFN1E1C0
      port map(D => N_207, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_1, E => \DES_SM_0[6]_net_1\, Q => 
        \BIT_OS_VAL_5[2]\);
    
    \INDEX_CNT_RNIQP083[2]\ : MX2
      port map(A => N_4047, B => N_4057, S => 
        \INDEX_CNT[2]_net_1\, Y => N_4062);
    
    \REG40M.BIT_OS_VAL_31[1]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_31_18[1]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_20, E => \DES_SM_4[6]_net_1\, Q
         => \BIT_OS_VAL_31[1]\);
    
    \REG40M.SEQCNTS_30_RNIVHVA[3]\ : MX2
      port map(A => \SEQCNTS_14[3]\, B => \SEQCNTS_30[3]\, S => 
        \CLKPHASE[4]_net_1\, Y => N_3856);
    
    \DES_SM_0_RNIKRD5U[8]\ : NOR2A
      port map(A => I_7, B => \DES_SM_0[8]_net_1\, Y => 
        \N_SEQCNTS_1_0[2]\);
    
    \REG40M.BIT_OS_VAL_25[0]\ : DFN1E1C0
      port map(D => N_228, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_20, E => \DES_SM[6]_net_1\, Q => 
        \BIT_OS_VAL_25[0]\);
    
    \REG40M.SEQCNTS_29[0]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[0]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_16_0, E => N_288, Q => \SEQCNTS_29[0]\);
    
    \REG40M.SEQCNTS_28[4]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[4]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_15, E => N_290, Q => \SEQCNTS_28[4]\);
    
    \REG40M.BIT_OS_VAL_29[0]\ : DFN1E1C0
      port map(D => N_216, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_4, E => \DES_SM_1[6]_net_1\, Q => 
        \BIT_OS_VAL_29[0]\);
    
    \WAITCNT_RNIV9DL_0[8]\ : NOR2
      port map(A => \WAITCNT[12]_net_1\, B => \WAITCNT[8]_net_1\, 
        Y => \DES_SM_ns_0_0_0_a2_0[0]\);
    
    \REG40M.SEQCNTS_28[1]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[1]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_15, E => N_290, Q => \SEQCNTS_28[1]\);
    
    \REG40M.BIT_OS_VAL_2[0]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_2_18[0]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_18, E => \DES_SM_4[6]_net_1\, Q
         => \BIT_OS_VAL_2[0]\);
    
    \REG40M.BIT_OS_VAL_23[3]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_23_18[3]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_17_0, E => \DES_SM_3[6]_net_1\, Q
         => \BIT_OS_VAL_23[3]\);
    
    \REG40M.BIT_OS_CNT_3_RNIIV1F[8]\ : OR3
      port map(A => \BIT_OS_CNT_3[4]\, B => \BIT_OS_CNT_3[8]\, C
         => \BIT_OS_CNT_3[5]\, Y => N_BIT_OS_VAL_3114lto8_2);
    
    \REG40M.BIT_OS_CNT_0_RNO[1]\ : XA1B
      port map(A => \BIT_OS_CNT_0[0]\, B => \BIT_OS_CNT_0[1]\, C
         => N_4530_2, Y => N_121);
    
    \CLKPHASE_1_RNIKJMG2[2]\ : MX2
      port map(A => N_3669, B => N_3681, S => 
        \CLKPHASE_1[2]_net_1\, Y => N_3685);
    
    \REG40M.SEQCNTS_9[2]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[2]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_20, E => N_328, Q => \SEQCNTS_9[2]\);
    
    \BEST_BIT_OS_VAL_RNO_22[2]\ : MX2
      port map(A => \BIT_OS_VAL_3[2]\, B => \BIT_OS_VAL_4[2]\, S
         => \INDEX_CNT_0[0]_net_1\, Y => N_3936);
    
    \REG40M.SEQCNTS_11[2]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[2]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_20, E => N_324, Q => \SEQCNTS_11[2]\);
    
    \INDEX_CNT_1_RNICONV1[3]\ : MX2
      port map(A => N_4001, B => N_4006, S => 
        \INDEX_CNT_1[3]_net_1\, Y => N_4011);
    
    \DES_SM_1_RNI14SU1[8]\ : NOR3A
      port map(A => N_5730, B => \DES_SM_1[8]_net_1\, C => 
        \INDEX_CNT_4[0]_net_1\, Y => \N_INDEX_CNT[0]\);
    
    \REG40M.SEQCNTS_26[2]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[2]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_12, E => N_294, Q => \SEQCNTS_26[2]\);
    
    \REG40M.BIT_OS_VAL_27_RNO[3]\ : MX2
      port map(A => \BIT_OS_VAL_27[3]\, B => N_209_0, S => 
        \un36_n_bit_os_val[4]\, Y => \N_BIT_OS_VAL_27_18[3]\);
    
    \INDEX_CNT_2_RNIBDCJ1[3]\ : MX2
      port map(A => N_4017, B => N_4022, S => 
        \INDEX_CNT_2[3]_net_1\, Y => N_4027);
    
    \RECD_SER_WORD_RNO[4]\ : OR3
      port map(A => \N_RECD_SER_WORD_iv_1[4]\, B => 
        \N_RECD_SER_WORD_iv_0[4]\, C => \N_RECD_SER_WORD_iv_5[4]\, 
        Y => \N_RECD_SER_WORD[4]\);
    
    \WAITCNT[12]\ : DFN1E0C0
      port map(D => WAITCNT_n12, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_21, E => N_5790, Q => 
        \WAITCNT[12]_net_1\);
    
    \REG40M.BIT_OS_VAL_21_RNO[2]\ : MX2
      port map(A => \BIT_OS_VAL_21[2]\, B => N_781, S => 
        \un36_n_bit_os_val[10]\, Y => N_179);
    
    \RECD_SER_WORD_RNO_7[7]\ : AO1
      port map(A => \ARB_BYTE[8]_net_1\, B => n_recd_ser_word165, 
        C => \ARB_BYTE_m_3[10]\, Y => \N_RECD_SER_WORD_iv_3[7]\);
    
    \MAX_CNT[5]\ : DFN1E0C0
      port map(D => N_5635, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_16, E => N_558, Q => \MAX_CNT[5]_net_1\);
    
    \INDEX_CNT_RNIAF3N4[2]\ : MX2
      port map(A => N_4082, B => N_4097, S => 
        \INDEX_CNT[2]_net_1\, Y => N_4102);
    
    \INDEX_CNT_RNI9JHU3[2]\ : MX2
      port map(A => N_4011, B => N_4026, S => 
        \INDEX_CNT[2]_net_1\, Y => N_4031);
    
    \REG40M.BIT_OS_CNT_4_RNI7QAI[2]\ : OR3C
      port map(A => \BIT_OS_CNT_4[1]\, B => \BIT_OS_CNT_4[2]\, C
         => \BIT_OS_CNT_4[0]\, Y => N_429);
    
    \MAX_CNT_RNO[7]\ : XA1C
      port map(A => \MAX_CNT[7]_net_1\, B => N_405, C => 
        un1_DES_SM_19, Y => N_5633);
    
    \REG40M.BIT_OS_VAL_10_RNIHQPM[2]\ : MX2
      port map(A => \BIT_OS_VAL_10[2]\, B => \BIT_OS_VAL_26[2]\, 
        S => \CLKPHASE_2[4]_net_1\, Y => N_3693);
    
    \REG40M.BIT_OS_CNT_6_RNO[1]\ : XA1B
      port map(A => \BIT_OS_CNT_6[0]\, B => \BIT_OS_CNT_6[1]\, C
         => N_4530_1, Y => N_85);
    
    \DES_SM_0[6]\ : DFN1C0
      port map(D => N_MAX_CNT_0_sqmuxa, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_27_1, Q => \DES_SM_0[6]_net_1\);
    
    \REG40M.BIT_OS_VAL_9_RNO[3]\ : MX2
      port map(A => \BIT_OS_VAL_9[3]\, B => N_209_0, S => 
        \un36_n_bit_os_val[22]\, Y => \N_BIT_OS_VAL_9_18[3]\);
    
    \REG40M.BIT_OS_CNT_4_RNO[0]\ : NOR2
      port map(A => \BIT_OS_CNT_4[0]\, B => N_4530, Y => N_507);
    
    \CLKPHASE_2_RNIKC1I1[3]\ : MX2
      port map(A => N_3602, B => N_3606, S => 
        \CLKPHASE_2[3]_net_1\, Y => N_3610);
    
    \REG40M.BIT_OS_VAL_25[3]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_25_18[3]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_20, E => \DES_SM[6]_net_1\, Q => 
        \BIT_OS_VAL_25[3]\);
    
    \REG40M.SEQCNTS_30[3]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[3]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_8, E => N_286, Q => \SEQCNTS_30[3]\);
    
    \REG40M.BIT_OS_VAL_10[1]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_10_18[1]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_6, E => \DES_SM_1[6]_net_1\, Q
         => \BIT_OS_VAL_10[1]\);
    
    \RECD_SER_WORD_RNO_0[3]\ : AO1
      port map(A => \ARB_BYTE[9]_net_1\, B => n_recd_ser_word170, 
        C => \ARB_BYTE_m[10]\, Y => \N_RECD_SER_WORD_iv_1[3]\);
    
    \DES_SM_RNILO5VH1[8]\ : NOR2A
      port map(A => I_12, B => \DES_SM[8]_net_1\, Y => 
        \N_SEQCNTS_1[4]\);
    
    \CLKPHASE_RNIP0JI_0[3]\ : NOR2A
      port map(A => N_211, B => N_90, Y => \un36_n_bit_os_val[3]\);
    
    \REG40M.SEQCNTS_13[3]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[3]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_1, E => N_320, Q => \SEQCNTS_13[3]\);
    
    \REG40M.SEQCNTS_5_RNIUJ5U[2]\ : MX2
      port map(A => \SEQCNTS_5[2]\, B => \SEQCNTS_6[2]\, S => 
        \INDEX_CNT_2[0]_net_1\, Y => N_4015);
    
    \CLKPHASE_RNI8FQ75[1]\ : MX2
      port map(A => N_3830, B => N_3865, S => \CLKPHASE[1]_net_1\, 
        Y => N_3870);
    
    \ARB_BYTE_RNIEV161_0[2]\ : NOR3B
      port map(A => \ARB_BYTE[2]_net_1\, B => N_562_3, C => 
        \ARB_BYTE[5]_net_1\, Y => BIT_OS_CNT_7lde_0_a3_1);
    
    \CLKPHASE_RNITSGNF1[0]\ : NOR3B
      port map(A => \un107_bit_os_val[2]\, B => 
        un1_DES_SM_1034_i_a2_3_2, C => \un107_bit_os_val[0]\, Y
         => N_758);
    
    \CLKPHASE_0_RNIUCJI4[1]\ : MX2
      port map(A => N_3756, B => N_3791, S => 
        \CLKPHASE_0[1]_net_1\, Y => N_3796);
    
    \REG40M.SEQCNTS_22_RNI1PMK[1]\ : MX2
      port map(A => \SEQCNTS_6[1]\, B => \SEQCNTS_22[1]\, S => 
        \CLKPHASE_5[4]_net_1\, Y => N_3849);
    
    \DES_SM_RNICU2EH7_3[8]\ : AO1
      port map(A => \un36_n_bit_os_val[0]\, B => N_782, C => 
        N_717, Y => N_284);
    
    \DES_SM_1[6]\ : DFN1C0
      port map(D => N_MAX_CNT_0_sqmuxa, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_27_1, Q => \DES_SM_1[6]_net_1\);
    
    \WAITCNT_RNO[12]\ : XA1C
      port map(A => \WAITCNT[12]_net_1\, B => N_5785, C => N_4539, 
        Y => WAITCNT_n12);
    
    \CLKPHASE_1_RNIPTE92[2]\ : MX2
      port map(A => N_3734, B => N_3749, S => 
        \CLKPHASE_1[2]_net_1\, Y => N_3754);
    
    \TUNE_CLKPHASE[4]\ : DFN1E1C0
      port map(D => N_1, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_13, E => \DES_SM[1]_net_1\, Q => 
        \TUNE_CLKPHASE[4]_net_1\);
    
    \REG40M.SEQCNTS_25_RNI473Q[2]\ : MX2
      port map(A => \SEQCNTS_25[2]\, B => \SEQCNTS_26[2]\, S => 
        \INDEX_CNT_4[0]_net_1\, Y => N_4040);
    
    \REG40M.SEQCNTS_21_RNIR64E[1]\ : MX2
      port map(A => \SEQCNTS_5[1]\, B => \SEQCNTS_21[1]\, S => 
        \CLKPHASE_1[4]_net_1\, Y => N_3774);
    
    \REG40M.SEQCNTS_19_RNI4PGG[3]\ : MX2
      port map(A => \SEQCNTS_3[3]\, B => \SEQCNTS_19[3]\, S => 
        \CLKPHASE_1[4]_net_1\, Y => N_3741);
    
    \REG40M.BIT_OS_VAL_2_RNI0AQR[1]\ : MX2
      port map(A => \BIT_OS_VAL_2[1]\, B => \BIT_OS_VAL_18[1]\, S
         => \CLKPHASE_1[4]_net_1\, Y => N_3688);
    
    \REG40M.BIT_OS_VAL_5_RNI1E0G[1]\ : MX2
      port map(A => \BIT_OS_VAL_5[1]\, B => \BIT_OS_VAL_21[1]\, S
         => \CLKPHASE_5[4]_net_1\, Y => N_3640);
    
    \BEST_SEQCNT_RNO[2]\ : NOR2A
      port map(A => \un6_n_best_seqcnt[2]\, B => 
        \DES_SM_1[8]_net_1\, Y => \N_BEST_SEQCNT[2]\);
    
    \INDEX_CNT_0_RNIK48A1[3]\ : MX2
      port map(A => N_4121, B => N_4126, S => 
        \INDEX_CNT_0[3]_net_1\, Y => N_4131);
    
    \DES_SM_RNICT161[7]\ : NOR2B
      port map(A => N_776, B => N_563_2, Y => 
        BIT_OS_CNT_5lde_0_a3_2);
    
    \REG40M.BIT_OS_CNT_1[8]\ : DFN1E1C0
      port map(D => N_125, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_4, E => BIT_OS_CNT_1e, Q => 
        \BIT_OS_CNT_1[8]\);
    
    \BEST_BIT_OS_VAL_RNO_28[0]\ : MX2
      port map(A => \BIT_OS_VAL_23[0]\, B => \BIT_OS_VAL_24[0]\, 
        S => \INDEX_CNT_2[0]_net_1\, Y => N_3974);
    
    \CLKPHASE_2_RNIAABG1[3]\ : MX2
      port map(A => N_3815, B => N_3820, S => 
        \CLKPHASE_2[3]_net_1\, Y => N_3825);
    
    \ADJ_Q[11]\ : DFN1C0
      port map(D => \ADJ_Q[9]_net_1\, CLK => CCC_160M_ADJ, CLR
         => P_MASTER_POR_B_c_26, Q => \ADJ_Q[11]_net_1\);
    
    \REG40M.SEQCNTS_4[2]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[2]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_13, E => N_338, Q => \SEQCNTS_4[2]\);
    
    \INDEX_CNT_0[2]\ : DFN1E0C0
      port map(D => \N_INDEX_CNT[2]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_17_0, E => N_5149, Q => 
        \INDEX_CNT_0[2]_net_1\);
    
    un41_n_seqcnts_I_7 : XOR2
      port map(A => N_4, B => \un39_n_seqcnts[2]\, Y => I_7);
    
    \REG40M.SEQCNTS_25_RNICE6Q[4]\ : MX2
      port map(A => \SEQCNTS_9[4]\, B => \SEQCNTS_25[4]\, S => 
        \CLKPHASE_4[4]_net_1\, Y => N_3767);
    
    \WAITCNT_RNO[9]\ : XA1C
      port map(A => \WAITCNT[9]_net_1\, B => N_5779, C => N_4539, 
        Y => N_5810);
    
    \REG40M.BIT_OS_CNT_6_RNO[3]\ : NOR3A
      port map(A => N_378, B => N_524, C => N_4530_1, Y => N_81);
    
    \REG40M.BIT_OS_CNT_4[1]\ : DFN1E1C0
      port map(D => N_5624, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_9, E => BIT_OS_CNT_4e, Q => 
        \BIT_OS_CNT_4[1]\);
    
    \ARB_BYTE_RNICT161[1]\ : NOR3C
      port map(A => \ARB_BYTE[4]_net_1\, B => \ARB_BYTE[1]_net_1\, 
        C => N_560_2, Y => BIT_OS_CNT_2lde_0_a3_1);
    
    \REG40M.BIT_OS_CNT_5_RNO[2]\ : XA1C
      port map(A => \BIT_OS_CNT_5[2]\, B => N_367, C => N_4530, Y
         => N_5630);
    
    \REG40M.BIT_OS_CNT_0[3]\ : DFN1E1C0
      port map(D => N_117, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_3, E => BIT_OS_CNT_0e, Q => 
        \BIT_OS_CNT_0[3]\);
    
    \DES_SM_0_RNIAB7UH7_3[8]\ : AO1
      port map(A => \un36_n_bit_os_val[16]\, B => N_782_0, C => 
        N_717_0, Y => N_316);
    
    \BEST_BIT_OS_VAL_RNO_25[3]\ : MX2
      port map(A => \BIT_OS_VAL_15[3]\, B => \BIT_OS_VAL_16[3]\, 
        S => \INDEX_CNT_2[0]_net_1\, Y => N_3953);
    
    \BEST_BIT_OS_VAL_RNO_14[3]\ : MX2
      port map(A => N_3977, B => N_3981, S => 
        \INDEX_CNT_2[3]_net_1\, Y => N_3985);
    
    \REG40M.SEQCNTS_11[4]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[4]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_20, E => N_324, Q => \SEQCNTS_11[4]\);
    
    un1_CLKPHASE_I_24 : NOR2B
      port map(A => \DWACT_ADD_CI_0_g_array_1[0]\, B => 
        \CLKPHASE[2]_net_1\, Y => \DWACT_ADD_CI_0_g_array_12[0]\);
    
    \CLKPHASE_RNIP0JI_2[3]\ : NOR2
      port map(A => N_5672, B => N_90, Y => 
        \un36_n_bit_os_val[19]\);
    
    \BEST_BIT_OS_VAL_RNO_19[1]\ : MX2
      port map(A => \BIT_OS_VAL_17[1]\, B => \BIT_OS_VAL_18[1]\, 
        S => \INDEX_CNT_3[0]_net_1\, Y => N_3907);
    
    \CLKPHASE_0_RNIID1G2[2]\ : MX2
      port map(A => N_3635, B => N_3647, S => 
        \CLKPHASE_0[2]_net_1\, Y => N_3651);
    
    \REG40M.BIT_OS_VAL_16[2]\ : DFN1E1C0
      port map(D => N_189, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_16_0, E => \DES_SM_3[6]_net_1\, Q => 
        \BIT_OS_VAL_16[2]\);
    
    \DES_SM_RNI1S8UM[6]\ : NOR2A
      port map(A => N_761, B => \un107_bit_os_val[1]\, Y => N_762);
    
    \SYNC_SM.n_best_clkphase14_0_I_3\ : NOR2A
      port map(A => \un6_n_best_seqcnt[0]\, B => 
        \BEST_SEQCNT[0]_net_1\, Y => N_4_1);
    
    \WAITCNT_RNIQFQA1[5]\ : NOR3C
      port map(A => \WAITCNT[11]_net_1\, B => \WAITCNT[5]_net_1\, 
        C => un1_DES_SM_471_i_0_a2_0_0_a2_4, Y => 
        un1_DES_SM_471_i_0_a2_0_0_a2_8);
    
    \REG40M.BIT_OS_CNT_0[0]\ : DFN1E1C0
      port map(D => N_547, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_2, E => BIT_OS_CNT_0e, Q => 
        \BIT_OS_CNT_0[0]\);
    
    \REG40M.SEQCNTS_13_RNINIFE[3]\ : MX2
      port map(A => \SEQCNTS_13[3]\, B => \SEQCNTS_29[3]\, S => 
        \CLKPHASE_2[4]_net_1\, Y => N_3781);
    
    \REG40M.BIT_OS_CNT_7[7]\ : DFN1E1C0
      port map(D => BIT_OS_CNT_7_n7, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_14, E => BIT_OS_CNT_7e, Q => 
        \BIT_OS_CNT_7[7]\);
    
    \REG40M.SEQCNTS_21[0]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[0]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_3, E => N_304, Q => \SEQCNTS_21[0]\);
    
    \REG40M.BIT_OS_CNT_5_RNO_0[8]\ : OR2A
      port map(A => \BIT_OS_CNT_5[7]\, B => N_409, Y => N_421);
    
    \REG40M.SEQCNTS_17_RNI8D3M[3]\ : MX2
      port map(A => \SEQCNTS_17[3]\, B => \SEQCNTS_18[3]\, S => 
        \INDEX_CNT_4[0]_net_1\, Y => N_4036);
    
    \REG40M.BIT_OS_CNT_3_RNO[6]\ : XA1B
      port map(A => BIT_OS_CNT_3_c5, B => \BIT_OS_CNT_3[6]\, C
         => N_4530_1, Y => BIT_OS_CNT_3_n6);
    
    \REG40M.BIT_OS_CNT_3[2]\ : DFN1E1C0
      port map(D => BIT_OS_CNT_3_n2, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_7, E => BIT_OS_CNT_3e, Q => 
        \BIT_OS_CNT_3[2]\);
    
    \ARB_BYTE_RNI3N9F[0]\ : NOR2A
      port map(A => \ARB_BYTE[0]_net_1\, B => \ARB_BYTE[3]_net_1\, 
        Y => N_772);
    
    un1_DES_SM_1003_i_0_a3 : NOR2A
      port map(A => \DES_SM[8]_net_1\, B => \DES_SM[4]_net_1\, Y
         => N_5792);
    
    \REG40M.BIT_OS_CNT_3_RNO[8]\ : XA1B
      port map(A => BIT_OS_CNT_3_432_0, B => \BIT_OS_CNT_3[8]\, C
         => N_4530_1, Y => BIT_OS_CNT_3_n8);
    
    \CLKPHASE_2[4]\ : DFN1C0
      port map(D => \TUNE_CLKPHASE_RNITINS2[4]_net_1\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_24_0, Q => 
        \CLKPHASE_2[4]_net_1\);
    
    \BEST_BIT_OS_VAL_RNO_7[0]\ : MX2
      port map(A => N_3878, B => N_3882, S => 
        \INDEX_CNT_0[3]_net_1\, Y => N_3886);
    
    \CLKPHASE_2_RNI66BG1[3]\ : MX2
      port map(A => N_3814, B => N_3819, S => 
        \CLKPHASE_2[3]_net_1\, Y => N_3824);
    
    \CLKPHASE_1_RNI1V7F1[3]\ : MX2
      port map(A => N_3813, B => N_3818, S => 
        \CLKPHASE_1[3]_net_1\, Y => N_3823);
    
    \CLKPHASE_2_RNI23621[3]\ : MX2
      port map(A => N_3800, B => N_3805, S => 
        \CLKPHASE_2[3]_net_1\, Y => N_3810);
    
    \INDEX_CNT_1_RNIPM5H1[3]\ : MX2
      port map(A => N_4013, B => N_4018, S => 
        \INDEX_CNT_1[3]_net_1\, Y => N_4023);
    
    \DES_SM_RNIDLMT71[8]\ : NOR2A
      port map(A => I_9, B => \DES_SM[8]_net_1\, Y => 
        \N_SEQCNTS_1[3]\);
    
    un3_n_index_cnt_I_6 : NOR2B
      port map(A => \INDEX_CNT[1]_net_1\, B => 
        \INDEX_CNT[0]_net_1\, Y => N_4_0);
    
    \REG40M.SEQCNTS_10[2]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[2]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_18, E => N_326, Q => \SEQCNTS_10[2]\);
    
    \REG40M.BIT_OS_CNT_3_RNO[4]\ : NOR2A
      port map(A => BIT_OS_CNT_3_n4_tz, B => N_4530, Y => 
        BIT_OS_CNT_3_n4);
    
    \REG40M.BIT_OS_VAL_6_RNIU8TE[0]\ : MX2
      port map(A => \BIT_OS_VAL_6[0]\, B => \BIT_OS_VAL_22[0]\, S
         => \CLKPHASE_2[4]_net_1\, Y => N_3699);
    
    \REG40M.BIT_OS_VAL_15[1]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_15_18[1]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_15, E => \DES_SM_2[6]_net_1\, Q
         => \BIT_OS_VAL_15[1]\);
    
    \REG40M.SEQCNTS_3[4]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[4]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_11, E => N_340, Q => \SEQCNTS_3[4]\);
    
    \ARB_WRD_40M_FIXED[9]\ : DFN1C0
      port map(D => \Q[9]_net_1\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_26, Q => \ARB_WRD_40M_FIXED[9]_net_1\);
    
    \REG40M.SEQCNTS_30[4]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[4]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_8, E => N_286, Q => \SEQCNTS_30[4]\);
    
    \REG40M.BIT_OS_VAL_29_RNIMHLG[0]\ : MX2
      port map(A => \BIT_OS_VAL_13[0]\, B => \BIT_OS_VAL_29[0]\, 
        S => \CLKPHASE_5[4]_net_1\, Y => N_3643);
    
    \REG40M.BIT_OS_CNT_4[8]\ : DFN1E1C0
      port map(D => N_35, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_9, E => BIT_OS_CNT_4e, Q => 
        \BIT_OS_CNT_4[8]\);
    
    \REG40M.BIT_OS_CNT_2_RNO[6]\ : XA1B
      port map(A => BIT_OS_CNT_2_c5, B => \BIT_OS_CNT_2[6]\, C
         => N_4530_0, Y => BIT_OS_CNT_2_n6);
    
    \SYNC_SM.n_best_clkphase14_0_I_6\ : OA1A
      port map(A => \BEST_SEQCNT[3]_net_1\, B => 
        \un6_n_best_seqcnt[3]\, C => N_3_0, Y => N_7);
    
    \REG40M.SEQCNTS_15[1]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[1]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_4, E => N_316, Q => \SEQCNTS_15[1]\);
    
    \REG40M.BIT_OS_VAL_17[2]\ : DFN1E1C0
      port map(D => N_187, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_18, E => \DES_SM_3[6]_net_1\, Q => 
        \BIT_OS_VAL_17[2]\);
    
    \DES_SM_RNO[7]\ : AO1B
      port map(A => \DES_SM_ns_i_a2_i_a3_0[1]\, B => N_116, C => 
        N_54, Y => N_49);
    
    \REG40M.BIT_OS_CNT_1_RNIUUE8[2]\ : OR3C
      port map(A => \BIT_OS_CNT_1[1]\, B => \BIT_OS_CNT_1[2]\, C
         => \BIT_OS_CNT_1[0]\, Y => N_428);
    
    \REG40M.SEQCNTS_15[2]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[2]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_4, E => N_316, Q => \SEQCNTS_15[2]\);
    
    \REG40M.BIT_OS_VAL_4_RNO[3]\ : MX2
      port map(A => N_209_0, B => \BIT_OS_VAL_4[3]\, S => N_5674, 
        Y => \N_BIT_OS_VAL_4_18[3]\);
    
    \BEST_CLKPHASE[0]\ : DFN1E1C0
      port map(D => \N_BEST_CLKPHASE[0]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_10, E => un1_N_CCC_RESET_EN_0_sqmuxa, 
        Q => \BEST_CLKPHASE[0]_net_1\);
    
    \REG40M.SEQCNTS_1_RNIPS9K[4]\ : MX2
      port map(A => \SEQCNTS_1[4]\, B => \SEQCNTS_2[4]\, S => 
        \INDEX_CNT_1[0]_net_1\, Y => N_4002);
    
    \DES_SM_0_RNISKC8K[8]\ : NOR2A
      port map(A => I_5, B => \DES_SM_0[8]_net_1\, Y => 
        \N_SEQCNTS_1_0[1]\);
    
    \REG40M.SEQCNTS_11_RNIQ6U81[2]\ : MX2
      port map(A => \SEQCNTS_11[2]\, B => \SEQCNTS_12[2]\, S => 
        \INDEX_CNT_4[0]_net_1\, Y => N_4075);
    
    \REG40M.BIT_OS_VAL_5_RNO[1]\ : MX2B
      port map(A => \BIT_OS_VAL_5[1]\, B => N_206, S => 
        \un36_n_bit_os_val[26]\, Y => \N_BIT_OS_VAL_5_18[1]\);
    
    \CLKPHASE_2_RNIIIBG1[3]\ : MX2
      port map(A => N_3817, B => N_3822, S => 
        \CLKPHASE_2[3]_net_1\, Y => N_3827);
    
    \ARB_BYTE_RNIAIJU[2]\ : NOR3B
      port map(A => \ARB_BYTE[5]_net_1\, B => N_771, C => 
        \ARB_BYTE[2]_net_1\, Y => N_561_3);
    
    \CLKPHASE_0_RNIA5411[3]\ : MX2
      port map(A => N_3639, B => N_3643, S => 
        \CLKPHASE_0[3]_net_1\, Y => N_3647);
    
    \BEST_BIT_OS_VAL_RNO_9[0]\ : MX2
      port map(A => N_3906, B => N_3910, S => 
        \INDEX_CNT_2[3]_net_1\, Y => N_3914);
    
    \WAITCNT_RNIH5MR[3]\ : NOR3C
      port map(A => \WAITCNT[4]_net_1\, B => \WAITCNT[3]_net_1\, 
        C => \WAITCNT[13]_net_1\, Y => 
        un1_DES_SM_471_i_0_a2_0_0_a2_6);
    
    \REG40M.SEQCNTS_19_RNI6RGG[4]\ : MX2
      port map(A => \SEQCNTS_3[4]\, B => \SEQCNTS_19[4]\, S => 
        \CLKPHASE_1[4]_net_1\, Y => N_3742);
    
    \DES_SM_RNI5LBTT[8]\ : NOR2A
      port map(A => I_7, B => \DES_SM[8]_net_1\, Y => 
        \N_SEQCNTS_1[2]\);
    
    un1_N_CCC_RESET_EN_0_sqmuxa_0_0_o2 : NOR2B
      port map(A => \DES_SM[8]_net_1\, B => OP_MODE_c_0, Y => 
        N_5784_i);
    
    \REG40M.BIT_OS_CNT_4_RNI0IBO7[4]\ : OR2
      port map(A => N_360, B => N_437, Y => N_781);
    
    \DES_SM_RNICU2EH7[8]\ : AO1
      port map(A => \un36_n_bit_os_val[9]\, B => N_782, C => 
        N_717, Y => N_302);
    
    \ARB_BYTE_RNI82M33_0[1]\ : AO1
      port map(A => BIT_OS_CNT_0lde_0_a3_1, B => 
        BIT_OS_CNT_0lde_0_a3_0, C => N_4530_1, Y => BIT_OS_CNT_0e);
    
    \REG40M.BIT_OS_VAL_7_RNO[2]\ : MX2
      port map(A => \BIT_OS_VAL_7[2]\, B => N_781, S => 
        \un36_n_bit_os_val[24]\, Y => N_205);
    
    \REG40M.SEQCNTS_7_RNIDD051[0]\ : MX2
      port map(A => \SEQCNTS_7[0]\, B => \SEQCNTS_8[0]\, S => 
        \INDEX_CNT[0]_net_1\, Y => N_4083);
    
    \REG40M.BIT_OS_VAL_18_RNO[1]\ : MX2B
      port map(A => \BIT_OS_VAL_18[1]\, B => N_206_0, S => 
        \un36_n_bit_os_val[13]\, Y => \N_BIT_OS_VAL_18_18[1]\);
    
    \REG40M.BIT_OS_VAL_0_RNISTDN[1]\ : MX2
      port map(A => \BIT_OS_VAL_0[1]\, B => \BIT_OS_VAL_16[1]\, S
         => \CLKPHASE_1[4]_net_1\, Y => N_3660);
    
    \REG40M.SEQCNTS_21_RNIN77G[0]\ : MX2
      port map(A => \SEQCNTS_21[0]\, B => \SEQCNTS_22[0]\, S => 
        \INDEX_CNT_3[0]_net_1\, Y => N_4048);
    
    \REG40M.BIT_OS_VAL_12[2]\ : DFN1E1C0
      port map(D => N_195, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_10, E => \DES_SM_2[6]_net_1\, Q => 
        \BIT_OS_VAL_12[2]\);
    
    \REG40M.SEQCNTS_6[4]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[4]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_16, E => N_334, Q => \SEQCNTS_6[4]\);
    
    \REG40M.BIT_OS_VAL_20[1]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_20_18[1]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_13, E => \DES_SM_2[6]_net_1\, Q
         => \BIT_OS_VAL_20[1]\);
    
    \REG40M.BIT_OS_CNT_3_RNI21431[6]\ : NOR2B
      port map(A => BIT_OS_CNT_3_c5, B => \BIT_OS_CNT_3[6]\, Y
         => BIT_OS_CNT_3_c6);
    
    \REG40M.BIT_OS_CNT_6[2]\ : DFN1E1C0
      port map(D => N_83, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_12, E => BIT_OS_CNT_6e, Q => 
        \BIT_OS_CNT_6[2]\);
    
    \BEST_BIT_OS_VAL_RNO_2[0]\ : MX2
      port map(A => N_3958, B => N_3986, S => 
        \INDEX_CNT[4]_net_1\, Y => N_3990);
    
    \REG40M.BIT_OS_CNT_6_RNIRQTO[8]\ : OR3
      port map(A => \BIT_OS_CNT_6[4]\, B => \BIT_OS_CNT_6[5]\, C
         => \BIT_OS_CNT_6[8]\, Y => N_BIT_OS_VAL_3126lto8_0_o3_0);
    
    \INDEX_CNT[0]\ : DFN1E0C0
      port map(D => \N_INDEX_CNT[0]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_16_0, E => N_5149, Q => 
        \INDEX_CNT[0]_net_1\);
    
    \ARB_BYTE_RNI3N9F_0[0]\ : NOR2A
      port map(A => \ARB_BYTE[3]_net_1\, B => \ARB_BYTE[0]_net_1\, 
        Y => N_771);
    
    \REG40M.BIT_OS_CNT_1[6]\ : DFN1E1C0
      port map(D => N_129, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_4, E => BIT_OS_CNT_1e, Q => 
        \BIT_OS_CNT_1[6]\);
    
    \REG40M.BIT_OS_CNT_0[5]\ : DFN1E1C0
      port map(D => N_113, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_3, E => BIT_OS_CNT_0e, Q => 
        \BIT_OS_CNT_0[5]\);
    
    \WAITCNT_RNO[4]\ : XA1C
      port map(A => \WAITCNT[4]_net_1\, B => N_5774, C => N_4539, 
        Y => N_37);
    
    \ARB_WRD_40M_FIXED[8]\ : DFN1C0
      port map(D => \Q[8]_net_1\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_26, Q => \ARB_WRD_40M_FIXED[8]_net_1\);
    
    \BIT_OS_SEL_3[0]\ : DFN1C0
      port map(D => \BEST_BIT_OS_VAL[0]_net_1\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_27_0, Q => BIT_OS_SEL_3(0));
    
    \REG40M.BIT_OS_CNT_7_RNO[8]\ : XA1B
      port map(A => BIT_OS_CNT_7_360_0, B => \BIT_OS_CNT_7[8]\, C
         => N_4530_2, Y => BIT_OS_CNT_7_n8);
    
    \CLKPHASE_RNI0GB33[2]\ : MX2
      port map(A => N_3698, B => N_3710, S => \CLKPHASE[2]_net_1\, 
        Y => N_3714);
    
    \BEST_BIT_OS_VAL_RNO_5[3]\ : MX2
      port map(A => N_3945, B => N_3957, S => 
        \INDEX_CNT_0[2]_net_1\, Y => N_3961);
    
    \SYNC_SM.N_TUNE_CLKPHASE_2_0_0_ADD_5x5_slow_I3_S\ : XNOR3
      port map(A => \BEST_SEQCNT[4]_net_1\, B => 
        \BEST_CLKPHASE[3]_net_1\, C => I2_un1_CO1, Y => 
        \N_TUNE_CLKPHASE_2[3]\);
    
    \CLKPHASE_RNI28EF1[3]\ : MX2
      port map(A => N_3837, B => N_3842, S => \CLKPHASE[3]_net_1\, 
        Y => N_3847);
    
    \CLKPHASE_RNIP0JI_2[1]\ : NOR2B
      port map(A => N_5712, B => N_215, Y => 
        \un36_n_bit_os_val[4]\);
    
    \RECD_SER_WORD_RNO_4[2]\ : NOR3C
      port map(A => n_recd_ser_word168_2, B => 
        n_recd_ser_word169_0, C => \ARB_BYTE[7]_net_1\, Y => 
        \ARB_BYTE_m_1[7]\);
    
    \RECD_SER_WORD[7]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[7]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_30, Q => \RECD_SER_WORD[7]_net_1\);
    
    \SYNC_SM.N_TUNE_CLKPHASE_2_0_0_ALL_PLL_LOCK\ : NOR2B
      port map(A => CCC_MAIN_LOCK, B => CCC_RX_CLK_LOCK, Y => 
        ALL_PLL_LOCK_c);
    
    \REG40M.BIT_OS_VAL_3_RNI3N911[0]\ : MX2
      port map(A => \BIT_OS_VAL_3[0]\, B => \BIT_OS_VAL_19[0]\, S
         => \CLKPHASE_4[4]_net_1\, Y => N_3611);
    
    un41_n_seqcnts_I_6 : NOR2B
      port map(A => \un39_n_seqcnts[1]\, B => \un39_n_seqcnts[0]\, 
        Y => N_4);
    
    \ARB_BYTE[10]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[10]_net_1\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_32_0, Q => 
        \ARB_BYTE[10]_net_1\);
    
    \WAITCNT[9]\ : DFN1E0C0
      port map(D => N_5810, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_9, E => N_5790, Q => \WAITCNT[9]_net_1\);
    
    \REG40M.SEQCNTS_30_RNI1KVA[4]\ : MX2
      port map(A => \SEQCNTS_14[4]\, B => \SEQCNTS_30[4]\, S => 
        \CLKPHASE[4]_net_1\, Y => N_3857);
    
    \RECD_SER_WORD_RNIIIBK[5]\ : NOR2B
      port map(A => \RECD_SER_WORD[5]_net_1\, B => DCB_SALT_SEL_c, 
        Y => \ELK_RX_SER_WORD_0[5]\);
    
    \CLKPHASE_RNIP0JI_6[0]\ : NOR2B
      port map(A => N_5711, B => N_214, Y => 
        \un36_n_bit_os_val[16]\);
    
    \CLKPHASE_RNIP0JI_1[0]\ : NOR3B
      port map(A => \CLKPHASE[0]_net_1\, B => N_204, C => N_90, Y
         => \un36_n_bit_os_val[10]\);
    
    \CLKPHASE[2]\ : DFN1C0
      port map(D => \TUNE_CLKPHASE_RNIDA643[2]_net_1\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_24_0, Q => 
        \CLKPHASE[2]_net_1\);
    
    \BEST_BIT_OS_VAL_RNO_9[1]\ : MX2
      port map(A => N_3907, B => N_3911, S => 
        \INDEX_CNT_2[3]_net_1\, Y => N_3915);
    
    \REG40M.SEQCNTS_27[0]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[0]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_13, E => N_292, Q => \SEQCNTS_27[0]\);
    
    \RECD_SER_WORD_RNO_0[1]\ : AO1
      port map(A => n_recd_ser_word170, B => \ARB_BYTE[7]_net_1\, 
        C => \ARB_BYTE_m[8]\, Y => \N_RECD_SER_WORD_iv_1[1]\);
    
    \DES_SM_0_RNIAB7UH7_5[8]\ : AO1
      port map(A => \un36_n_bit_os_val[24]\, B => N_782_0, C => 
        N_717_0, Y => N_332);
    
    \TUNE_CLKPHASE_RNI79F03[1]\ : AO1A
      port map(A => N_5780, B => \TUNE_CLKPHASE[1]_net_1\, C => 
        N_5793, Y => \TUNE_CLKPHASE_RNI79F03[1]_net_1\);
    
    \CLKPHASE_RNICU2EH7_0[1]\ : AO1
      port map(A => \un36_n_bit_os_val[6]\, B => N_782, C => 
        N_717, Y => N_296);
    
    \CLKPHASE_0_RNIUNTU[3]\ : MX2
      port map(A => N_3641, B => N_3645, S => 
        \CLKPHASE_0[3]_net_1\, Y => N_3649);
    
    \RECD_SER_WORD_RNIHHBK_0[4]\ : NOR2A
      port map(A => \RECD_SER_WORD[4]_net_1\, B => DCB_SALT_SEL_c, 
        Y => TFC_RX_SER_WORD(4));
    
    \DES_SM_RNICU2EH7_1[8]\ : AO1
      port map(A => \un36_n_bit_os_val[12]\, B => N_782, C => 
        N_717, Y => N_308);
    
    \REG40M.SEQCNTS_20_RNI3JAG[4]\ : MX2
      port map(A => \SEQCNTS_4[4]\, B => \SEQCNTS_20[4]\, S => 
        \CLKPHASE_5[4]_net_1\, Y => N_3817);
    
    \REG40M.BIT_OS_VAL_10_RNIJSPM[3]\ : MX2
      port map(A => \BIT_OS_VAL_10[3]\, B => \BIT_OS_VAL_26[3]\, 
        S => \CLKPHASE_2[4]_net_1\, Y => N_3694);
    
    \RECD_SER_WORD_RNO_4[3]\ : NOR3C
      port map(A => n_recd_ser_word168_2, B => 
        n_recd_ser_word169_0, C => \ARB_BYTE[8]_net_1\, Y => 
        \ARB_BYTE_m_1[8]\);
    
    \ARB_BYTE_RNI2M9F[0]\ : NOR2A
      port map(A => \ARB_BYTE[2]_net_1\, B => \ARB_BYTE[0]_net_1\, 
        Y => BIT_OS_CNT_3lde_0_a3_0);
    
    un1_DES_SM_1003_i_0 : OR2
      port map(A => N_128, B => N_5792, Y => N_5724);
    
    \RECD_SER_WORD_RNI01N81[0]\ : NOR2
      port map(A => \ELK_RX_SER_WORD_0[0]\, B => 
        \ELK_RX_SER_WORD_0[6]\, Y => ELK0_SYNC_DET_1_2);
    
    un1_CLKPHASE_I_28 : AND2
      port map(A => \CLKPHASE[2]_net_1\, B => \CLKPHASE[3]_net_1\, 
        Y => \DWACT_ADD_CI_0_pog_array_1[0]\);
    
    CONFIG_ONCE_TRIG_RNO : AO1A
      port map(A => \DES_SM_0[8]_net_1\, B => 
        N_CONFIG_ONCE_TRIG_i_a3_0, C => N_140, Y => N_58);
    
    \INDEX_CNT_0[0]\ : DFN1E0C0
      port map(D => \N_INDEX_CNT[0]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_16_0, E => N_5149, Q => 
        \INDEX_CNT_0[0]_net_1\);
    
    \REG40M.BIT_OS_VAL_3_RNO[0]\ : MX2
      port map(A => N_5666, B => \BIT_OS_VAL_3[0]\, S => N_5675, 
        Y => \N_BIT_OS_VAL_3_18[0]\);
    
    \INDEX_CNT_1_RNIC9VM1[3]\ : MX2
      port map(A => N_4034, B => N_4039, S => 
        \INDEX_CNT_1[3]_net_1\, Y => N_4044);
    
    \REG40M.BIT_OS_VAL_28_RNO[1]\ : MX2B
      port map(A => \BIT_OS_VAL_28[1]\, B => N_206, S => 
        \un36_n_bit_os_val[3]\, Y => \N_BIT_OS_VAL_28_18[1]\);
    
    \REG40M.BIT_OS_VAL_18[0]\ : DFN1E1C0
      port map(D => N_249, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_19, E => \DES_SM_4[6]_net_1\, Q => 
        \BIT_OS_VAL_18[0]\);
    
    \REG40M.SEQCNTS_13_RNIRD7C[1]\ : MX2
      port map(A => \SEQCNTS_13[1]\, B => \SEQCNTS_14[1]\, S => 
        \INDEX_CNT_3[0]_net_1\, Y => N_4019);
    
    \CLKPHASE_0_RNIDA401[3]\ : MX2
      port map(A => N_3848, B => N_3853, S => 
        \CLKPHASE_0[3]_net_1\, Y => N_3858);
    
    \REG40M.BIT_OS_VAL_26[2]\ : DFN1E1C0
      port map(D => N_169, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_21, E => \DES_SM[6]_net_1\, Q => 
        \BIT_OS_VAL_26[2]\);
    
    \REG40M.BIT_OS_VAL_13[1]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_13_18[1]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_12, E => \DES_SM_2[6]_net_1\, Q
         => \BIT_OS_VAL_13[1]\);
    
    \REG40M.SEQCNTS_6[1]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[1]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_16, E => N_334, Q => \SEQCNTS_6[1]\);
    
    \Q[14]\ : DFN1C0
      port map(D => \ADJ_Q[14]_net_1\, CLK => CCC_160M_FXD, CLR
         => P_MASTER_POR_B_c_23, Q => \Q[14]_net_1\);
    
    \REG40M.BIT_OS_CNT_2_RNIK7CV[1]\ : OR3
      port map(A => N_BIT_OS_VAL_3110lt8, B => 
        N_BIT_OS_VAL_3110lto8_1, C => N_BIT_OS_VAL_3110lto8_2, Y
         => N_BIT_OS_VAL_3110);
    
    \REG40M.SEQCNTS_29[3]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[3]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_16_0, E => N_288, Q => \SEQCNTS_29[3]\);
    
    \CLKPHASE_RNIQVDF1[3]\ : MX2
      port map(A => N_3835, B => N_3840, S => \CLKPHASE[3]_net_1\, 
        Y => N_3845);
    
    \REG40M.SEQCNTS_29_RNI26G41[1]\ : MX2
      port map(A => N_4049, B => \SEQCNTS_29[1]\, S => 
        \INDEX_CNT_2[3]_net_1\, Y => N_4054);
    
    \REG40M.BIT_OS_CNT_0_RNI4NQD[1]\ : OR3
      port map(A => N_750, B => N_BIT_OS_VAL_312lto8_0_o3_1, C
         => N_BIT_OS_VAL_312lto8_0_o3_2, Y => N_BIT_OS_VAL_312);
    
    \RECD_SER_WORD_RNO_4[4]\ : NOR3C
      port map(A => n_recd_ser_word168_2, B => 
        n_recd_ser_word169_0, C => \ARB_BYTE[9]_net_1\, Y => 
        \ARB_BYTE_m_1[9]\);
    
    \BEST_BIT_OS_VAL_RNO_20[0]\ : MX2
      port map(A => \BIT_OS_VAL_25[0]\, B => \BIT_OS_VAL_26[0]\, 
        S => \INDEX_CNT_3[0]_net_1\, Y => N_3910);
    
    \BEST_BIT_OS_VAL_RNO_22[1]\ : MX2
      port map(A => \BIT_OS_VAL_3[1]\, B => \BIT_OS_VAL_4[1]\, S
         => \INDEX_CNT_0[0]_net_1\, Y => N_3935);
    
    \REG40M.BIT_OS_CNT_0_RNIUO55[1]\ : NOR3C
      port map(A => \BIT_OS_CNT_0[2]\, B => \BIT_OS_CNT_0[1]\, C
         => \BIT_OS_CNT_0[3]\, Y => N_750);
    
    \REG40M.BIT_OS_CNT_5_RNIQRQS[3]\ : OR2A
      port map(A => \BIT_OS_CNT_5[3]\, B => N_373, Y => N_376);
    
    \REG40M.BIT_OS_CNT_1_RNISM4U2[4]\ : AO1A
      port map(A => N_BIT_OS_VAL_3110, B => N_BIT_OS_VAL_316, C
         => N_BIT_OS_VAL_3114, Y => N_82);
    
    \REG40M.SEQCNTS_24[3]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[3]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_8, E => N_298, Q => \SEQCNTS_24[3]\);
    
    \REG40M.SEQCNTS_13_RNI1K7C[4]\ : MX2
      port map(A => \SEQCNTS_13[4]\, B => \SEQCNTS_14[4]\, S => 
        \INDEX_CNT_3[0]_net_1\, Y => N_4022);
    
    \REG40M.BIT_OS_CNT_4[4]\ : DFN1E1C0
      port map(D => N_5623, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_9, E => BIT_OS_CNT_4e, Q => 
        \BIT_OS_CNT_4[4]\);
    
    \REG40M.SEQCNTS_15_RNIQEAD[0]\ : MX2
      port map(A => \SEQCNTS_15[0]\, B => \SEQCNTS_16[0]\, S => 
        \INDEX_CNT_0[0]_net_1\, Y => N_4088);
    
    \CLKPHASE_1_RNIHE5C1[3]\ : MX2
      port map(A => N_3742, B => N_3747, S => 
        \CLKPHASE_1[3]_net_1\, Y => N_3752);
    
    \REG40M.SEQCNTS_27[1]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[1]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_13, E => N_292, Q => \SEQCNTS_27[1]\);
    
    \REG40M.BIT_OS_VAL_25[1]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_25_18[1]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_20, E => \DES_SM[6]_net_1\, Q => 
        \BIT_OS_VAL_25[1]\);
    
    \CLKPHASE_RNIB6EBB[0]\ : MX2
      port map(A => N_3658, B => N_3718, S => \CLKPHASE[0]_net_1\, 
        Y => \un107_bit_os_val[3]\);
    
    \BEST_BIT_OS_VAL_RNO_29[3]\ : MX2
      port map(A => \BIT_OS_VAL_31[3]\, B => \BIT_OS_VAL_0[3]\, S
         => \INDEX_CNT_3[0]_net_1\, Y => N_3981);
    
    \REG40M.BIT_OS_VAL_30[0]\ : DFN1E1C0
      port map(D => N_213, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_18, E => \DES_SM_4[6]_net_1\, Q => 
        \BIT_OS_VAL_30[0]\);
    
    \REG40M.BIT_OS_CNT_0_RNIHDE3[0]\ : OR2B
      port map(A => \BIT_OS_CNT_0[1]\, B => \BIT_OS_CNT_0[0]\, Y
         => N_368);
    
    \MAX_CNT_RNO[5]\ : XA1C
      port map(A => \MAX_CNT[5]_net_1\, B => N_385, C => 
        un1_DES_SM_19, Y => N_5635);
    
    \WAITCNT_RNO_0[8]\ : OA1C
      port map(A => \WAITCNT[7]_net_1\, B => N_5777, C => 
        \WAITCNT[8]_net_1\, Y => N_5807);
    
    \REG40M.BIT_OS_CNT_4_RNIMFEO[0]\ : OR2A
      port map(A => \BIT_OS_CNT_4[0]\, B => N_363, Y => N_379);
    
    \BEST_CLKPHASE_RNO[2]\ : NOR2A
      port map(A => I_7_0, B => \DES_SM_1[8]_net_1\, Y => 
        \N_BEST_CLKPHASE[2]\);
    
    \REG40M.BIT_OS_VAL_29_RNIOJLG[1]\ : MX2
      port map(A => \BIT_OS_VAL_13[1]\, B => \BIT_OS_VAL_29[1]\, 
        S => \CLKPHASE_5[4]_net_1\, Y => N_3644);
    
    \CLKPHASE[1]\ : DFN1C0
      port map(D => \TUNE_CLKPHASE_RNI79F03[1]_net_1\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_24_0, Q => 
        \CLKPHASE[1]_net_1\);
    
    \PHASE_ADJ[1]\ : DFN1C0
      port map(D => \CLKPHASE[1]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c, Q => PHASE_ADJ_160_L(1));
    
    \REG40M.SEQCNTS_30_RNIRDVA[1]\ : MX2
      port map(A => \SEQCNTS_14[1]\, B => \SEQCNTS_30[1]\, S => 
        \CLKPHASE[4]_net_1\, Y => N_3854);
    
    \REG40M.BIT_OS_VAL_27[2]\ : DFN1E1C0
      port map(D => N_167, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_2, E => \DES_SM_0[6]_net_1\, Q => 
        \BIT_OS_VAL_27[2]\);
    
    \DES_SM_RNIK5SE_0[8]\ : NOR2A
      port map(A => \DES_SM[8]_net_1\, B => \DES_SM[6]_net_1\, Y
         => N_717);
    
    \REG40M.BIT_OS_VAL_14_RNO[0]\ : MX2
      port map(A => N_5666_0, B => \BIT_OS_VAL_14[0]\, S => 
        N_5673, Y => \N_BIT_OS_VAL_14_18[0]\);
    
    \RECD_SER_WORD_RNO_3[4]\ : NOR3C
      port map(A => n_recd_ser_word167_1, B => 
        n_recd_ser_word171_0, C => \ARB_BYTE[11]_net_1\, Y => 
        \ARB_BYTE_m[11]\);
    
    \REG40M.SEQCNTS_23_RNIUFDH[1]\ : MX2
      port map(A => \SEQCNTS_7[1]\, B => \SEQCNTS_23[1]\, S => 
        \CLKPHASE_0[4]_net_1\, Y => N_3729);
    
    \REG40M.BIT_OS_CNT_6_RNIG9ND4[7]\ : OR2
      port map(A => N_BIT_OS_VAL_3126, B => N_BIT_OS_VAL_3130, Y
         => N_360);
    
    \INDEX_CNT_RNIAE2N4[2]\ : MX2
      port map(A => N_4078, B => N_4093, S => 
        \INDEX_CNT[2]_net_1\, Y => N_4098);
    
    \CLKPHASE_0_RNIJ80G2[2]\ : MX2
      port map(A => N_3843, B => N_3858, S => 
        \CLKPHASE_0[2]_net_1\, Y => N_3863);
    
    \INDEX_CNT_0_RNI3ATE3[2]\ : MX2
      port map(A => N_4115, B => N_4130, S => 
        \INDEX_CNT_0[2]_net_1\, Y => N_4135);
    
    \WAITCNT_RNIOU3P[1]\ : NOR3C
      port map(A => \WAITCNT[1]_net_1\, B => \WAITCNT[7]_net_1\, 
        C => un1_DES_SM_471_i_0_a2_0_0_a2_2, Y => 
        un1_DES_SM_471_i_0_a2_0_0_a2_7);
    
    \REG40M.SEQCNTS_4[0]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[0]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_13, E => N_338, Q => \SEQCNTS_4[0]\);
    
    \REG40M.SEQCNTS_14[1]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[1]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_2, E => N_318, Q => \SEQCNTS_14[1]\);
    
    \REG40M.SEQCNTS_31_RNIGO4I[3]\ : NOR2A
      port map(A => \SEQCNTS_31[3]\, B => \INDEX_CNT[0]_net_1\, Y
         => N_4126);
    
    \WAITCNT[10]\ : DFN1E0C0
      port map(D => N_5811, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_21, E => N_5790, Q => 
        \WAITCNT[10]_net_1\);
    
    \WAITCNT_RNI7V292[8]\ : NOR3C
      port map(A => \DES_SM_ns_0_0_0_a2_1[0]\, B => 
        \DES_SM_ns_0_0_0_a2_0[0]\, C => \DES_SM_ns_0_0_0_a2_2[0]\, 
        Y => \DES_SM_ns_0_0_0_a2_4[0]\);
    
    \BEST_BIT_OS_VAL_RNO_5[2]\ : MX2
      port map(A => N_3944, B => N_3956, S => 
        \INDEX_CNT_0[2]_net_1\, Y => N_3960);
    
    \REG40M.SEQCNTS_16_RNI7JH7[4]\ : NOR2B
      port map(A => \SEQCNTS_16[4]\, B => \CLKPHASE[4]_net_1\, Y
         => N_3802);
    
    \DES_SM[7]\ : DFN1C0
      port map(D => N_49, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_27, Q => \DES_SM[7]_net_1\);
    
    \ARB_WRD_40M_FIXED[14]\ : DFN1C0
      port map(D => \Q[14]_net_1\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_28, Q => \ARB_WRD_40M_FIXED[14]_net_1\);
    
    \REG40M.BIT_OS_VAL_22[2]\ : DFN1E1C0
      port map(D => N_177, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_15, E => \DES_SM_3[6]_net_1\, Q => 
        \BIT_OS_VAL_22[2]\);
    
    \REG40M.BIT_OS_VAL_30_RNIDNSP[0]\ : MX2
      port map(A => \BIT_OS_VAL_14[0]\, B => \BIT_OS_VAL_30[0]\, 
        S => \CLKPHASE_3[4]_net_1\, Y => N_3703);
    
    \REG40M.BIT_OS_CNT_3[0]\ : DFN1E1C0
      port map(D => N_5619, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_7, E => BIT_OS_CNT_3e, Q => 
        \BIT_OS_CNT_3[0]\);
    
    \INDEX_CNT_RNI9AST1[3]\ : MX2
      port map(A => N_4104, B => N_4109, S => 
        \INDEX_CNT[3]_net_1\, Y => N_4114);
    
    \CLKPHASE_RNICT4B[1]\ : NOR2A
      port map(A => \CLKPHASE[1]_net_1\, B => N_5668, Y => N_5712);
    
    \REG40M.BIT_OS_VAL_7_RNI4N9J[1]\ : MX2
      port map(A => \BIT_OS_VAL_7[1]\, B => \BIT_OS_VAL_23[1]\, S
         => \CLKPHASE_4[4]_net_1\, Y => N_3604);
    
    \BEST_BIT_OS_VAL_RNO_23[2]\ : MX2
      port map(A => \BIT_OS_VAL_11[2]\, B => \BIT_OS_VAL_12[2]\, 
        S => \INDEX_CNT_1[0]_net_1\, Y => N_3940);
    
    \BEST_BIT_OS_VAL_RNO_21[2]\ : MX2
      port map(A => \BIT_OS_VAL_21[2]\, B => \BIT_OS_VAL_22[2]\, 
        S => \INDEX_CNT[0]_net_1\, Y => N_3920);
    
    \BEST_BIT_OS_VAL_RNO_11[0]\ : MX2
      port map(A => N_3934, B => N_3938, S => 
        \INDEX_CNT_0[3]_net_1\, Y => N_3942);
    
    \REG40M.BIT_OS_VAL_9_RNO[2]\ : MX2
      port map(A => \BIT_OS_VAL_9[2]\, B => N_781, S => 
        \un36_n_bit_os_val[22]\, Y => N_201);
    
    \ARB_BYTE[1]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[1]_net_1\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_27, Q => 
        \ARB_BYTE[1]_net_1\);
    
    \REG40M.BIT_OS_CNT_6_RNO[4]\ : XA1C
      port map(A => N_378, B => \BIT_OS_CNT_6[4]\, C => N_4530_1, 
        Y => N_79);
    
    \DES_SM_0[8]\ : DFN1P0
      port map(D => \DES_SM_ns[0]\, CLK => CLK_40M_GL, PRE => 
        P_MASTER_POR_B_c_27_1, Q => \DES_SM_0[8]_net_1\);
    
    \REG40M.BIT_OS_CNT_3_RNI7K1F[2]\ : NOR3C
      port map(A => \BIT_OS_CNT_3[2]\, B => \BIT_OS_CNT_3[3]\, C
         => \BIT_OS_CNT_3[1]\, Y => N_BIT_OS_VAL_3114lt8);
    
    \REG40M.SEQCNTS_14[4]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[4]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_2, E => N_318, Q => \SEQCNTS_14[4]\);
    
    \REG40M.SEQCNTS_18[3]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[3]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_8, E => N_310, Q => \SEQCNTS_18[3]\);
    
    \REG40M.BIT_OS_CNT_3[8]\ : DFN1E1C0
      port map(D => BIT_OS_CNT_3_n8, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_7, E => BIT_OS_CNT_3e, Q => 
        \BIT_OS_CNT_3[8]\);
    
    \REG40M.SEQCNTS_11_RNIM2U81[0]\ : MX2
      port map(A => \SEQCNTS_11[0]\, B => \SEQCNTS_12[0]\, S => 
        \INDEX_CNT_4[0]_net_1\, Y => N_4073);
    
    \REG40M.BIT_OS_CNT_7_RNO[1]\ : XA1B
      port map(A => \BIT_OS_CNT_7[1]\, B => \BIT_OS_CNT_7[0]\, C
         => N_4530_2, Y => BIT_OS_CNT_7_n1);
    
    \MAX_CNT_RNIG67M[5]\ : NOR2
      port map(A => \MAX_CNT[5]_net_1\, B => \MAX_CNT[7]_net_1\, 
        Y => DES_SM_tr2_i_a3_2);
    
    \DES_SM_RNIFA8R[0]\ : MX2A
      port map(A => \DES_SM[0]_net_1\, B => OP_MODE_c_0, S => 
        \DES_SM_0[8]_net_1\, Y => N_5780);
    
    \REG40M.BIT_OS_CNT_7_RNIULQ12[6]\ : NOR2B
      port map(A => BIT_OS_CNT_7_c5, B => \BIT_OS_CNT_7[6]\, Y
         => BIT_OS_CNT_7_c6);
    
    \DES_SM_RNO_0[7]\ : NOR2B
      port map(A => CCC_RX_CLK_LOCK, B => N_70, Y => 
        \DES_SM_ns_i_a2_i_a3_0[1]\);
    
    \CLKPHASE_1_RNIDA5C1[3]\ : MX2
      port map(A => N_3741, B => N_3746, S => 
        \CLKPHASE_1[3]_net_1\, Y => N_3751);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \RECD_SER_WORD_RNIEEBK[1]\ : NOR2B
      port map(A => \RECD_SER_WORD[1]_net_1\, B => DCB_SALT_SEL_c, 
        Y => ELK_RX_SER_WORD_0(1));
    
    \DES_SM_2[6]\ : DFN1C0
      port map(D => N_MAX_CNT_0_sqmuxa, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_27_1, Q => \DES_SM_2[6]_net_1\);
    
    \ARB_WRD_40M_FIXED[1]\ : DFN1C0
      port map(D => \Q[1]_net_1\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_26, Q => \ARB_WRD_40M_FIXED[1]_net_1\);
    
    \REG40M.BIT_OS_VAL_30[3]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_30_18[3]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_18, E => \DES_SM_4[6]_net_1\, Q
         => \BIT_OS_VAL_30[3]\);
    
    \REG40M.BIT_OS_VAL_1_RNIV2HO[2]\ : MX2
      port map(A => \BIT_OS_VAL_1[2]\, B => \BIT_OS_VAL_17[2]\, S
         => \CLKPHASE_0[4]_net_1\, Y => N_3629);
    
    \CLKPHASE_RNIO7B33[2]\ : MX2
      port map(A => N_3697, B => N_3709, S => \CLKPHASE[2]_net_1\, 
        Y => N_3713);
    
    \REG40M.BIT_OS_VAL_5_RNI5I0G[3]\ : MX2
      port map(A => \BIT_OS_VAL_5[3]\, B => \BIT_OS_VAL_21[3]\, S
         => \CLKPHASE_5[4]_net_1\, Y => N_3642);
    
    \REG40M.BIT_OS_CNT_5[4]\ : DFN1E1C0
      port map(D => N_5628, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_11, E => BIT_OS_CNT_5e, Q => 
        \BIT_OS_CNT_5[4]\);
    
    \INDEX_CNT[1]\ : DFN1E0C0
      port map(D => \N_INDEX_CNT[1]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_17, E => N_5149, Q => 
        \INDEX_CNT[1]_net_1\);
    
    \DES_SM_0_RNISRO581[8]\ : NOR2A
      port map(A => I_9, B => \DES_SM_0[8]_net_1\, Y => 
        \N_SEQCNTS_1_0[3]\);
    
    \CLKPHASE_1_RNI0S4U[3]\ : MX2
      port map(A => N_3773, B => N_3778, S => 
        \CLKPHASE_1[3]_net_1\, Y => N_3783);
    
    \REG40M.BIT_OS_VAL_24_RNO[0]\ : MX2
      port map(A => \BIT_OS_VAL_24[0]\, B => N_5666_0, S => 
        \un36_n_bit_os_val[7]\, Y => N_231);
    
    \REG40M.BIT_OS_CNT_4_RNO[3]\ : NOR3A
      port map(A => N_379, B => N_504, C => N_4530_0, Y => N_45);
    
    \RECD_SER_WORD_RNO_1[7]\ : AO1
      port map(A => \ARB_BYTE[11]_net_1\, B => n_recd_ser_word168, 
        C => \ARB_BYTE_m_1[12]\, Y => \N_RECD_SER_WORD_iv_0[7]\);
    
    \REG40M.BIT_OS_VAL_6[0]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_6_18[0]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_2, E => \DES_SM_0[6]_net_1\, Q
         => \BIT_OS_VAL_6[0]\);
    
    \REG40M.BIT_OS_CNT_5_RNI7ODE[6]\ : OR2
      port map(A => \BIT_OS_CNT_5[7]\, B => \BIT_OS_CNT_5[6]\, Y
         => N_BIT_OS_VAL_3122lto8_0_o3_1);
    
    \CLKPHASE_RNIVNJCG7[0]\ : OR3
      port map(A => un1_DES_SM_1034_i_o2_1, B => N_754, C => 
        un1_DES_SM_1034_i_o2_2, Y => N_782_0);
    
    \ADJ_Q[3]\ : DFN1C0
      port map(D => \ADJ_Q[1]_net_1\, CLK => CCC_160M_ADJ, CLR
         => P_MASTER_POR_B_c_34_0, Q => \ADJ_Q[3]_net_1\);
    
    \REG40M.BIT_OS_VAL_11_RNO[0]\ : MX2
      port map(A => \BIT_OS_VAL_11[0]\, B => N_5666_0, S => 
        \un36_n_bit_os_val[20]\, Y => N_267);
    
    \REG40M.BIT_OS_CNT_6_RNI32RH1[5]\ : OR3B
      port map(A => \BIT_OS_CNT_6[4]\, B => \BIT_OS_CNT_6[5]\, C
         => N_378, Y => N_387);
    
    \REG40M.BIT_OS_CNT_1_RNO[4]\ : XA1C
      port map(A => \BIT_OS_CNT_1[4]\, B => N_380, C => N_4530_1, 
        Y => N_133);
    
    \INDEX_CNT_0_RNIBR7A1[3]\ : MX2
      port map(A => N_4118, B => N_4123, S => 
        \INDEX_CNT_0[3]_net_1\, Y => N_4128);
    
    \BIT_OS_SEL_4[2]\ : DFN1C0
      port map(D => \BEST_BIT_OS_VAL[2]_net_1\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_27_0, Q => BIT_OS_SEL_4(2));
    
    \REG40M.SEQCNTS_9[0]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[0]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_20, E => N_328, Q => \SEQCNTS_9[0]\);
    
    \REG40M.SEQCNTS_22_RNI7VMK[4]\ : MX2
      port map(A => \SEQCNTS_6[4]\, B => \SEQCNTS_22[4]\, S => 
        \CLKPHASE_5[4]_net_1\, Y => N_3852);
    
    \REG40M.BIT_OS_CNT_3_RNI4H1F[2]\ : NOR3C
      port map(A => \BIT_OS_CNT_3[1]\, B => \BIT_OS_CNT_3[0]\, C
         => \BIT_OS_CNT_3[2]\, Y => BIT_OS_CNT_3_c2);
    
    \INDEX_CNT_0_RNISMFL3[2]\ : MX2
      port map(A => N_4008, B => N_4023, S => 
        \INDEX_CNT_0[2]_net_1\, Y => N_4028);
    
    \DES_SM_RNI74OM_2[7]\ : NOR3A
      port map(A => \DES_SM[7]_net_1\, B => \ARB_BYTE[7]_net_1\, 
        C => \ARB_BYTE[6]_net_1\, Y => N_560_2);
    
    \BEST_BIT_OS_VAL_RNO_4[0]\ : MX2
      port map(A => N_3914, B => N_3922, S => 
        \INDEX_CNT_0[2]_net_1\, Y => N_3926);
    
    \REG40M.BIT_OS_CNT_0[2]\ : DFN1E1C0
      port map(D => N_119, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_3, E => BIT_OS_CNT_0e, Q => 
        \BIT_OS_CNT_0[2]\);
    
    \CLKPHASE_RNIP0JI_2[0]\ : NOR3A
      port map(A => \CLKPHASE[0]_net_1\, B => N_90, C => N_5663, 
        Y => \un36_n_bit_os_val[26]\);
    
    \PHASE_ADJ[0]\ : DFN1C0
      port map(D => \CLKPHASE[0]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c, Q => PHASE_ADJ_160_L(0));
    
    \DES_SM_RNICU2EH7_6[8]\ : AO1
      port map(A => \un36_n_bit_os_val[11]\, B => N_782, C => 
        N_717, Y => N_306);
    
    \ARB_WRD_40M_FIXED[3]\ : DFN1C0
      port map(D => \Q[3]_net_1\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_26, Q => \ARB_WRD_40M_FIXED[3]_net_1\);
    
    \WAITCNT_RNI46UD2[10]\ : OR2A
      port map(A => \WAITCNT[10]_net_1\, B => N_5781, Y => N_5782);
    
    \REG40M.SEQCNTS_1[0]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[0]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_8, E => N_344, Q => \SEQCNTS_1[0]\);
    
    \REG40M.SEQCNTS_23_RNIOAAH[0]\ : MX2
      port map(A => \SEQCNTS_23[0]\, B => \SEQCNTS_24[0]\, S => 
        \INDEX_CNT_0[0]_net_1\, Y => N_4118);
    
    \REG40M.SEQCNTS_15[4]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[4]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_4, E => N_316, Q => \SEQCNTS_15[4]\);
    
    \REG40M.BIT_OS_CNT_3_RNI1N2P[4]\ : NOR3C
      port map(A => \BIT_OS_CNT_3[3]\, B => BIT_OS_CNT_3_c2, C
         => \BIT_OS_CNT_3[4]\, Y => BIT_OS_CNT_3_c4);
    
    \BIT_OS_SEL_0[1]\ : DFN1C0
      port map(D => \BEST_BIT_OS_VAL[1]_net_1\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_27_0, Q => BIT_OS_SEL_0(1));
    
    \BEST_BIT_OS_VAL_RNO_13[0]\ : MX2
      port map(A => N_3962, B => N_3966, S => 
        \INDEX_CNT_1[3]_net_1\, Y => N_3970);
    
    \CLKPHASE_0_RNIND1C[2]\ : OR3A
      port map(A => \CLKPHASE_0[1]_net_1\, B => 
        \CLKPHASE_0[2]_net_1\, C => N_80, Y => N_5678);
    
    \MAX_CNT_RNO[2]\ : NOR3A
      port map(A => N_370, B => N_535, C => un1_DES_SM_19, Y => 
        N_5638);
    
    \DES_SM[0]\ : DFN1C0
      port map(D => \DES_SM_RNO[0]_net_1\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_26, Q => \DES_SM[0]_net_1\);
    
    \REG40M.SEQCNTS_31_RNIDL4I[0]\ : NOR2A
      port map(A => \SEQCNTS_31[0]\, B => \INDEX_CNT[0]_net_1\, Y
         => N_4123);
    
    \REG40M.BIT_OS_VAL_28[0]\ : DFN1E1C0
      port map(D => N_219, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_2, E => \DES_SM_0[6]_net_1\, Q => 
        \BIT_OS_VAL_28[0]\);
    
    \REG40M.BIT_OS_CNT_6_RNO[2]\ : NOR3A
      port map(A => N_430, B => N_525, C => N_4530_1, Y => N_83);
    
    \REG40M.BIT_OS_CNT_4_RNO_0[8]\ : OR2A
      port map(A => \BIT_OS_CNT_4[7]\, B => N_410, Y => N_420);
    
    \INDEX_CNT_1_RNIPO2O1[3]\ : MX2
      port map(A => N_4037, B => N_4042, S => 
        \INDEX_CNT_1[3]_net_1\, Y => N_4047);
    
    \RECD_SER_WORD_RNIFFBK[2]\ : NOR2B
      port map(A => \RECD_SER_WORD[2]_net_1\, B => DCB_SALT_SEL_c, 
        Y => ELK_RX_SER_WORD_0(2));
    
    \SYNC_SM.N_TUNE_CLKPHASE_2_0_0_ADD_5x5_slow_I1_S\ : XNOR3
      port map(A => \BEST_SEQCNT[2]_net_1\, B => 
        \BEST_CLKPHASE[1]_net_1\, C => I0_un1_CO1, Y => 
        \N_TUNE_CLKPHASE_2[1]\);
    
    \CLKPHASE_0_RNIORR71[3]\ : MX2
      port map(A => N_3759, B => N_3764, S => 
        \CLKPHASE_0[3]_net_1\, Y => N_3769);
    
    \REG40M.BIT_OS_VAL_17[3]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_17_18[3]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_18, E => \DES_SM_3[6]_net_1\, Q
         => \BIT_OS_VAL_17[3]\);
    
    \REG40M.BIT_OS_VAL_23[1]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_23_18[1]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_17_0, E => \DES_SM_3[6]_net_1\, Q
         => \BIT_OS_VAL_23[1]\);
    
    \MAX_CNT_RNO_0[8]\ : OR2A
      port map(A => \MAX_CNT[7]_net_1\, B => N_405, Y => N_422);
    
    \REG40M.SEQCNTS_15_RNIAOS9[0]\ : MX2
      port map(A => \SEQCNTS_31[0]\, B => \SEQCNTS_15[0]\, S => 
        \CLKPHASE_0[4]_net_1\, Y => N_3723);
    
    \REG40M.BIT_OS_CNT_6_RNO_0[2]\ : AOI1
      port map(A => \BIT_OS_CNT_6[1]\, B => \BIT_OS_CNT_6[0]\, C
         => \BIT_OS_CNT_6[2]\, Y => N_525);
    
    \ADJ_Q[7]\ : DFN1C0
      port map(D => \ADJ_Q[5]_net_1\, CLK => CCC_160M_ADJ, CLR
         => P_MASTER_POR_B_c_34_0, Q => \ADJ_Q[7]_net_1\);
    
    \CLKPHASE_0_RNISVR71[3]\ : MX2
      port map(A => N_3760, B => N_3765, S => 
        \CLKPHASE_0[3]_net_1\, Y => N_3770);
    
    \RECD_SER_WORD_RNO_5[1]\ : NOR3C
      port map(A => n_recd_ser_word165_2, B => 
        n_recd_ser_word166_0, C => \ARB_BYTE[3]_net_1\, Y => 
        \ARB_BYTE_m_0[3]\);
    
    \REG40M.BIT_OS_CNT_6_RNIU7711[0]\ : OR2A
      port map(A => \BIT_OS_CNT_6[0]\, B => N_365, Y => N_378);
    
    \RECD_SER_WORD_RNO_8[6]\ : NOR3C
      port map(A => n_recd_ser_word165_2, B => 
        n_recd_ser_word167_1, C => \ARB_BYTE[9]_net_1\, Y => 
        \ARB_BYTE_m_3[9]\);
    
    un41_n_seqcnts_I_10 : AND3
      port map(A => \un39_n_seqcnts[0]\, B => \un39_n_seqcnts[1]\, 
        C => \un39_n_seqcnts[2]\, Y => \DWACT_FINC_E[0]\);
    
    \CLKPHASE_0_RNIMGRD2[2]\ : MX2
      port map(A => N_3638, B => N_3650, S => 
        \CLKPHASE_0[2]_net_1\, Y => N_3654);
    
    \BIT_OS_SEL_RNINMQF_0[1]\ : NOR2A
      port map(A => \BIT_OS_SEL[1]_net_1\, B => 
        \BIT_OS_SEL[0]_net_1\, Y => n_recd_ser_word166_0);
    
    \BEST_BIT_OS_VAL_RNO_3[3]\ : MX2
      port map(A => N_3889, B => N_3901, S => 
        \INDEX_CNT_0[2]_net_1\, Y => N_3905);
    
    \REG40M.SEQCNTS_18[2]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[2]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_8, E => N_310, Q => \SEQCNTS_18[2]\);
    
    \REG40M.SEQCNTS_10[3]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[3]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_18, E => N_326, Q => \SEQCNTS_10[3]\);
    
    \CLKPHASE_0_RNI69V31[3]\ : MX2
      port map(A => N_3673, B => N_3677, S => 
        \CLKPHASE_0[3]_net_1\, Y => N_3681);
    
    \RECD_SER_WORD_RNO_6[2]\ : OA1
      port map(A => \BIT_OS_SEL[3]_net_1\, B => 
        n_recd_ser_word164, C => \ARB_BYTE[2]_net_1\, Y => 
        \ARB_BYTE_m_1[2]\);
    
    \DES_SM_RNO_0[4]\ : NOR3C
      port map(A => N_5072_2, B => DES_SM_tr7_0, C => N_215, Y
         => N_5072);
    
    \BEST_CLKPHASE_RNO[1]\ : NOR2A
      port map(A => I_5_0, B => \DES_SM_1[8]_net_1\, Y => 
        \N_BEST_CLKPHASE[1]\);
    
    \CLKPHASE_0_RNI8OLNH7[2]\ : AO1
      port map(A => \un36_n_bit_os_val[21]\, B => N_782_0, C => 
        N_717_0, Y => N_326);
    
    \REG40M.SEQCNTS_22[1]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[1]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_5, E => N_302, Q => \SEQCNTS_22[1]\);
    
    \REG40M.SEQCNTS_16[3]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[3]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_5, E => N_314, Q => \SEQCNTS_16[3]\);
    
    \REG40M.BIT_OS_CNT_1[0]\ : DFN1E1C0
      port map(D => N_557, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_4, E => BIT_OS_CNT_1e, Q => 
        \BIT_OS_CNT_1[0]\);
    
    \TUNE_CLKPHASE[0]\ : DFN1E1P0
      port map(D => I0_un1_S, CLK => CLK_40M_GL, PRE => 
        P_MASTER_POR_B_c_12, E => \DES_SM[1]_net_1\, Q => 
        \TUNE_CLKPHASE[0]_net_1\);
    
    \REG40M.SEQCNTS_21[3]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[3]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_3, E => N_304, Q => \SEQCNTS_21[3]\);
    
    \DES_SM_3[6]\ : DFN1C0
      port map(D => N_MAX_CNT_0_sqmuxa, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_27_1, Q => \DES_SM_3[6]_net_1\);
    
    \RECD_SER_WORD_RNO_1[6]\ : AO1
      port map(A => \ARB_BYTE[10]_net_1\, B => n_recd_ser_word168, 
        C => \ARB_BYTE_m_1[11]\, Y => \N_RECD_SER_WORD_iv_0[6]\);
    
    \BEST_BIT_OS_VAL_RNO_13[1]\ : MX2
      port map(A => N_3963, B => N_3967, S => 
        \INDEX_CNT_1[3]_net_1\, Y => N_3971);
    
    \REG40M.BIT_OS_VAL_13_RNO[0]\ : MX2
      port map(A => \BIT_OS_VAL_13[0]\, B => N_5666, S => 
        \un36_n_bit_os_val[18]\, Y => N_261);
    
    \RECD_SER_WORD_RNO_2[0]\ : OR3
      port map(A => \ARB_BYTE_m[2]\, B => \ARB_BYTE_m[0]\, C => 
        \N_RECD_SER_WORD_iv_3[0]\, Y => \N_RECD_SER_WORD_iv_5[0]\);
    
    \REG40M.BIT_OS_VAL_2_RNI4EQR[3]\ : MX2
      port map(A => \BIT_OS_VAL_2[3]\, B => \BIT_OS_VAL_18[3]\, S
         => \CLKPHASE_1[4]_net_1\, Y => N_3690);
    
    \REG40M.BIT_OS_VAL_21_RNO[0]\ : MX2
      port map(A => \BIT_OS_VAL_21[0]\, B => N_5666, S => 
        \un36_n_bit_os_val[10]\, Y => N_240);
    
    \REG40M.SEQCNTS_25_RNI693Q[3]\ : MX2
      port map(A => \SEQCNTS_25[3]\, B => \SEQCNTS_26[3]\, S => 
        \INDEX_CNT_4[0]_net_1\, Y => N_4041);
    
    \REG40M.BIT_OS_CNT_1_RNO[3]\ : NOR3A
      port map(A => N_380, B => N_554, C => N_4530_1, Y => N_135);
    
    \TUNE_CLKPHASE_RNIDA643[2]\ : AO1A
      port map(A => N_5780, B => \TUNE_CLKPHASE[2]_net_1\, C => 
        N_5794, Y => \TUNE_CLKPHASE_RNIDA643[2]_net_1\);
    
    \REG40M.SEQCNTS_25_RNI253Q[1]\ : MX2
      port map(A => \SEQCNTS_25[1]\, B => \SEQCNTS_26[1]\, S => 
        \INDEX_CNT_4[0]_net_1\, Y => N_4039);
    
    \INDEX_CNT_1_RNI85VM1[3]\ : MX2
      port map(A => N_4033, B => N_4038, S => 
        \INDEX_CNT_1[3]_net_1\, Y => N_4043);
    
    \DES_SM_RNIGJIS[0]\ : NOR2A
      port map(A => N_123, B => \DES_SM[0]_net_1\, Y => 
        un1_DES_SM_471_i_0_0_0_a3_0);
    
    \REG40M.BIT_OS_CNT_4_RNO_0[6]\ : OA1C
      port map(A => \BIT_OS_CNT_4[5]\, B => N_382, C => 
        \BIT_OS_CNT_4[6]\, Y => N_501);
    
    \REG40M.SEQCNTS_13[2]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[2]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_1, E => N_320, Q => \SEQCNTS_13[2]\);
    
    \BEST_BIT_OS_VAL_RNO_7[1]\ : MX2
      port map(A => N_3879, B => N_3883, S => 
        \INDEX_CNT_0[3]_net_1\, Y => N_3887);
    
    \REG40M.BIT_OS_VAL_12[1]\ : DFN1E1C0
      port map(D => \N_BIT_OS_VAL_12_18[1]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_10, E => \DES_SM_1[6]_net_1\, Q
         => \BIT_OS_VAL_12[1]\);
    
    \RECD_SER_WORD_RNO_5[3]\ : NOR3C
      port map(A => n_recd_ser_word165_2, B => 
        n_recd_ser_word166_0, C => \ARB_BYTE[5]_net_1\, Y => 
        \ARB_BYTE_m_2[5]\);
    
    un41_n_seqcnts_I_8 : AND3
      port map(A => \un39_n_seqcnts[0]\, B => \un39_n_seqcnts[1]\, 
        C => \un39_n_seqcnts[2]\, Y => N_3_1);
    
    un1_CLKPHASE_I_20 : XOR2
      port map(A => \CLKPHASE[4]_net_1\, B => 
        \DWACT_ADD_CI_0_g_array_2[0]\, Y => I_20);
    
    \BIT_OS_SEL_2[1]\ : DFN1C0
      port map(D => \BEST_BIT_OS_VAL[1]_net_1\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_27_0, Q => BIT_OS_SEL_2(1));
    
    \BEST_BIT_OS_VAL_RNO_16[0]\ : MX2
      port map(A => \BIT_OS_VAL_9[0]\, B => \BIT_OS_VAL_10[0]\, S
         => \INDEX_CNT_0[0]_net_1\, Y => N_3882);
    
    \RECD_SER_WORD[5]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[5]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_30, Q => \RECD_SER_WORD[5]_net_1\);
    
    \CLKPHASE_RNIO61T9[0]\ : MX2
      port map(A => N_3795, B => N_3870, S => \CLKPHASE[0]_net_1\, 
        Y => \un39_n_seqcnts[2]\);
    
    \REG40M.SEQCNTS_23[1]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[1]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_6, E => N_300, Q => \SEQCNTS_23[1]\);
    
    \REG40M.BIT_OS_VAL_1_RNO[2]\ : MX2
      port map(A => N_781_0, B => \BIT_OS_VAL_1[2]\, S => N_5676, 
        Y => N_5654);
    
    \REG40M.BIT_OS_CNT_1[7]\ : DFN1E1C0
      port map(D => N_127, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_4, E => BIT_OS_CNT_1e, Q => 
        \BIT_OS_CNT_1[7]\);
    
    \REG40M.BIT_OS_CNT_0_RNO[5]\ : XA1C
      port map(A => \BIT_OS_CNT_0[5]\, B => N_383, C => N_4530_2, 
        Y => N_113);
    
    \BIT_OS_SEL_4[1]\ : DFN1C0
      port map(D => \BEST_BIT_OS_VAL[1]_net_1\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_27_0, Q => BIT_OS_SEL_4(1));
    
    \ARB_BYTE_RNIFBTD1[0]\ : NOR3C
      port map(A => BIT_OS_CNT_3lde_0_a3_1, B => 
        BIT_OS_CNT_3lde_0_a3_0, C => N_776, Y => 
        BIT_OS_CNT_3lde_0_a3_3);
    
    \CLKPHASE_1[4]\ : DFN1C0
      port map(D => \TUNE_CLKPHASE_RNITINS2[4]_net_1\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_24_0, Q => 
        \CLKPHASE_1[4]_net_1\);
    
    \REG40M.BIT_OS_CNT_6_RNO[7]\ : NOR3A
      port map(A => N_419, B => N_4530_2, C => 
        BIT_OS_CNT_6_n7_i_0, Y => N_73);
    
    \REG40M.SEQCNTS_21[1]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[1]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_3, E => N_304, Q => \SEQCNTS_21[1]\);
    
    \REG40M.BIT_OS_CNT_3[5]\ : DFN1E1C0
      port map(D => BIT_OS_CNT_3_n5, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_7, E => BIT_OS_CNT_3e, Q => 
        \BIT_OS_CNT_3[5]\);
    
    \RECD_SER_WORD_RNIJJBK_0[6]\ : NOR2A
      port map(A => \RECD_SER_WORD[6]_net_1\, B => DCB_SALT_SEL_c, 
        Y => TFC_RX_SER_WORD(6));
    
    \REG40M.SEQCNTS_27[3]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1[3]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_13, E => N_292, Q => \SEQCNTS_27[3]\);
    
    \REG40M.BIT_OS_VAL_10_RNO[0]\ : MX2
      port map(A => \BIT_OS_VAL_10[0]\, B => N_5666, S => 
        \un36_n_bit_os_val[21]\, Y => N_270);
    
    \CLKPHASE_RNI7L0A5[1]\ : MX2
      port map(A => N_3831, B => N_3866, S => \CLKPHASE[1]_net_1\, 
        Y => N_3871);
    
    \CLKPHASE[4]\ : DFN1C0
      port map(D => \TUNE_CLKPHASE_RNITINS2[4]_net_1\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_24_0, Q => 
        \CLKPHASE[4]_net_1\);
    
    \WAITCNT[3]\ : DFN1E0C0
      port map(D => N_39, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_9, E => N_5790, Q => \WAITCNT[3]_net_1\);
    
    \REG40M.SEQCNTS_20_RNITOMJ[0]\ : MX2
      port map(A => \SEQCNTS_19[0]\, B => \SEQCNTS_20[0]\, S => 
        \INDEX_CNT_4[0]_net_1\, Y => N_4103);
    
    \REG40M.SEQCNTS_25_RNI8B3Q[4]\ : MX2
      port map(A => \SEQCNTS_25[4]\, B => \SEQCNTS_26[4]\, S => 
        \INDEX_CNT_4[0]_net_1\, Y => N_4042);
    
    \REG40M.BIT_OS_VAL_8_RNO[3]\ : MX2
      port map(A => \BIT_OS_VAL_8[3]\, B => N_209_0, S => 
        \un36_n_bit_os_val[23]\, Y => \N_BIT_OS_VAL_8_18[3]\);
    
    \CLKPHASE_0_RNIDPFH4[1]\ : MX2
      port map(A => N_3755, B => N_3790, S => 
        \CLKPHASE_0[1]_net_1\, Y => N_3795);
    
    \REG40M.SEQCNTS_31[0]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[0]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_9, E => N_284, Q => \SEQCNTS_31[0]\);
    
    \REG40M.SEQCNTS_23[0]\ : DFN1E1C0
      port map(D => \N_SEQCNTS_1_0[0]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_6, E => N_300, Q => \SEQCNTS_23[0]\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity TOP_MASTER_DES320M is

    port( BIT_OS_SEL_7_0        : out   std_logic;
          BIT_OS_SEL_6          : out   std_logic_vector(2 downto 1);
          BIT_OS_SEL_5          : out   std_logic_vector(2 downto 0);
          BIT_OS_SEL_4          : out   std_logic_vector(2 downto 0);
          BIT_OS_SEL_3          : out   std_logic_vector(2 downto 0);
          BIT_OS_SEL_2          : out   std_logic_vector(2 downto 0);
          BIT_OS_SEL_1          : out   std_logic_vector(2 downto 0);
          BIT_OS_SEL_0          : out   std_logic_vector(2 downto 0);
          OP_MODE_c_0           : in    std_logic;
          BIT_OS_SEL            : out   std_logic_vector(2 downto 0);
          TFC_RX_SER_WORD       : out   std_logic_vector(7 downto 0);
          ELK_RX_SER_WORD_0     : out   std_logic_vector(7 downto 0);
          P_MASTER_POR_B_c_27_0 : in    std_logic;
          P_MASTER_POR_B_c_27_1 : in    std_logic;
          P_MASTER_POR_B_c_16_0 : in    std_logic;
          P_MASTER_POR_B_c_17_0 : in    std_logic;
          P_MASTER_POR_B_c_24_0 : in    std_logic;
          TFC_SYNC_DET_1        : out   std_logic;
          ELK0_SYNC_DET_1       : out   std_logic;
          DCB_SALT_SEL_c        : in    std_logic;
          TFC_IN_R              : in    std_logic;
          ELK0_IN_R             : in    std_logic;
          TFC_IN_F              : in    std_logic;
          ELK0_IN_F             : in    std_logic;
          ALL_PLL_LOCK_c        : out   std_logic;
          CCC_MAIN_LOCK         : in    std_logic;
          P_MASTER_POR_B_c_31_0 : in    std_logic;
          P_MASTER_POR_B_c_26   : in    std_logic;
          P_MASTER_POR_B_c_32   : in    std_logic;
          P_MASTER_POR_B_c_24   : in    std_logic;
          P_MASTER_POR_B_c_5    : in    std_logic;
          P_MASTER_POR_B_c_4    : in    std_logic;
          P_MASTER_POR_B_c_2    : in    std_logic;
          P_MASTER_POR_B_c_3    : in    std_logic;
          P_MASTER_POR_B_c_9    : in    std_logic;
          P_MASTER_POR_B_c_21   : in    std_logic;
          P_MASTER_POR_B_c_15   : in    std_logic;
          P_MASTER_POR_B_c_16   : in    std_logic;
          P_MASTER_POR_B_c_12   : in    std_logic;
          P_MASTER_POR_B_c_11   : in    std_logic;
          P_MASTER_POR_B_c_7    : in    std_logic;
          ALIGN_ACTIVE          : out   std_logic;
          P_MASTER_POR_B_c_27   : in    std_logic;
          P_MASTER_POR_B_c_10   : in    std_logic;
          P_MASTER_POR_B_c_17   : in    std_logic;
          P_MASTER_POR_B_c_1    : in    std_logic;
          P_MASTER_POR_B_c_20   : in    std_logic;
          P_MASTER_POR_B_c_8    : in    std_logic;
          P_MASTER_POR_B_c_29   : in    std_logic;
          P_MASTER_POR_B_c_30   : in    std_logic;
          P_MASTER_POR_B_c_28   : in    std_logic;
          P_MASTER_POR_B_c_34_0 : in    std_logic;
          P_MASTER_POR_B_c_32_0 : in    std_logic;
          CCC_160M_FXD          : in    std_logic;
          P_MASTER_POR_B_c_23   : in    std_logic;
          P_MASTER_POR_B_c      : in    std_logic;
          CLK_40M_BUF_RECD      : in    std_logic;
          CLK_40M_GL            : in    std_logic;
          P_MASTER_POR_B_c_22_0 : in    std_logic;
          P_MASTER_POR_B_c_14   : in    std_logic;
          P_MASTER_POR_B_c_6    : in    std_logic;
          P_MASTER_POR_B_c_25   : in    std_logic;
          P_MASTER_POR_B_c_13   : in    std_logic;
          P_MASTER_POR_B_c_22   : in    std_logic;
          P_MASTER_POR_B_c_31   : in    std_logic;
          P_MASTER_POR_B_c_33   : in    std_logic;
          P_MASTER_POR_B_c_18   : in    std_logic;
          P_MASTER_POR_B_c_19   : in    std_logic;
          P_MASTER_POR_B_c_34   : in    std_logic;
          CCC_160M_ADJ          : out   std_logic
        );

end TOP_MASTER_DES320M;

architecture DEF_ARCH of TOP_MASTER_DES320M is 

  component CCC_DYN_TRIPLE_160M
    port( AUX_SUPDATE      : in    std_logic := 'U';
          AUX_SSHIFT       : in    std_logic := 'U';
          AUX_SDIN         : in    std_logic := 'U';
          AUX_MODE         : in    std_logic := 'U';
          CCC_RX_CLK_LOCK  : out   std_logic;
          CCC_160M_2ADJ_1  : out   std_logic;
          CCC_160M_1ADJ_1  : out   std_logic;
          CCC_160M_ADJ_1   : out   std_logic;
          CLK_40M_BUF_RECD : in    std_logic := 'U';
          CLK_40M_GL       : in    std_logic := 'U'
        );
  end component;

  component GP_CCC_SCONFIG
    port( PHASE_ADJ_160_L       : in    std_logic_vector(4 downto 0) := (others => 'U');
          P_MASTER_POR_B_c_34   : in    std_logic := 'U';
          P_MASTER_POR_B_c_19   : in    std_logic := 'U';
          P_MASTER_POR_B_c_18   : in    std_logic := 'U';
          P_MASTER_POR_B_c_33   : in    std_logic := 'U';
          P_MASTER_POR_B_c_31   : in    std_logic := 'U';
          P_MASTER_POR_B_c_22   : in    std_logic := 'U';
          AUX_SSHIFT            : out   std_logic;
          P_MASTER_POR_B_c_13   : in    std_logic := 'U';
          AUX_SUPDATE           : out   std_logic;
          P_MASTER_POR_B_c_25   : in    std_logic := 'U';
          P_MASTER_POR_B_c_6    : in    std_logic := 'U';
          AUX_SDIN              : out   std_logic;
          P_MASTER_POR_B_c_14   : in    std_logic := 'U';
          CCC2_CONFIG_TRIG_i_0  : in    std_logic := 'U';
          AUX_MODE              : out   std_logic;
          P_MASTER_POR_B_c_22_0 : in    std_logic := 'U';
          CLK_40M_GL            : in    std_logic := 'U'
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component MASTER_DES320M
    port( PHASE_ADJ_160_L       : out   std_logic_vector(4 downto 0);
          ELK_RX_SER_WORD_0     : out   std_logic_vector(7 downto 0);
          TFC_RX_SER_WORD       : out   std_logic_vector(7 downto 0);
          BIT_OS_SEL            : out   std_logic_vector(2 downto 0);
          OP_MODE_c_0           : in    std_logic := 'U';
          BIT_OS_SEL_0          : out   std_logic_vector(2 downto 0);
          BIT_OS_SEL_1          : out   std_logic_vector(2 downto 0);
          BIT_OS_SEL_2          : out   std_logic_vector(2 downto 0);
          BIT_OS_SEL_3          : out   std_logic_vector(2 downto 0);
          BIT_OS_SEL_4          : out   std_logic_vector(2 downto 0);
          BIT_OS_SEL_5          : out   std_logic_vector(2 downto 0);
          BIT_OS_SEL_6          : out   std_logic_vector(2 downto 1);
          BIT_OS_SEL_7_0        : out   std_logic;
          P_MASTER_POR_B_c      : in    std_logic := 'U';
          P_MASTER_POR_B_c_23   : in    std_logic := 'U';
          P_MASTER_POR_B_c_34   : in    std_logic := 'U';
          CCC_160M_FXD          : in    std_logic := 'U';
          P_MASTER_POR_B_c_33   : in    std_logic := 'U';
          P_MASTER_POR_B_c_32_0 : in    std_logic := 'U';
          P_MASTER_POR_B_c_34_0 : in    std_logic := 'U';
          P_MASTER_POR_B_c_28   : in    std_logic := 'U';
          P_MASTER_POR_B_c_30   : in    std_logic := 'U';
          P_MASTER_POR_B_c_29   : in    std_logic := 'U';
          P_MASTER_POR_B_c_8    : in    std_logic := 'U';
          P_MASTER_POR_B_c_19   : in    std_logic := 'U';
          P_MASTER_POR_B_c_18   : in    std_logic := 'U';
          P_MASTER_POR_B_c_20   : in    std_logic := 'U';
          P_MASTER_POR_B_c_1    : in    std_logic := 'U';
          P_MASTER_POR_B_c_17   : in    std_logic := 'U';
          P_MASTER_POR_B_c_13   : in    std_logic := 'U';
          P_MASTER_POR_B_c_10   : in    std_logic := 'U';
          P_MASTER_POR_B_c_27   : in    std_logic := 'U';
          ALIGN_ACTIVE          : out   std_logic;
          P_MASTER_POR_B_c_7    : in    std_logic := 'U';
          P_MASTER_POR_B_c_11   : in    std_logic := 'U';
          P_MASTER_POR_B_c_12   : in    std_logic := 'U';
          P_MASTER_POR_B_c_14   : in    std_logic := 'U';
          P_MASTER_POR_B_c_16   : in    std_logic := 'U';
          P_MASTER_POR_B_c_15   : in    std_logic := 'U';
          P_MASTER_POR_B_c_21   : in    std_logic := 'U';
          P_MASTER_POR_B_c_9    : in    std_logic := 'U';
          P_MASTER_POR_B_c_3    : in    std_logic := 'U';
          P_MASTER_POR_B_c_2    : in    std_logic := 'U';
          P_MASTER_POR_B_c_4    : in    std_logic := 'U';
          P_MASTER_POR_B_c_6    : in    std_logic := 'U';
          P_MASTER_POR_B_c_5    : in    std_logic := 'U';
          P_MASTER_POR_B_c_24   : in    std_logic := 'U';
          CCC2_CONFIG_TRIG_i_0  : out   std_logic;
          P_MASTER_POR_B_c_32   : in    std_logic := 'U';
          P_MASTER_POR_B_c_26   : in    std_logic := 'U';
          P_MASTER_POR_B_c_31_0 : in    std_logic := 'U';
          CCC_160M_ADJ          : in    std_logic := 'U';
          CCC_MAIN_LOCK         : in    std_logic := 'U';
          ALL_PLL_LOCK_c        : out   std_logic;
          ELK0_IN_F             : in    std_logic := 'U';
          TFC_IN_F              : in    std_logic := 'U';
          ELK0_IN_R             : in    std_logic := 'U';
          TFC_IN_R              : in    std_logic := 'U';
          DCB_SALT_SEL_c        : in    std_logic := 'U';
          ELK0_SYNC_DET_1       : out   std_logic;
          TFC_SYNC_DET_1        : out   std_logic;
          CCC_RX_CLK_LOCK       : in    std_logic := 'U';
          P_MASTER_POR_B_c_24_0 : in    std_logic := 'U';
          P_MASTER_POR_B_c_17_0 : in    std_logic := 'U';
          P_MASTER_POR_B_c_16_0 : in    std_logic := 'U';
          P_MASTER_POR_B_c_27_1 : in    std_logic := 'U';
          P_MASTER_POR_B_c_27_0 : in    std_logic := 'U';
          CLK_40M_GL            : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal CCC_160M_2ADJ, CCC_160M_1ADJ, \CCC_160M_ADJ\, 
        \PHASE_ADJ_160_L[0]\, \PHASE_ADJ_160_L[1]\, 
        \PHASE_ADJ_160_L[2]\, \PHASE_ADJ_160_L[3]\, 
        \PHASE_ADJ_160_L[4]\, AUX_SSHIFT, AUX_SUPDATE, AUX_SDIN, 
        CCC2_CONFIG_TRIG_i_0, AUX_MODE, CCC_RX_CLK_LOCK, \GND\, 
        \VCC\ : std_logic;

    for all : CCC_DYN_TRIPLE_160M
	Use entity work.CCC_DYN_TRIPLE_160M(DEF_ARCH);
    for all : GP_CCC_SCONFIG
	Use entity work.GP_CCC_SCONFIG(DEF_ARCH);
    for all : MASTER_DES320M
	Use entity work.MASTER_DES320M(DEF_ARCH);
begin 

    CCC_160M_ADJ <= \CCC_160M_ADJ\;

    U13B_CCC : CCC_DYN_TRIPLE_160M
      port map(AUX_SUPDATE => AUX_SUPDATE, AUX_SSHIFT => 
        AUX_SSHIFT, AUX_SDIN => AUX_SDIN, AUX_MODE => AUX_MODE, 
        CCC_RX_CLK_LOCK => CCC_RX_CLK_LOCK, CCC_160M_2ADJ_1 => 
        CCC_160M_2ADJ, CCC_160M_1ADJ_1 => CCC_160M_1ADJ, 
        CCC_160M_ADJ_1 => \CCC_160M_ADJ\, CLK_40M_BUF_RECD => 
        CLK_40M_BUF_RECD, CLK_40M_GL => CLK_40M_GL);
    
    U13A_ADJ_160M : GP_CCC_SCONFIG
      port map(PHASE_ADJ_160_L(4) => \PHASE_ADJ_160_L[4]\, 
        PHASE_ADJ_160_L(3) => \PHASE_ADJ_160_L[3]\, 
        PHASE_ADJ_160_L(2) => \PHASE_ADJ_160_L[2]\, 
        PHASE_ADJ_160_L(1) => \PHASE_ADJ_160_L[1]\, 
        PHASE_ADJ_160_L(0) => \PHASE_ADJ_160_L[0]\, 
        P_MASTER_POR_B_c_34 => P_MASTER_POR_B_c_34, 
        P_MASTER_POR_B_c_19 => P_MASTER_POR_B_c_19, 
        P_MASTER_POR_B_c_18 => P_MASTER_POR_B_c_18, 
        P_MASTER_POR_B_c_33 => P_MASTER_POR_B_c_33, 
        P_MASTER_POR_B_c_31 => P_MASTER_POR_B_c_31, 
        P_MASTER_POR_B_c_22 => P_MASTER_POR_B_c_22, AUX_SSHIFT
         => AUX_SSHIFT, P_MASTER_POR_B_c_13 => 
        P_MASTER_POR_B_c_13, AUX_SUPDATE => AUX_SUPDATE, 
        P_MASTER_POR_B_c_25 => P_MASTER_POR_B_c_25, 
        P_MASTER_POR_B_c_6 => P_MASTER_POR_B_c_6, AUX_SDIN => 
        AUX_SDIN, P_MASTER_POR_B_c_14 => P_MASTER_POR_B_c_14, 
        CCC2_CONFIG_TRIG_i_0 => CCC2_CONFIG_TRIG_i_0, AUX_MODE
         => AUX_MODE, P_MASTER_POR_B_c_22_0 => 
        P_MASTER_POR_B_c_22_0, CLK_40M_GL => CLK_40M_GL);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    U13C_MASTER_DESER : MASTER_DES320M
      port map(PHASE_ADJ_160_L(4) => \PHASE_ADJ_160_L[4]\, 
        PHASE_ADJ_160_L(3) => \PHASE_ADJ_160_L[3]\, 
        PHASE_ADJ_160_L(2) => \PHASE_ADJ_160_L[2]\, 
        PHASE_ADJ_160_L(1) => \PHASE_ADJ_160_L[1]\, 
        PHASE_ADJ_160_L(0) => \PHASE_ADJ_160_L[0]\, 
        ELK_RX_SER_WORD_0(7) => ELK_RX_SER_WORD_0(7), 
        ELK_RX_SER_WORD_0(6) => ELK_RX_SER_WORD_0(6), 
        ELK_RX_SER_WORD_0(5) => ELK_RX_SER_WORD_0(5), 
        ELK_RX_SER_WORD_0(4) => ELK_RX_SER_WORD_0(4), 
        ELK_RX_SER_WORD_0(3) => ELK_RX_SER_WORD_0(3), 
        ELK_RX_SER_WORD_0(2) => ELK_RX_SER_WORD_0(2), 
        ELK_RX_SER_WORD_0(1) => ELK_RX_SER_WORD_0(1), 
        ELK_RX_SER_WORD_0(0) => ELK_RX_SER_WORD_0(0), 
        TFC_RX_SER_WORD(7) => TFC_RX_SER_WORD(7), 
        TFC_RX_SER_WORD(6) => TFC_RX_SER_WORD(6), 
        TFC_RX_SER_WORD(5) => TFC_RX_SER_WORD(5), 
        TFC_RX_SER_WORD(4) => TFC_RX_SER_WORD(4), 
        TFC_RX_SER_WORD(3) => TFC_RX_SER_WORD(3), 
        TFC_RX_SER_WORD(2) => TFC_RX_SER_WORD(2), 
        TFC_RX_SER_WORD(1) => TFC_RX_SER_WORD(1), 
        TFC_RX_SER_WORD(0) => TFC_RX_SER_WORD(0), BIT_OS_SEL(2)
         => BIT_OS_SEL(2), BIT_OS_SEL(1) => BIT_OS_SEL(1), 
        BIT_OS_SEL(0) => BIT_OS_SEL(0), OP_MODE_c_0 => 
        OP_MODE_c_0, BIT_OS_SEL_0(2) => BIT_OS_SEL_0(2), 
        BIT_OS_SEL_0(1) => BIT_OS_SEL_0(1), BIT_OS_SEL_0(0) => 
        BIT_OS_SEL_0(0), BIT_OS_SEL_1(2) => BIT_OS_SEL_1(2), 
        BIT_OS_SEL_1(1) => BIT_OS_SEL_1(1), BIT_OS_SEL_1(0) => 
        BIT_OS_SEL_1(0), BIT_OS_SEL_2(2) => BIT_OS_SEL_2(2), 
        BIT_OS_SEL_2(1) => BIT_OS_SEL_2(1), BIT_OS_SEL_2(0) => 
        BIT_OS_SEL_2(0), BIT_OS_SEL_3(2) => BIT_OS_SEL_3(2), 
        BIT_OS_SEL_3(1) => BIT_OS_SEL_3(1), BIT_OS_SEL_3(0) => 
        BIT_OS_SEL_3(0), BIT_OS_SEL_4(2) => BIT_OS_SEL_4(2), 
        BIT_OS_SEL_4(1) => BIT_OS_SEL_4(1), BIT_OS_SEL_4(0) => 
        BIT_OS_SEL_4(0), BIT_OS_SEL_5(2) => BIT_OS_SEL_5(2), 
        BIT_OS_SEL_5(1) => BIT_OS_SEL_5(1), BIT_OS_SEL_5(0) => 
        BIT_OS_SEL_5(0), BIT_OS_SEL_6(2) => BIT_OS_SEL_6(2), 
        BIT_OS_SEL_6(1) => BIT_OS_SEL_6(1), BIT_OS_SEL_7_0 => 
        BIT_OS_SEL_7_0, P_MASTER_POR_B_c => P_MASTER_POR_B_c, 
        P_MASTER_POR_B_c_23 => P_MASTER_POR_B_c_23, 
        P_MASTER_POR_B_c_34 => P_MASTER_POR_B_c_34, CCC_160M_FXD
         => CCC_160M_FXD, P_MASTER_POR_B_c_33 => 
        P_MASTER_POR_B_c_33, P_MASTER_POR_B_c_32_0 => 
        P_MASTER_POR_B_c_32_0, P_MASTER_POR_B_c_34_0 => 
        P_MASTER_POR_B_c_34_0, P_MASTER_POR_B_c_28 => 
        P_MASTER_POR_B_c_28, P_MASTER_POR_B_c_30 => 
        P_MASTER_POR_B_c_30, P_MASTER_POR_B_c_29 => 
        P_MASTER_POR_B_c_29, P_MASTER_POR_B_c_8 => 
        P_MASTER_POR_B_c_8, P_MASTER_POR_B_c_19 => 
        P_MASTER_POR_B_c_19, P_MASTER_POR_B_c_18 => 
        P_MASTER_POR_B_c_18, P_MASTER_POR_B_c_20 => 
        P_MASTER_POR_B_c_20, P_MASTER_POR_B_c_1 => 
        P_MASTER_POR_B_c_1, P_MASTER_POR_B_c_17 => 
        P_MASTER_POR_B_c_17, P_MASTER_POR_B_c_13 => 
        P_MASTER_POR_B_c_13, P_MASTER_POR_B_c_10 => 
        P_MASTER_POR_B_c_10, P_MASTER_POR_B_c_27 => 
        P_MASTER_POR_B_c_27, ALIGN_ACTIVE => ALIGN_ACTIVE, 
        P_MASTER_POR_B_c_7 => P_MASTER_POR_B_c_7, 
        P_MASTER_POR_B_c_11 => P_MASTER_POR_B_c_11, 
        P_MASTER_POR_B_c_12 => P_MASTER_POR_B_c_12, 
        P_MASTER_POR_B_c_14 => P_MASTER_POR_B_c_14, 
        P_MASTER_POR_B_c_16 => P_MASTER_POR_B_c_16, 
        P_MASTER_POR_B_c_15 => P_MASTER_POR_B_c_15, 
        P_MASTER_POR_B_c_21 => P_MASTER_POR_B_c_21, 
        P_MASTER_POR_B_c_9 => P_MASTER_POR_B_c_9, 
        P_MASTER_POR_B_c_3 => P_MASTER_POR_B_c_3, 
        P_MASTER_POR_B_c_2 => P_MASTER_POR_B_c_2, 
        P_MASTER_POR_B_c_4 => P_MASTER_POR_B_c_4, 
        P_MASTER_POR_B_c_6 => P_MASTER_POR_B_c_6, 
        P_MASTER_POR_B_c_5 => P_MASTER_POR_B_c_5, 
        P_MASTER_POR_B_c_24 => P_MASTER_POR_B_c_24, 
        CCC2_CONFIG_TRIG_i_0 => CCC2_CONFIG_TRIG_i_0, 
        P_MASTER_POR_B_c_32 => P_MASTER_POR_B_c_32, 
        P_MASTER_POR_B_c_26 => P_MASTER_POR_B_c_26, 
        P_MASTER_POR_B_c_31_0 => P_MASTER_POR_B_c_31_0, 
        CCC_160M_ADJ => \CCC_160M_ADJ\, CCC_MAIN_LOCK => 
        CCC_MAIN_LOCK, ALL_PLL_LOCK_c => ALL_PLL_LOCK_c, 
        ELK0_IN_F => ELK0_IN_F, TFC_IN_F => TFC_IN_F, ELK0_IN_R
         => ELK0_IN_R, TFC_IN_R => TFC_IN_R, DCB_SALT_SEL_c => 
        DCB_SALT_SEL_c, ELK0_SYNC_DET_1 => ELK0_SYNC_DET_1, 
        TFC_SYNC_DET_1 => TFC_SYNC_DET_1, CCC_RX_CLK_LOCK => 
        CCC_RX_CLK_LOCK, P_MASTER_POR_B_c_24_0 => 
        P_MASTER_POR_B_c_24_0, P_MASTER_POR_B_c_17_0 => 
        P_MASTER_POR_B_c_17_0, P_MASTER_POR_B_c_16_0 => 
        P_MASTER_POR_B_c_16_0, P_MASTER_POR_B_c_27_1 => 
        P_MASTER_POR_B_c_27_1, P_MASTER_POR_B_c_27_0 => 
        P_MASTER_POR_B_c_27_0, CLK_40M_GL => CLK_40M_GL);
    
    GND_i : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SLAVE_DES320S_1_17_14 is

    port( ELK_RX_SER_WORD_16     : out   std_logic_vector(7 downto 0);
          BIT_OS_SEL_3           : in    std_logic_vector(2 downto 0);
          BIT_OS_SEL_2_0         : in    std_logic;
          BIT_OS_SEL_1           : in    std_logic_vector(2 downto 1);
          CLK_40M_GL             : in    std_logic;
          CCC_160M_FXD           : in    std_logic;
          ELK_IN_R               : in    std_logic;
          ELK_IN_F               : in    std_logic;
          MASTER_DCB_POR_B_i_0_i : in    std_logic;
          CCC_160M_ADJ           : in    std_logic
        );

end SLAVE_DES320S_1_17_14;

architecture DEF_ARCH of SLAVE_DES320S_1_17_14 is 

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal N_17, \ARB_BYTE[0]_net_1\, \ARB_BYTE[4]_net_1\, N_18, 
        \ARB_BYTE[1]_net_1\, \ARB_BYTE[5]_net_1\, N_19, 
        \ARB_BYTE[2]_net_1\, \ARB_BYTE[6]_net_1\, N_20, 
        \ARB_BYTE[3]_net_1\, \ARB_BYTE[7]_net_1\, N_21, 
        \ARB_BYTE[8]_net_1\, N_22, \ARB_BYTE[9]_net_1\, N_23, 
        \ARB_BYTE[10]_net_1\, N_24, \ARB_BYTE[11]_net_1\, N_31, 
        \ARB_BYTE[12]_net_1\, N_32, \ARB_BYTE[13]_net_1\, N_33, 
        N_34, N_35, N_36, N_37, N_38, N_39, N_40, N_56, 
        \ARB_BYTE[14]_net_1\, N_64, \N_RECD_SER_WORD[0]\, 
        \N_RECD_SER_WORD[1]\, \N_RECD_SER_WORD[2]\, 
        \N_RECD_SER_WORD[3]\, \N_RECD_SER_WORD[4]\, 
        \N_RECD_SER_WORD[5]\, \N_RECD_SER_WORD[6]\, 
        \N_RECD_SER_WORD[7]\, \ADJ_SER_IN_F_0DEL\, 
        \ADJ_SER_IN_R_0DEL\, \ADJ_SER_IN_F_1DEL\, 
        \ADJ_SER_IN_R_1DEL\, \Q[0]_net_1\, \ADJ_Q[0]_net_1\, 
        \Q[1]_net_1\, \ADJ_Q[1]_net_1\, \Q[2]_net_1\, 
        \ADJ_Q[2]_net_1\, \Q[3]_net_1\, \ADJ_Q[3]_net_1\, 
        \Q[4]_net_1\, \ADJ_Q[4]_net_1\, \Q[5]_net_1\, 
        \ADJ_Q[5]_net_1\, \Q[6]_net_1\, \ADJ_Q[6]_net_1\, 
        \Q[7]_net_1\, \ADJ_Q[7]_net_1\, \Q[8]_net_1\, 
        \ADJ_Q[8]_net_1\, \Q[9]_net_1\, \ADJ_Q[9]_net_1\, 
        \Q[10]_net_1\, \ADJ_Q[10]_net_1\, \Q[11]_net_1\, 
        \ADJ_Q[11]_net_1\, \Q[12]_net_1\, \ADJ_Q[12]_net_1\, 
        \Q[13]_net_1\, \ADJ_Q[13]_net_1\, \Q[14]_net_1\, 
        \ADJ_Q[14]_net_1\, \ARB_WRD_40M_FIXED[0]_net_1\, 
        \ARB_WRD_40M_FIXED[1]_net_1\, 
        \ARB_WRD_40M_FIXED[2]_net_1\, 
        \ARB_WRD_40M_FIXED[3]_net_1\, 
        \ARB_WRD_40M_FIXED[4]_net_1\, 
        \ARB_WRD_40M_FIXED[5]_net_1\, 
        \ARB_WRD_40M_FIXED[6]_net_1\, 
        \ARB_WRD_40M_FIXED[7]_net_1\, 
        \ARB_WRD_40M_FIXED[8]_net_1\, 
        \ARB_WRD_40M_FIXED[9]_net_1\, 
        \ARB_WRD_40M_FIXED[10]_net_1\, 
        \ARB_WRD_40M_FIXED[11]_net_1\, 
        \ARB_WRD_40M_FIXED[12]_net_1\, 
        \ARB_WRD_40M_FIXED[13]_net_1\, 
        \ARB_WRD_40M_FIXED[14]_net_1\, \GND\, \VCC\ : std_logic;

begin 


    \RECD_SER_WORD_RNO[5]\ : MX2
      port map(A => N_38, B => N_39, S => BIT_OS_SEL_3(0), Y => 
        \N_RECD_SER_WORD[5]\);
    
    \ARB_WRD_40M_FIXED[9]\ : DFN1C0
      port map(D => \Q[9]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[9]_net_1\);
    
    \ADJ_Q[4]\ : DFN1C0
      port map(D => \ADJ_Q[2]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[4]_net_1\);
    
    \ARB_BYTE[6]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[6]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[6]_net_1\);
    
    ADJ_SER_IN_F_1DEL : DFN1C0
      port map(D => \ADJ_SER_IN_F_0DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_F_1DEL\);
    
    \ARB_BYTE_RNI97U91[4]\ : MX2
      port map(A => \ARB_BYTE[4]_net_1\, B => \ARB_BYTE[8]_net_1\, 
        S => BIT_OS_SEL_1(2), Y => N_21);
    
    \ARB_BYTE[0]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[0]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[0]_net_1\);
    
    \Q[11]\ : DFN1C0
      port map(D => \ADJ_Q[11]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[11]_net_1\);
    
    \ADJ_Q[8]\ : DFN1C0
      port map(D => \ADJ_Q[6]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[8]_net_1\);
    
    \ADJ_Q[6]\ : DFN1C0
      port map(D => \ADJ_Q[4]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[6]_net_1\);
    
    \ADJ_Q[12]\ : DFN1C0
      port map(D => \ADJ_Q[10]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[12]_net_1\);
    
    \RECD_SER_WORD_RNO_1[0]\ : MX2
      port map(A => \ARB_BYTE[0]_net_1\, B => \ARB_BYTE[4]_net_1\, 
        S => BIT_OS_SEL_1(2), Y => N_17);
    
    \Q[1]\ : DFN1C0
      port map(D => \ADJ_Q[1]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[1]_net_1\);
    
    \ARB_BYTE_RNI9CFT2[10]\ : MX2
      port map(A => N_21, B => N_23, S => BIT_OS_SEL_1(1), Y => 
        N_37);
    
    \ARB_BYTE_RNI31U91[1]\ : MX2
      port map(A => \ARB_BYTE[1]_net_1\, B => \ARB_BYTE[5]_net_1\, 
        S => BIT_OS_SEL_1(2), Y => N_18);
    
    \ARB_BYTE[4]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[4]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[4]_net_1\);
    
    \ADJ_Q[2]\ : DFN1C0
      port map(D => \ADJ_Q[0]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[2]_net_1\);
    
    \RECD_SER_WORD_RNO_1[7]\ : MX2
      port map(A => \ARB_BYTE[10]_net_1\, B => 
        \ARB_BYTE[14]_net_1\, S => BIT_OS_SEL_3(2), Y => N_56);
    
    \RECD_SER_WORD[4]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[4]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_16(4));
    
    \Q[5]\ : DFN1C0
      port map(D => \ADJ_Q[5]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[5]_net_1\);
    
    \ADJ_Q[11]\ : DFN1C0
      port map(D => \ADJ_Q[9]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[11]_net_1\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \ADJ_Q[3]\ : DFN1C0
      port map(D => \ADJ_Q[1]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[3]_net_1\);
    
    \Q[10]\ : DFN1C0
      port map(D => \ADJ_Q[10]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[10]_net_1\);
    
    \ARB_WRD_40M_FIXED[6]\ : DFN1C0
      port map(D => \Q[6]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[6]_net_1\);
    
    \ARB_WRD_40M_FIXED[1]\ : DFN1C0
      port map(D => \Q[1]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[1]_net_1\);
    
    \ARB_BYTE_RNIO3841[12]\ : MX2
      port map(A => \ARB_BYTE[8]_net_1\, B => 
        \ARB_BYTE[12]_net_1\, S => BIT_OS_SEL_1(2), Y => N_31);
    
    \RECD_SER_WORD[3]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[3]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_16(3));
    
    \ARB_BYTE_RNIDGFT2[11]\ : MX2
      port map(A => N_22, B => N_24, S => BIT_OS_SEL_1(1), Y => 
        N_38);
    
    \RECD_SER_WORD[0]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[0]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_16(0));
    
    \RECD_SER_WORD_RNO[3]\ : MX2
      port map(A => N_36, B => N_37, S => BIT_OS_SEL_3(0), Y => 
        \N_RECD_SER_WORD[3]\);
    
    \Q[0]\ : DFN1C0
      port map(D => \ADJ_Q[0]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[0]_net_1\);
    
    \ARB_BYTE_RNIM1841[11]\ : MX2
      port map(A => \ARB_BYTE[7]_net_1\, B => 
        \ARB_BYTE[11]_net_1\, S => BIT_OS_SEL_1(2), Y => N_24);
    
    \RECD_SER_WORD_RNO_0[7]\ : MX2
      port map(A => N_31, B => N_56, S => BIT_OS_SEL_3(1), Y => 
        N_64);
    
    \Q[7]\ : DFN1C0
      port map(D => \ADJ_Q[7]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[7]_net_1\);
    
    \ARB_BYTE[14]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[14]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[14]_net_1\);
    
    \ARB_WRD_40M_FIXED[2]\ : DFN1C0
      port map(D => \Q[2]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[2]_net_1\);
    
    \ARB_WRD_40M_FIXED[14]\ : DFN1C0
      port map(D => \Q[14]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[14]_net_1\);
    
    \RECD_SER_WORD_RNO[2]\ : MX2
      port map(A => N_35, B => N_36, S => BIT_OS_SEL_3(0), Y => 
        \N_RECD_SER_WORD[2]\);
    
    \ARB_BYTE_RNIMB533[1]\ : MX2
      port map(A => N_18, B => N_20, S => BIT_OS_SEL_1(1), Y => 
        N_34);
    
    \ARB_BYTE_RNIPBS82[10]\ : MX2
      port map(A => N_23, B => N_31, S => BIT_OS_SEL_2_0, Y => 
        N_39);
    
    \ARB_BYTE[2]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[2]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[2]_net_1\);
    
    \ARB_BYTE_RNIB9U91[5]\ : MX2
      port map(A => \ARB_BYTE[5]_net_1\, B => \ARB_BYTE[9]_net_1\, 
        S => BIT_OS_SEL_1(2), Y => N_22);
    
    \ADJ_Q[7]\ : DFN1C0
      port map(D => \ADJ_Q[5]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[7]_net_1\);
    
    \ARB_BYTE[8]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[8]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[8]_net_1\);
    
    \RECD_SER_WORD[5]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[5]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_16(5));
    
    \ARB_BYTE_RNIQ5841[13]\ : MX2
      port map(A => \ARB_BYTE[9]_net_1\, B => 
        \ARB_BYTE[13]_net_1\, S => BIT_OS_SEL_1(2), Y => N_32);
    
    \ARB_BYTE[12]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[12]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[12]_net_1\);
    
    \RECD_SER_WORD[1]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[1]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_16(1));
    
    \Q[3]\ : DFN1C0
      port map(D => \ADJ_Q[3]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[3]_net_1\);
    
    ADJ_SER_IN_F_0DEL : DFN1C0
      port map(D => ELK_IN_F, CLK => CCC_160M_ADJ, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_F_0DEL\);
    
    \RECD_SER_WORD_RNO[7]\ : MX2
      port map(A => N_40, B => N_64, S => BIT_OS_SEL_3(0), Y => 
        \N_RECD_SER_WORD[7]\);
    
    \RECD_SER_WORD_RNO[1]\ : MX2
      port map(A => N_34, B => N_35, S => BIT_OS_SEL_3(0), Y => 
        \N_RECD_SER_WORD[1]\);
    
    \ARB_WRD_40M_FIXED[4]\ : DFN1C0
      port map(D => \Q[4]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[4]_net_1\);
    
    \RECD_SER_WORD_RNO[0]\ : MX2
      port map(A => N_33, B => N_34, S => BIT_OS_SEL_3(0), Y => 
        \N_RECD_SER_WORD[0]\);
    
    \Q[6]\ : DFN1C0
      port map(D => \ADJ_Q[6]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[6]_net_1\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \ARB_WRD_40M_FIXED[8]\ : DFN1C0
      port map(D => \Q[8]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[8]_net_1\);
    
    \ARB_BYTE_RNIQF533[2]\ : MX2
      port map(A => N_19, B => N_21, S => BIT_OS_SEL_1(1), Y => 
        N_35);
    
    \ARB_BYTE[11]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[11]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[11]_net_1\);
    
    \Q[9]\ : DFN1C0
      port map(D => \ADJ_Q[9]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[9]_net_1\);
    
    \Q[14]\ : DFN1C0
      port map(D => \ADJ_Q[14]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[14]_net_1\);
    
    ADJ_SER_IN_R_0DEL : DFN1C0
      port map(D => ELK_IN_R, CLK => CCC_160M_ADJ, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_R_0DEL\);
    
    \Q[13]\ : DFN1C0
      port map(D => \ADJ_Q[13]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[13]_net_1\);
    
    \ARB_BYTE[9]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[9]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[9]_net_1\);
    
    ADJ_SER_IN_R_1DEL : DFN1C0
      port map(D => \ADJ_SER_IN_R_0DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_R_1DEL\);
    
    \ARB_BYTE[10]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[10]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[10]_net_1\);
    
    \ADJ_Q[9]\ : DFN1C0
      port map(D => \ADJ_Q[7]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[9]_net_1\);
    
    \RECD_SER_WORD[7]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[7]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_16(7));
    
    \ARB_WRD_40M_FIXED[5]\ : DFN1C0
      port map(D => \Q[5]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[5]_net_1\);
    
    \ARB_WRD_40M_FIXED[12]\ : DFN1C0
      port map(D => \Q[12]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[12]_net_1\);
    
    \ARB_WRD_40M_FIXED[11]\ : DFN1C0
      port map(D => \Q[11]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[11]_net_1\);
    
    \ARB_WRD_40M_FIXED[0]\ : DFN1C0
      port map(D => \Q[0]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[0]_net_1\);
    
    \ADJ_Q[10]\ : DFN1C0
      port map(D => \ADJ_Q[8]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[10]_net_1\);
    
    \Q[2]\ : DFN1C0
      port map(D => \ADJ_Q[2]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[2]_net_1\);
    
    \ARB_BYTE_RNI75U91[3]\ : MX2
      port map(A => \ARB_BYTE[3]_net_1\, B => \ARB_BYTE[7]_net_1\, 
        S => BIT_OS_SEL_1(2), Y => N_20);
    
    \ADJ_Q[1]\ : DFN1C0
      port map(D => \ADJ_SER_IN_F_1DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[1]_net_1\);
    
    \RECD_SER_WORD[6]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[6]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_16(6));
    
    \RECD_SER_WORD[2]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[2]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_16(2));
    
    \ADJ_Q[13]\ : DFN1C0
      port map(D => \ADJ_Q[11]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[13]_net_1\);
    
    \ARB_BYTE_RNITFS82[13]\ : MX2
      port map(A => N_24, B => N_32, S => BIT_OS_SEL_2_0, Y => 
        N_40);
    
    \ARB_BYTE_RNIKV741[10]\ : MX2
      port map(A => \ARB_BYTE[6]_net_1\, B => 
        \ARB_BYTE[10]_net_1\, S => BIT_OS_SEL_1(2), Y => N_23);
    
    \ARB_BYTE_RNI53U91[2]\ : MX2
      port map(A => \ARB_BYTE[2]_net_1\, B => \ARB_BYTE[6]_net_1\, 
        S => BIT_OS_SEL_1(2), Y => N_19);
    
    \Q[8]\ : DFN1C0
      port map(D => \ADJ_Q[8]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[8]_net_1\);
    
    \ARB_BYTE[5]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[5]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[5]_net_1\);
    
    \ADJ_Q[14]\ : DFN1C0
      port map(D => \ADJ_Q[12]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[14]_net_1\);
    
    \RECD_SER_WORD_RNO[4]\ : MX2
      port map(A => N_37, B => N_38, S => BIT_OS_SEL_3(0), Y => 
        \N_RECD_SER_WORD[4]\);
    
    \Q[12]\ : DFN1C0
      port map(D => \ADJ_Q[12]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[12]_net_1\);
    
    \ARB_BYTE[13]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[13]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[13]_net_1\);
    
    \ARB_WRD_40M_FIXED[3]\ : DFN1C0
      port map(D => \Q[3]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[3]_net_1\);
    
    \ARB_BYTE_RNIUJ533[3]\ : MX2
      port map(A => N_20, B => N_22, S => BIT_OS_SEL_1(1), Y => 
        N_36);
    
    \ARB_BYTE[7]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[7]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[7]_net_1\);
    
    \RECD_SER_WORD_RNO_0[0]\ : MX2
      port map(A => N_17, B => N_19, S => BIT_OS_SEL_1(1), Y => 
        N_33);
    
    \Q[4]\ : DFN1C0
      port map(D => \ADJ_Q[4]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[4]_net_1\);
    
    \ARB_WRD_40M_FIXED[7]\ : DFN1C0
      port map(D => \Q[7]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[7]_net_1\);
    
    \RECD_SER_WORD_RNO[6]\ : MX2
      port map(A => N_39, B => N_40, S => BIT_OS_SEL_3(0), Y => 
        \N_RECD_SER_WORD[6]\);
    
    \ARB_BYTE[3]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[3]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[3]_net_1\);
    
    \ADJ_Q[5]\ : DFN1C0
      port map(D => \ADJ_Q[3]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[5]_net_1\);
    
    \ARB_BYTE[1]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[1]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[1]_net_1\);
    
    \ARB_WRD_40M_FIXED[13]\ : DFN1C0
      port map(D => \Q[13]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[13]_net_1\);
    
    \ADJ_Q[0]\ : DFN1C0
      port map(D => \ADJ_SER_IN_R_1DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[0]_net_1\);
    
    \ARB_WRD_40M_FIXED[10]\ : DFN1C0
      port map(D => \Q[10]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[10]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SER320M_3_34_16 is

    port( ELK_TX_DAT                 : in    std_logic_vector(7 downto 0);
          MASTER_SALT_POR_B_i_0_i_14 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_10 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_0  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_16 : in    std_logic;
          ELK_OUT_R                  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_1  : in    std_logic;
          ELK_OUT_F                  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_8  : in    std_logic;
          CCC_160M_FXD               : in    std_logic;
          CLK_40M_GL                 : in    std_logic
        );

end SER320M_3_34_16;

architecture DEF_ARCH of SER320M_3_34_16 is 

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \N_SER_CMD_WORD_R[0]\, \START_RISE\, 
        \N_SER_CMD_WORD_F[0]\, \N_SER_CMD_WORD_R[3]\, 
        \SER_CMD_WORD_R[2]_net_1\, \N_SER_CMD_WORD_R[2]\, 
        \SER_CMD_WORD_R[1]_net_1\, \N_SER_CMD_WORD_R[1]\, 
        \SER_CMD_WORD_R[0]_net_1\, \N_SER_CMD_WORD_F[3]\, 
        \SER_CMD_WORD_F[2]_net_1\, \N_SER_CMD_WORD_F[2]\, 
        \SER_CMD_WORD_F[1]_net_1\, \N_SER_CMD_WORD_F[1]\, 
        \SER_CMD_WORD_F[0]_net_1\, N_START_RISE, 
        \CLK40M_GEN_DEL0\, \SER_OUT_FI\, \SER_OUT_RI\, 
        \SER_CMD_WORD_F[3]_net_1\, \SER_CMD_WORD_R[3]_net_1\, 
        \GND\, \VCC\ : std_logic;

begin 


    SER_OUT_FI : DFN1C0
      port map(D => \SER_CMD_WORD_F[3]_net_1\, CLK => 
        CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_10, Q => 
        \SER_OUT_FI\);
    
    \SER_CMD_WORD_F[3]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[3]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_14, Q => 
        \SER_CMD_WORD_F[3]_net_1\);
    
    \SER_CMD_WORD_R[1]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[1]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_10, Q => 
        \SER_CMD_WORD_R[1]_net_1\);
    
    \SER_CMD_WORD_R[2]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[2]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_10, Q => 
        \SER_CMD_WORD_R[2]_net_1\);
    
    \SER_CMD_WORD_R_RNO[3]\ : MX2
      port map(A => \SER_CMD_WORD_R[2]_net_1\, B => ELK_TX_DAT(7), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_R[3]\);
    
    \SER_CMD_WORD_R_RNO[0]\ : NOR2B
      port map(A => \START_RISE\, B => ELK_TX_DAT(1), Y => 
        \N_SER_CMD_WORD_R[0]\);
    
    \SER_CMD_WORD_F[0]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[0]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_14, Q => 
        \SER_CMD_WORD_F[0]_net_1\);
    
    \SER_CMD_WORD_R_RNO[1]\ : MX2
      port map(A => \SER_CMD_WORD_R[0]_net_1\, B => ELK_TX_DAT(3), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_R[1]\);
    
    \SER_CMD_WORD_F_RNO[2]\ : MX2
      port map(A => \SER_CMD_WORD_F[1]_net_1\, B => ELK_TX_DAT(4), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_F[2]\);
    
    \SER_CMD_WORD_F_RNO[3]\ : MX2
      port map(A => \SER_CMD_WORD_F[2]_net_1\, B => ELK_TX_DAT(6), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_F[3]\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    CLK40M_GEN_DEL0 : DFN1C0
      port map(D => CLK_40M_GL, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_8, Q => \CLK40M_GEN_DEL0\);
    
    SER_OUT_RI : DFN1C0
      port map(D => \SER_CMD_WORD_R[3]_net_1\, CLK => 
        CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_10, Q => 
        \SER_OUT_RI\);
    
    \SER_CMD_WORD_F[2]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[2]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_14, Q => 
        \SER_CMD_WORD_F[2]_net_1\);
    
    \SER_CMD_WORD_F_RNO[1]\ : MX2
      port map(A => \SER_CMD_WORD_F[0]_net_1\, B => ELK_TX_DAT(2), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_F[1]\);
    
    \SER_CMD_WORD_R[0]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[0]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_10, Q => 
        \SER_CMD_WORD_R[0]_net_1\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    START_RISE : DFN1C0
      port map(D => N_START_RISE, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_0, Q => \START_RISE\);
    
    \SER_CMD_WORD_R[3]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[3]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_10, Q => 
        \SER_CMD_WORD_R[3]_net_1\);
    
    \SER_CMD_WORD_F_RNO[0]\ : NOR2B
      port map(A => \START_RISE\, B => ELK_TX_DAT(0), Y => 
        \N_SER_CMD_WORD_F[0]\);
    
    SER_OUT_RDEL : DFN1C0
      port map(D => \SER_OUT_RI\, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_16, Q => ELK_OUT_R);
    
    \SER_CMD_WORD_F[1]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[1]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_14, Q => 
        \SER_CMD_WORD_F[1]_net_1\);
    
    START_RISE_RNO : NOR2B
      port map(A => \CLK40M_GEN_DEL0\, B => CLK_40M_GL, Y => 
        N_START_RISE);
    
    \SER_CMD_WORD_R_RNO[2]\ : MX2
      port map(A => \SER_CMD_WORD_R[1]_net_1\, B => ELK_TX_DAT(5), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_R[2]\);
    
    SER_OUT_FDEL : DFN1C0
      port map(D => \SER_OUT_FI\, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_1, Q => ELK_OUT_F);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity DDR_BIDIR_LVDS_DUAL_CLK_16 is

    port( DCB_SALT_SEL_c_i : in    std_logic;
          ELK16_DAT_P      : inout std_logic := 'Z';
          ELK16_DAT_N      : inout std_logic := 'Z';
          ELK_OUT_R        : in    std_logic;
          ELK_OUT_F        : in    std_logic;
          CCC_160M_FXD     : in    std_logic;
          CCC_160M_ADJ     : in    std_logic;
          ELK_IN_DDR_R     : out   std_logic;
          ELK_IN_DDR_F     : out   std_logic
        );

end DDR_BIDIR_LVDS_DUAL_CLK_16;

architecture DEF_ARCH of DDR_BIDIR_LVDS_DUAL_CLK_16 is 

  component DDR_REG
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          QR  : out   std_logic;
          QF  : out   std_logic
        );
  end component;

  component DDR_OUT
    port( DR  : in    std_logic := 'U';
          DF  : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component BIBUF_LVDS
    port( PADP : inout   std_logic;
          PADN : inout   std_logic;
          D    : in    std_logic := 'U';
          E    : in    std_logic := 'U';
          Y    : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal DDR_BIDIR_LVDS_DUAL_CLK_16_GND, BIBUF_LVDS_0_Y, 
        DDR_OUT_0_Q, \VCC\ : std_logic;

begin 


    DDR_REG_0 : DDR_REG
      port map(D => BIBUF_LVDS_0_Y, CLK => CCC_160M_ADJ, CLR => 
        DDR_BIDIR_LVDS_DUAL_CLK_16_GND, QR => ELK_IN_DDR_R, QF
         => ELK_IN_DDR_F);
    
    DDR_OUT_0 : DDR_OUT
      port map(DR => ELK_OUT_R, DF => ELK_OUT_F, CLK => 
        CCC_160M_FXD, CLR => DDR_BIDIR_LVDS_DUAL_CLK_16_GND, Q
         => DDR_OUT_0_Q);
    
    BIBUF_LVDS_0 : BIBUF_LVDS
      port map(PADP => ELK16_DAT_P, PADN => ELK16_DAT_N, D => 
        DDR_OUT_0_Q, E => DCB_SALT_SEL_c_i, Y => BIBUF_LVDS_0_Y);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    GND_i : GND
      port map(Y => DDR_BIDIR_LVDS_DUAL_CLK_16_GND);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SYNC_DAT_SEL_16 is

    port( ELK_TX_DAT                : out   std_logic_vector(7 downto 0);
          PATT_ELK_DAT_16           : in    std_logic_vector(7 downto 0);
          OP_MODE_c_2_0             : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_9 : in    std_logic;
          CLK_40M_GL                : in    std_logic
        );

end SYNC_DAT_SEL_16;

architecture DEF_ARCH of SYNC_DAT_SEL_16 is 

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \N_SERDAT[0]\, \N_SERDAT[1]\, \N_SERDAT[2]\, 
        \N_SERDAT[3]\, \N_SERDAT[4]\, \N_SERDAT[5]\, 
        \N_SERDAT[6]\, \N_SERDAT[7]\, \GND\, \VCC\ : std_logic;

begin 


    \SERDAT_RNO[4]\ : NOR2A
      port map(A => PATT_ELK_DAT_16(4), B => OP_MODE_c_2_0, Y => 
        \N_SERDAT[4]\);
    
    \SERDAT_RNO[0]\ : NOR2A
      port map(A => PATT_ELK_DAT_16(0), B => OP_MODE_c_2_0, Y => 
        \N_SERDAT[0]\);
    
    \SERDAT[6]\ : DFN1C0
      port map(D => \N_SERDAT[6]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_9, Q => ELK_TX_DAT(6));
    
    \SERDAT[4]\ : DFN1C0
      port map(D => \N_SERDAT[4]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_9, Q => ELK_TX_DAT(4));
    
    \SERDAT_RNO[7]\ : OR2
      port map(A => PATT_ELK_DAT_16(7), B => OP_MODE_c_2_0, Y => 
        \N_SERDAT[7]\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \SERDAT_RNO[3]\ : OR2
      port map(A => PATT_ELK_DAT_16(3), B => OP_MODE_c_2_0, Y => 
        \N_SERDAT[3]\);
    
    \SERDAT_RNO[2]\ : OR2
      port map(A => PATT_ELK_DAT_16(2), B => OP_MODE_c_2_0, Y => 
        \N_SERDAT[2]\);
    
    \SERDAT[5]\ : DFN1C0
      port map(D => \N_SERDAT[5]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_9, Q => ELK_TX_DAT(5));
    
    \SERDAT[7]\ : DFN1C0
      port map(D => \N_SERDAT[7]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_9, Q => ELK_TX_DAT(7));
    
    GND_i : GND
      port map(Y => \GND\);
    
    \SERDAT_RNO[5]\ : NOR2A
      port map(A => PATT_ELK_DAT_16(5), B => OP_MODE_c_2_0, Y => 
        \N_SERDAT[5]\);
    
    \SERDAT[0]\ : DFN1C0
      port map(D => \N_SERDAT[0]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_9, Q => ELK_TX_DAT(0));
    
    \SERDAT_RNO[6]\ : NOR2A
      port map(A => PATT_ELK_DAT_16(6), B => OP_MODE_c_2_0, Y => 
        \N_SERDAT[6]\);
    
    \SERDAT[1]\ : DFN1C0
      port map(D => \N_SERDAT[1]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_9, Q => ELK_TX_DAT(1));
    
    \SERDAT_RNO[1]\ : OR2
      port map(A => PATT_ELK_DAT_16(1), B => OP_MODE_c_2_0, Y => 
        \N_SERDAT[1]\);
    
    \SERDAT[3]\ : DFN1C0
      port map(D => \N_SERDAT[3]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_9, Q => ELK_TX_DAT(3));
    
    \SERDAT[2]\ : DFN1C0
      port map(D => \N_SERDAT[2]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_9, Q => ELK_TX_DAT(2));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity ELINK_SLAVE_15_11 is

    port( BIT_OS_SEL_1               : in    std_logic_vector(2 downto 1);
          BIT_OS_SEL_2_0             : in    std_logic;
          BIT_OS_SEL_3               : in    std_logic_vector(2 downto 0);
          ELK_RX_SER_WORD_16         : out   std_logic_vector(7 downto 0);
          OP_MODE_c_2_0              : in    std_logic;
          PATT_ELK_DAT_16            : in    std_logic_vector(7 downto 0);
          MASTER_DCB_POR_B_i_0_i     : in    std_logic;
          ELK16_DAT_N                : inout std_logic := 'Z';
          ELK16_DAT_P                : inout std_logic := 'Z';
          DCB_SALT_SEL_c_i           : in    std_logic;
          CCC_160M_FXD               : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_8  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_1  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_16 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_0  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_10 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_14 : in    std_logic;
          CLK_40M_GL                 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_9  : in    std_logic;
          DEV_RST_B_c_1              : in    std_logic;
          CCC_160M_ADJ               : in    std_logic
        );

end ELINK_SLAVE_15_11;

architecture DEF_ARCH of ELINK_SLAVE_15_11 is 

  component SLAVE_DES320S_1_17_14
    port( ELK_RX_SER_WORD_16     : out   std_logic_vector(7 downto 0);
          BIT_OS_SEL_3           : in    std_logic_vector(2 downto 0) := (others => 'U');
          BIT_OS_SEL_2_0         : in    std_logic := 'U';
          BIT_OS_SEL_1           : in    std_logic_vector(2 downto 1) := (others => 'U');
          CLK_40M_GL             : in    std_logic := 'U';
          CCC_160M_FXD           : in    std_logic := 'U';
          ELK_IN_R               : in    std_logic := 'U';
          ELK_IN_F               : in    std_logic := 'U';
          MASTER_DCB_POR_B_i_0_i : in    std_logic := 'U';
          CCC_160M_ADJ           : in    std_logic := 'U'
        );
  end component;

  component SER320M_3_34_16
    port( ELK_TX_DAT                 : in    std_logic_vector(7 downto 0) := (others => 'U');
          MASTER_SALT_POR_B_i_0_i_14 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_10 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_0  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_16 : in    std_logic := 'U';
          ELK_OUT_R                  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_1  : in    std_logic := 'U';
          ELK_OUT_F                  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_8  : in    std_logic := 'U';
          CCC_160M_FXD               : in    std_logic := 'U';
          CLK_40M_GL                 : in    std_logic := 'U'
        );
  end component;

  component DDR_BIDIR_LVDS_DUAL_CLK_16
    port( DCB_SALT_SEL_c_i : in    std_logic := 'U';
          ELK16_DAT_P      : inout   std_logic;
          ELK16_DAT_N      : inout   std_logic;
          ELK_OUT_R        : in    std_logic := 'U';
          ELK_OUT_F        : in    std_logic := 'U';
          CCC_160M_FXD     : in    std_logic := 'U';
          CCC_160M_ADJ     : in    std_logic := 'U';
          ELK_IN_DDR_R     : out   std_logic;
          ELK_IN_DDR_F     : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component SYNC_DAT_SEL_16
    port( ELK_TX_DAT                : out   std_logic_vector(7 downto 0);
          PATT_ELK_DAT_16           : in    std_logic_vector(7 downto 0) := (others => 'U');
          OP_MODE_c_2_0             : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_9 : in    std_logic := 'U';
          CLK_40M_GL                : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \ELK_IN_F\, ELK_IN_DDR_F, \ELK_IN_R\, ELK_IN_DDR_R, 
        \ELK_TX_DAT[0]\, \ELK_TX_DAT[1]\, \ELK_TX_DAT[2]\, 
        \ELK_TX_DAT[3]\, \ELK_TX_DAT[4]\, \ELK_TX_DAT[5]\, 
        \ELK_TX_DAT[6]\, \ELK_TX_DAT[7]\, ELK_OUT_R, ELK_OUT_F, 
        \GND\, \VCC\ : std_logic;

    for all : SLAVE_DES320S_1_17_14
	Use entity work.SLAVE_DES320S_1_17_14(DEF_ARCH);
    for all : SER320M_3_34_16
	Use entity work.SER320M_3_34_16(DEF_ARCH);
    for all : DDR_BIDIR_LVDS_DUAL_CLK_16
	Use entity work.DDR_BIDIR_LVDS_DUAL_CLK_16(DEF_ARCH);
    for all : SYNC_DAT_SEL_16
	Use entity work.SYNC_DAT_SEL_16(DEF_ARCH);
begin 


    U_SLAVE_1ELK : SLAVE_DES320S_1_17_14
      port map(ELK_RX_SER_WORD_16(7) => ELK_RX_SER_WORD_16(7), 
        ELK_RX_SER_WORD_16(6) => ELK_RX_SER_WORD_16(6), 
        ELK_RX_SER_WORD_16(5) => ELK_RX_SER_WORD_16(5), 
        ELK_RX_SER_WORD_16(4) => ELK_RX_SER_WORD_16(4), 
        ELK_RX_SER_WORD_16(3) => ELK_RX_SER_WORD_16(3), 
        ELK_RX_SER_WORD_16(2) => ELK_RX_SER_WORD_16(2), 
        ELK_RX_SER_WORD_16(1) => ELK_RX_SER_WORD_16(1), 
        ELK_RX_SER_WORD_16(0) => ELK_RX_SER_WORD_16(0), 
        BIT_OS_SEL_3(2) => BIT_OS_SEL_3(2), BIT_OS_SEL_3(1) => 
        BIT_OS_SEL_3(1), BIT_OS_SEL_3(0) => BIT_OS_SEL_3(0), 
        BIT_OS_SEL_2_0 => BIT_OS_SEL_2_0, BIT_OS_SEL_1(2) => 
        BIT_OS_SEL_1(2), BIT_OS_SEL_1(1) => BIT_OS_SEL_1(1), 
        CLK_40M_GL => CLK_40M_GL, CCC_160M_FXD => CCC_160M_FXD, 
        ELK_IN_R => \ELK_IN_R\, ELK_IN_F => \ELK_IN_F\, 
        MASTER_DCB_POR_B_i_0_i => MASTER_DCB_POR_B_i_0_i, 
        CCC_160M_ADJ => CCC_160M_ADJ);
    
    U_ELK1_CMD_TX : SER320M_3_34_16
      port map(ELK_TX_DAT(7) => \ELK_TX_DAT[7]\, ELK_TX_DAT(6)
         => \ELK_TX_DAT[6]\, ELK_TX_DAT(5) => \ELK_TX_DAT[5]\, 
        ELK_TX_DAT(4) => \ELK_TX_DAT[4]\, ELK_TX_DAT(3) => 
        \ELK_TX_DAT[3]\, ELK_TX_DAT(2) => \ELK_TX_DAT[2]\, 
        ELK_TX_DAT(1) => \ELK_TX_DAT[1]\, ELK_TX_DAT(0) => 
        \ELK_TX_DAT[0]\, MASTER_SALT_POR_B_i_0_i_14 => 
        MASTER_SALT_POR_B_i_0_i_14, MASTER_SALT_POR_B_i_0_i_10
         => MASTER_SALT_POR_B_i_0_i_10, MASTER_SALT_POR_B_i_0_i_0
         => MASTER_SALT_POR_B_i_0_i_0, MASTER_SALT_POR_B_i_0_i_16
         => MASTER_SALT_POR_B_i_0_i_16, ELK_OUT_R => ELK_OUT_R, 
        MASTER_SALT_POR_B_i_0_i_1 => MASTER_SALT_POR_B_i_0_i_1, 
        ELK_OUT_F => ELK_OUT_F, MASTER_SALT_POR_B_i_0_i_8 => 
        MASTER_SALT_POR_B_i_0_i_8, CCC_160M_FXD => CCC_160M_FXD, 
        CLK_40M_GL => CLK_40M_GL);
    
    U_DDR_ELK1 : DDR_BIDIR_LVDS_DUAL_CLK_16
      port map(DCB_SALT_SEL_c_i => DCB_SALT_SEL_c_i, ELK16_DAT_P
         => ELK16_DAT_P, ELK16_DAT_N => ELK16_DAT_N, ELK_OUT_R
         => ELK_OUT_R, ELK_OUT_F => ELK_OUT_F, CCC_160M_FXD => 
        CCC_160M_FXD, CCC_160M_ADJ => CCC_160M_ADJ, ELK_IN_DDR_R
         => ELK_IN_DDR_R, ELK_IN_DDR_F => ELK_IN_DDR_F);
    
    ELK_IN_F : DFN1C0
      port map(D => ELK_IN_DDR_F, CLK => CCC_160M_ADJ, CLR => 
        DEV_RST_B_c_1, Q => \ELK_IN_F\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    U_ELK1_SERDAT_SOURCE : SYNC_DAT_SEL_16
      port map(ELK_TX_DAT(7) => \ELK_TX_DAT[7]\, ELK_TX_DAT(6)
         => \ELK_TX_DAT[6]\, ELK_TX_DAT(5) => \ELK_TX_DAT[5]\, 
        ELK_TX_DAT(4) => \ELK_TX_DAT[4]\, ELK_TX_DAT(3) => 
        \ELK_TX_DAT[3]\, ELK_TX_DAT(2) => \ELK_TX_DAT[2]\, 
        ELK_TX_DAT(1) => \ELK_TX_DAT[1]\, ELK_TX_DAT(0) => 
        \ELK_TX_DAT[0]\, PATT_ELK_DAT_16(7) => PATT_ELK_DAT_16(7), 
        PATT_ELK_DAT_16(6) => PATT_ELK_DAT_16(6), 
        PATT_ELK_DAT_16(5) => PATT_ELK_DAT_16(5), 
        PATT_ELK_DAT_16(4) => PATT_ELK_DAT_16(4), 
        PATT_ELK_DAT_16(3) => PATT_ELK_DAT_16(3), 
        PATT_ELK_DAT_16(2) => PATT_ELK_DAT_16(2), 
        PATT_ELK_DAT_16(1) => PATT_ELK_DAT_16(1), 
        PATT_ELK_DAT_16(0) => PATT_ELK_DAT_16(0), OP_MODE_c_2_0
         => OP_MODE_c_2_0, MASTER_SALT_POR_B_i_0_i_9 => 
        MASTER_SALT_POR_B_i_0_i_9, CLK_40M_GL => CLK_40M_GL);
    
    ELK_IN_R : DFN1C0
      port map(D => ELK_IN_DDR_R, CLK => CCC_160M_ADJ, CLR => 
        DEV_RST_B_c_1, Q => \ELK_IN_R\);
    
    GND_i : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity tristate_buf_2 is

    port( P_USB_MASTER_EN_c : in    std_logic;
          USB_SIWU_BI       : in    std_logic;
          USB_SIWU_B        : out   std_logic
        );

end tristate_buf_2;

architecture DEF_ARCH of tristate_buf_2 is 

  component TRIBUFF_F_24U
    port( D   : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          PAD : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \GND\, \VCC\ : std_logic;

begin 


    \TRIBUFF_F_24U[0]\ : TRIBUFF_F_24U
      port map(D => USB_SIWU_BI, E => P_USB_MASTER_EN_c, PAD => 
        USB_SIWU_B);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    GND_i : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity DDR_BIDIR_LVDS_DUAL_CLK_0 is

    port( DCB_SALT_SEL_c_i : in    std_logic;
          ELK0_DAT_P       : inout std_logic := 'Z';
          ELK0_DAT_N       : inout std_logic := 'Z';
          ELK0_OUT_R_i_0   : in    std_logic;
          ELK0_OUT_F_i_0   : in    std_logic;
          CCC_160M_FXD     : in    std_logic;
          CCC_160M_ADJ     : in    std_logic;
          ELK0_IN_DDR_F_i  : out   std_logic;
          ELK0_IN_DDR_R_i  : out   std_logic
        );

end DDR_BIDIR_LVDS_DUAL_CLK_0;

architecture DEF_ARCH of DDR_BIDIR_LVDS_DUAL_CLK_0 is 

  component DDR_REG
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          QR  : out   std_logic;
          QF  : out   std_logic
        );
  end component;

  component DDR_OUT
    port( DR  : in    std_logic := 'U';
          DF  : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component BIBUF_LVDS
    port( PADP : inout   std_logic;
          PADN : inout   std_logic;
          D    : in    std_logic := 'U';
          E    : in    std_logic := 'U';
          Y    : out   std_logic
        );
  end component;

  component INV
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal ELK0_IN_DDR_R, ELK0_IN_DDR_F, 
        DDR_BIDIR_LVDS_DUAL_CLK_0_GND, BIBUF_LVDS_0_Y, 
        DDR_OUT_0_Q, \VCC\ : std_logic;

begin 


    DDR_REG_0 : DDR_REG
      port map(D => BIBUF_LVDS_0_Y, CLK => CCC_160M_ADJ, CLR => 
        DDR_BIDIR_LVDS_DUAL_CLK_0_GND, QR => ELK0_IN_DDR_R, QF
         => ELK0_IN_DDR_F);
    
    DDR_OUT_0 : DDR_OUT
      port map(DR => ELK0_OUT_R_i_0, DF => ELK0_OUT_F_i_0, CLK
         => CCC_160M_FXD, CLR => DDR_BIDIR_LVDS_DUAL_CLK_0_GND, Q
         => DDR_OUT_0_Q);
    
    BIBUF_LVDS_0 : BIBUF_LVDS
      port map(PADP => ELK0_DAT_P, PADN => ELK0_DAT_N, D => 
        DDR_OUT_0_Q, E => DCB_SALT_SEL_c_i, Y => BIBUF_LVDS_0_Y);
    
    DDR_REG_0_RNIDU52_0 : INV
      port map(A => ELK0_IN_DDR_R, Y => ELK0_IN_DDR_R_i);
    
    DDR_REG_0_RNIDU52 : INV
      port map(A => ELK0_IN_DDR_F, Y => ELK0_IN_DDR_F_i);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    GND_i : GND
      port map(Y => DDR_BIDIR_LVDS_DUAL_CLK_0_GND);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity LVDS_CLK_IN is

    port( CLK200_N : in    std_logic;
          CLK200_P : in    std_logic;
          Y        : out   std_logic
        );

end LVDS_CLK_IN;

architecture DEF_ARCH of LVDS_CLK_IN is 

  component INBUF_LVDS
    port( PADP : in    std_logic := 'U';
          PADN : in    std_logic := 'U';
          Y    : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \GND\, \VCC\ : std_logic;

begin 


    \INBUF_LVDS[0]\ : INBUF_LVDS
      port map(PADP => CLK200_P, PADN => CLK200_N, Y => Y);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    GND_i : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SLAVE_DES320S_1_17_17 is

    port( ELK_RX_SER_WORD_19     : out   std_logic_vector(7 downto 0);
          BIT_OS_SEL_2_0         : in    std_logic;
          BIT_OS_SEL_1           : in    std_logic_vector(2 downto 1);
          BIT_OS_SEL_0           : in    std_logic_vector(2 downto 1);
          BIT_OS_SEL_0_d0        : in    std_logic;
          CLK_40M_GL             : in    std_logic;
          CCC_160M_FXD           : in    std_logic;
          ELK_IN_R               : in    std_logic;
          ELK_IN_F               : in    std_logic;
          MASTER_DCB_POR_B_i_0_i : in    std_logic;
          CCC_160M_ADJ           : in    std_logic
        );

end SLAVE_DES320S_1_17_17;

architecture DEF_ARCH of SLAVE_DES320S_1_17_17 is 

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal N_17, \ARB_BYTE[0]_net_1\, \ARB_BYTE[4]_net_1\, N_18, 
        \ARB_BYTE[1]_net_1\, \ARB_BYTE[5]_net_1\, N_19, 
        \ARB_BYTE[2]_net_1\, \ARB_BYTE[6]_net_1\, N_20, 
        \ARB_BYTE[3]_net_1\, \ARB_BYTE[7]_net_1\, N_21, 
        \ARB_BYTE[8]_net_1\, N_22, \ARB_BYTE[9]_net_1\, N_23, 
        \ARB_BYTE[10]_net_1\, N_24, \ARB_BYTE[11]_net_1\, N_31, 
        \ARB_BYTE[12]_net_1\, N_32, \ARB_BYTE[13]_net_1\, N_33, 
        N_34, N_35, N_36, N_37, N_38, N_39, N_40, N_56, 
        \ARB_BYTE[14]_net_1\, N_64, \N_RECD_SER_WORD[0]\, 
        \N_RECD_SER_WORD[1]\, \N_RECD_SER_WORD[2]\, 
        \N_RECD_SER_WORD[3]\, \N_RECD_SER_WORD[4]\, 
        \N_RECD_SER_WORD[5]\, \N_RECD_SER_WORD[6]\, 
        \N_RECD_SER_WORD[7]\, \ADJ_SER_IN_F_0DEL\, 
        \ADJ_SER_IN_R_0DEL\, \ADJ_SER_IN_F_1DEL\, 
        \ADJ_SER_IN_R_1DEL\, \Q[0]_net_1\, \ADJ_Q[0]_net_1\, 
        \Q[1]_net_1\, \ADJ_Q[1]_net_1\, \Q[2]_net_1\, 
        \ADJ_Q[2]_net_1\, \Q[3]_net_1\, \ADJ_Q[3]_net_1\, 
        \Q[4]_net_1\, \ADJ_Q[4]_net_1\, \Q[5]_net_1\, 
        \ADJ_Q[5]_net_1\, \Q[6]_net_1\, \ADJ_Q[6]_net_1\, 
        \Q[7]_net_1\, \ADJ_Q[7]_net_1\, \Q[8]_net_1\, 
        \ADJ_Q[8]_net_1\, \Q[9]_net_1\, \ADJ_Q[9]_net_1\, 
        \Q[10]_net_1\, \ADJ_Q[10]_net_1\, \Q[11]_net_1\, 
        \ADJ_Q[11]_net_1\, \Q[12]_net_1\, \ADJ_Q[12]_net_1\, 
        \Q[13]_net_1\, \ADJ_Q[13]_net_1\, \Q[14]_net_1\, 
        \ADJ_Q[14]_net_1\, \ARB_WRD_40M_FIXED[0]_net_1\, 
        \ARB_WRD_40M_FIXED[1]_net_1\, 
        \ARB_WRD_40M_FIXED[2]_net_1\, 
        \ARB_WRD_40M_FIXED[3]_net_1\, 
        \ARB_WRD_40M_FIXED[4]_net_1\, 
        \ARB_WRD_40M_FIXED[5]_net_1\, 
        \ARB_WRD_40M_FIXED[6]_net_1\, 
        \ARB_WRD_40M_FIXED[7]_net_1\, 
        \ARB_WRD_40M_FIXED[8]_net_1\, 
        \ARB_WRD_40M_FIXED[9]_net_1\, 
        \ARB_WRD_40M_FIXED[10]_net_1\, 
        \ARB_WRD_40M_FIXED[11]_net_1\, 
        \ARB_WRD_40M_FIXED[12]_net_1\, 
        \ARB_WRD_40M_FIXED[13]_net_1\, 
        \ARB_WRD_40M_FIXED[14]_net_1\, \GND\, \VCC\ : std_logic;

begin 


    \RECD_SER_WORD_RNO[5]\ : MX2
      port map(A => N_38, B => N_39, S => BIT_OS_SEL_2_0, Y => 
        \N_RECD_SER_WORD[5]\);
    
    \ARB_WRD_40M_FIXED[9]\ : DFN1C0
      port map(D => \Q[9]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[9]_net_1\);
    
    \ADJ_Q[4]\ : DFN1C0
      port map(D => \ADJ_Q[2]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[4]_net_1\);
    
    \ARB_BYTE_RNIODBS1[5]\ : MX2
      port map(A => N_22, B => N_24, S => BIT_OS_SEL_0(1), Y => 
        N_38);
    
    \ARB_BYTE[6]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[6]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[6]_net_1\);
    
    ADJ_SER_IN_F_1DEL : DFN1C0
      port map(D => \ADJ_SER_IN_F_0DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_F_1DEL\);
    
    \ARB_BYTE[0]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[0]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[0]_net_1\);
    
    \Q[11]\ : DFN1C0
      port map(D => \ADJ_Q[11]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[11]_net_1\);
    
    \ARB_BYTE_RNIVDQ21[13]\ : MX2
      port map(A => \ARB_BYTE[9]_net_1\, B => 
        \ARB_BYTE[13]_net_1\, S => BIT_OS_SEL_0(2), Y => N_32);
    
    \ARB_BYTE_RNICJHS[11]\ : MX2
      port map(A => \ARB_BYTE[7]_net_1\, B => 
        \ARB_BYTE[11]_net_1\, S => BIT_OS_SEL_0_d0, Y => N_24);
    
    \ADJ_Q[8]\ : DFN1C0
      port map(D => \ADJ_Q[6]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[8]_net_1\);
    
    \ARB_BYTE_RNIM3ID2[13]\ : MX2
      port map(A => N_24, B => N_32, S => BIT_OS_SEL_0(1), Y => 
        N_40);
    
    \ARB_BYTE_RNIK9BS1[4]\ : MX2
      port map(A => N_21, B => N_23, S => BIT_OS_SEL_0(1), Y => 
        N_37);
    
    \ADJ_Q[6]\ : DFN1C0
      port map(D => \ADJ_Q[4]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[6]_net_1\);
    
    \ADJ_Q[12]\ : DFN1C0
      port map(D => \ADJ_Q[10]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[12]_net_1\);
    
    \RECD_SER_WORD_RNO_1[0]\ : MX2
      port map(A => \ARB_BYTE[0]_net_1\, B => \ARB_BYTE[4]_net_1\, 
        S => BIT_OS_SEL_0_d0, Y => N_17);
    
    \ARB_BYTE_RNIAHHS[6]\ : MX2
      port map(A => \ARB_BYTE[6]_net_1\, B => 
        \ARB_BYTE[10]_net_1\, S => BIT_OS_SEL_0_d0, Y => N_23);
    
    \Q[1]\ : DFN1C0
      port map(D => \ADJ_Q[1]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[1]_net_1\);
    
    \ARB_BYTE_RNIIVHD2[6]\ : MX2
      port map(A => N_23, B => N_31, S => BIT_OS_SEL_0(1), Y => 
        N_39);
    
    \ARB_BYTE[4]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[4]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[4]_net_1\);
    
    \ADJ_Q[2]\ : DFN1C0
      port map(D => \ADJ_Q[0]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[2]_net_1\);
    
    \RECD_SER_WORD_RNO_1[7]\ : MX2
      port map(A => \ARB_BYTE[10]_net_1\, B => 
        \ARB_BYTE[14]_net_1\, S => BIT_OS_SEL_1(2), Y => N_56);
    
    \RECD_SER_WORD[4]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[4]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_19(4));
    
    \Q[5]\ : DFN1C0
      port map(D => \ADJ_Q[5]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[5]_net_1\);
    
    \ADJ_Q[11]\ : DFN1C0
      port map(D => \ADJ_Q[9]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[11]_net_1\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \ADJ_Q[3]\ : DFN1C0
      port map(D => \ADJ_Q[1]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[3]_net_1\);
    
    \Q[10]\ : DFN1C0
      port map(D => \ADJ_Q[10]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[10]_net_1\);
    
    \ARB_WRD_40M_FIXED[6]\ : DFN1C0
      port map(D => \Q[6]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[6]_net_1\);
    
    \ARB_WRD_40M_FIXED[1]\ : DFN1C0
      port map(D => \Q[1]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[1]_net_1\);
    
    \RECD_SER_WORD[3]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[3]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_19(3));
    
    \RECD_SER_WORD[0]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[0]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_19(0));
    
    \RECD_SER_WORD_RNO[3]\ : MX2
      port map(A => N_36, B => N_37, S => BIT_OS_SEL_2_0, Y => 
        \N_RECD_SER_WORD[3]\);
    
    \Q[0]\ : DFN1C0
      port map(D => \ADJ_Q[0]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[0]_net_1\);
    
    \RECD_SER_WORD_RNO_0[7]\ : MX2
      port map(A => N_31, B => N_56, S => BIT_OS_SEL_1(1), Y => 
        N_64);
    
    \Q[7]\ : DFN1C0
      port map(D => \ADJ_Q[7]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[7]_net_1\);
    
    \ARB_BYTE[14]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[14]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[14]_net_1\);
    
    \ARB_WRD_40M_FIXED[2]\ : DFN1C0
      port map(D => \Q[2]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[2]_net_1\);
    
    \ARB_WRD_40M_FIXED[14]\ : DFN1C0
      port map(D => \Q[14]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[14]_net_1\);
    
    \RECD_SER_WORD_RNO[2]\ : MX2
      port map(A => N_35, B => N_36, S => BIT_OS_SEL_2_0, Y => 
        \N_RECD_SER_WORD[2]\);
    
    \ARB_BYTE[2]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[2]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[2]_net_1\);
    
    \ADJ_Q[7]\ : DFN1C0
      port map(D => \ADJ_Q[5]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[7]_net_1\);
    
    \ARB_BYTE[8]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[8]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[8]_net_1\);
    
    \RECD_SER_WORD[5]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[5]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_19(5));
    
    \ARB_BYTE[12]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[12]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[12]_net_1\);
    
    \RECD_SER_WORD[1]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[1]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_19(1));
    
    \Q[3]\ : DFN1C0
      port map(D => \ADJ_Q[3]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[3]_net_1\);
    
    \ARB_BYTE_RNIRHJH[2]\ : MX2
      port map(A => \ARB_BYTE[2]_net_1\, B => \ARB_BYTE[6]_net_1\, 
        S => BIT_OS_SEL_0_d0, Y => N_19);
    
    \ARB_BYTE_RNIVLJH[4]\ : MX2
      port map(A => \ARB_BYTE[4]_net_1\, B => \ARB_BYTE[8]_net_1\, 
        S => BIT_OS_SEL_0_d0, Y => N_21);
    
    ADJ_SER_IN_F_0DEL : DFN1C0
      port map(D => ELK_IN_F, CLK => CCC_160M_ADJ, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_F_0DEL\);
    
    \RECD_SER_WORD_RNO[7]\ : MX2
      port map(A => N_40, B => N_64, S => BIT_OS_SEL_2_0, Y => 
        \N_RECD_SER_WORD[7]\);
    
    \RECD_SER_WORD_RNO[1]\ : MX2
      port map(A => N_34, B => N_35, S => BIT_OS_SEL_2_0, Y => 
        \N_RECD_SER_WORD[1]\);
    
    \ARB_WRD_40M_FIXED[4]\ : DFN1C0
      port map(D => \Q[4]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[4]_net_1\);
    
    \RECD_SER_WORD_RNO[0]\ : MX2
      port map(A => N_33, B => N_34, S => BIT_OS_SEL_2_0, Y => 
        \N_RECD_SER_WORD[0]\);
    
    \Q[6]\ : DFN1C0
      port map(D => \ADJ_Q[6]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[6]_net_1\);
    
    \ARB_BYTE_RNI16DH1[1]\ : MX2
      port map(A => N_18, B => N_20, S => BIT_OS_SEL_0(1), Y => 
        N_34);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \ARB_WRD_40M_FIXED[8]\ : DFN1C0
      port map(D => \Q[8]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[8]_net_1\);
    
    \ARB_BYTE[11]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[11]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[11]_net_1\);
    
    \Q[9]\ : DFN1C0
      port map(D => \ADJ_Q[9]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[9]_net_1\);
    
    \Q[14]\ : DFN1C0
      port map(D => \ADJ_Q[14]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[14]_net_1\);
    
    ADJ_SER_IN_R_0DEL : DFN1C0
      port map(D => ELK_IN_R, CLK => CCC_160M_ADJ, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_R_0DEL\);
    
    \Q[13]\ : DFN1C0
      port map(D => \ADJ_Q[13]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[13]_net_1\);
    
    \ARB_BYTE_RNI1OJH[5]\ : MX2
      port map(A => \ARB_BYTE[5]_net_1\, B => \ARB_BYTE[9]_net_1\, 
        S => BIT_OS_SEL_0_d0, Y => N_22);
    
    \ARB_BYTE[9]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[9]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[9]_net_1\);
    
    ADJ_SER_IN_R_1DEL : DFN1C0
      port map(D => \ADJ_SER_IN_R_0DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_R_1DEL\);
    
    \ARB_BYTE[10]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[10]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[10]_net_1\);
    
    \ADJ_Q[9]\ : DFN1C0
      port map(D => \ADJ_Q[7]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[9]_net_1\);
    
    \RECD_SER_WORD[7]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[7]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_19(7));
    
    \ARB_WRD_40M_FIXED[5]\ : DFN1C0
      port map(D => \Q[5]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[5]_net_1\);
    
    \ARB_WRD_40M_FIXED[12]\ : DFN1C0
      port map(D => \Q[12]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[12]_net_1\);
    
    \ARB_WRD_40M_FIXED[11]\ : DFN1C0
      port map(D => \Q[11]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[11]_net_1\);
    
    \ARB_WRD_40M_FIXED[0]\ : DFN1C0
      port map(D => \Q[0]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[0]_net_1\);
    
    \ADJ_Q[10]\ : DFN1C0
      port map(D => \ADJ_Q[8]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[10]_net_1\);
    
    \Q[2]\ : DFN1C0
      port map(D => \ADJ_Q[2]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[2]_net_1\);
    
    \ARB_BYTE_RNI9EDH1[3]\ : MX2
      port map(A => N_20, B => N_22, S => BIT_OS_SEL_0(1), Y => 
        N_36);
    
    \ARB_BYTE_RNITBQ21[12]\ : MX2
      port map(A => \ARB_BYTE[8]_net_1\, B => 
        \ARB_BYTE[12]_net_1\, S => BIT_OS_SEL_0(2), Y => N_31);
    
    \ADJ_Q[1]\ : DFN1C0
      port map(D => \ADJ_SER_IN_F_1DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[1]_net_1\);
    
    \RECD_SER_WORD[6]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[6]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_19(6));
    
    \ARB_BYTE_RNI5ADH1[2]\ : MX2
      port map(A => N_19, B => N_21, S => BIT_OS_SEL_0(1), Y => 
        N_35);
    
    \RECD_SER_WORD[2]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[2]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_19(2));
    
    \ADJ_Q[13]\ : DFN1C0
      port map(D => \ADJ_Q[11]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[13]_net_1\);
    
    \ARB_BYTE_RNITJJH[3]\ : MX2
      port map(A => \ARB_BYTE[3]_net_1\, B => \ARB_BYTE[7]_net_1\, 
        S => BIT_OS_SEL_0_d0, Y => N_20);
    
    \Q[8]\ : DFN1C0
      port map(D => \ADJ_Q[8]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[8]_net_1\);
    
    \ARB_BYTE[5]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[5]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[5]_net_1\);
    
    \ADJ_Q[14]\ : DFN1C0
      port map(D => \ADJ_Q[12]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[14]_net_1\);
    
    \RECD_SER_WORD_RNO[4]\ : MX2
      port map(A => N_37, B => N_38, S => BIT_OS_SEL_2_0, Y => 
        \N_RECD_SER_WORD[4]\);
    
    \Q[12]\ : DFN1C0
      port map(D => \ADJ_Q[12]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[12]_net_1\);
    
    \ARB_BYTE[13]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[13]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[13]_net_1\);
    
    \ARB_WRD_40M_FIXED[3]\ : DFN1C0
      port map(D => \Q[3]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[3]_net_1\);
    
    \ARB_BYTE[7]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[7]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[7]_net_1\);
    
    \RECD_SER_WORD_RNO_0[0]\ : MX2
      port map(A => N_17, B => N_19, S => BIT_OS_SEL_0(1), Y => 
        N_33);
    
    \Q[4]\ : DFN1C0
      port map(D => \ADJ_Q[4]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[4]_net_1\);
    
    \ARB_WRD_40M_FIXED[7]\ : DFN1C0
      port map(D => \Q[7]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[7]_net_1\);
    
    \RECD_SER_WORD_RNO[6]\ : MX2
      port map(A => N_39, B => N_40, S => BIT_OS_SEL_2_0, Y => 
        \N_RECD_SER_WORD[6]\);
    
    \ARB_BYTE_RNIPFJH[1]\ : MX2
      port map(A => \ARB_BYTE[1]_net_1\, B => \ARB_BYTE[5]_net_1\, 
        S => BIT_OS_SEL_0_d0, Y => N_18);
    
    \ARB_BYTE[3]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[3]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[3]_net_1\);
    
    \ADJ_Q[5]\ : DFN1C0
      port map(D => \ADJ_Q[3]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[5]_net_1\);
    
    \ARB_BYTE[1]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[1]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[1]_net_1\);
    
    \ARB_WRD_40M_FIXED[13]\ : DFN1C0
      port map(D => \Q[13]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[13]_net_1\);
    
    \ADJ_Q[0]\ : DFN1C0
      port map(D => \ADJ_SER_IN_R_1DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[0]_net_1\);
    
    \ARB_WRD_40M_FIXED[10]\ : DFN1C0
      port map(D => \Q[10]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[10]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SER320M_3_34_19 is

    port( ELK_TX_DAT                 : in    std_logic_vector(7 downto 0);
          MASTER_SALT_POR_B_i_0_i_4  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_7  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_0  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_8  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_12 : in    std_logic;
          ELK_OUT_R                  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_16 : in    std_logic;
          ELK_OUT_F                  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_10 : in    std_logic;
          CCC_160M_FXD               : in    std_logic;
          CLK_40M_GL                 : in    std_logic
        );

end SER320M_3_34_19;

architecture DEF_ARCH of SER320M_3_34_19 is 

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \N_SER_CMD_WORD_R[0]\, \START_RISE\, 
        \N_SER_CMD_WORD_F[0]\, \N_SER_CMD_WORD_R[3]\, 
        \SER_CMD_WORD_R[2]_net_1\, \N_SER_CMD_WORD_R[2]\, 
        \SER_CMD_WORD_R[1]_net_1\, \N_SER_CMD_WORD_R[1]\, 
        \SER_CMD_WORD_R[0]_net_1\, \N_SER_CMD_WORD_F[3]\, 
        \SER_CMD_WORD_F[2]_net_1\, \N_SER_CMD_WORD_F[2]\, 
        \SER_CMD_WORD_F[1]_net_1\, \N_SER_CMD_WORD_F[1]\, 
        \SER_CMD_WORD_F[0]_net_1\, N_START_RISE, 
        \CLK40M_GEN_DEL0\, \SER_OUT_FI\, \SER_OUT_RI\, 
        \SER_CMD_WORD_F[3]_net_1\, \SER_CMD_WORD_R[3]_net_1\, 
        \GND\, \VCC\ : std_logic;

begin 


    SER_OUT_FI : DFN1C0
      port map(D => \SER_CMD_WORD_F[3]_net_1\, CLK => 
        CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_0, Q => 
        \SER_OUT_FI\);
    
    \SER_CMD_WORD_F[3]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[3]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_7, Q => 
        \SER_CMD_WORD_F[3]_net_1\);
    
    \SER_CMD_WORD_R[1]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[1]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_4, Q => 
        \SER_CMD_WORD_R[1]_net_1\);
    
    \SER_CMD_WORD_R[2]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[2]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_4, Q => 
        \SER_CMD_WORD_R[2]_net_1\);
    
    \SER_CMD_WORD_R_RNO[3]\ : MX2
      port map(A => \SER_CMD_WORD_R[2]_net_1\, B => ELK_TX_DAT(7), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_R[3]\);
    
    \SER_CMD_WORD_R_RNO[0]\ : NOR2B
      port map(A => \START_RISE\, B => ELK_TX_DAT(1), Y => 
        \N_SER_CMD_WORD_R[0]\);
    
    \SER_CMD_WORD_F[0]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[0]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_7, Q => 
        \SER_CMD_WORD_F[0]_net_1\);
    
    \SER_CMD_WORD_R_RNO[1]\ : MX2
      port map(A => \SER_CMD_WORD_R[0]_net_1\, B => ELK_TX_DAT(3), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_R[1]\);
    
    \SER_CMD_WORD_F_RNO[2]\ : MX2
      port map(A => \SER_CMD_WORD_F[1]_net_1\, B => ELK_TX_DAT(4), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_F[2]\);
    
    \SER_CMD_WORD_F_RNO[3]\ : MX2
      port map(A => \SER_CMD_WORD_F[2]_net_1\, B => ELK_TX_DAT(6), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_F[3]\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    CLK40M_GEN_DEL0 : DFN1C0
      port map(D => CLK_40M_GL, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_10, Q => \CLK40M_GEN_DEL0\);
    
    SER_OUT_RI : DFN1C0
      port map(D => \SER_CMD_WORD_R[3]_net_1\, CLK => 
        CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_0, Q => 
        \SER_OUT_RI\);
    
    \SER_CMD_WORD_F[2]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[2]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_7, Q => 
        \SER_CMD_WORD_F[2]_net_1\);
    
    \SER_CMD_WORD_F_RNO[1]\ : MX2
      port map(A => \SER_CMD_WORD_F[0]_net_1\, B => ELK_TX_DAT(2), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_F[1]\);
    
    \SER_CMD_WORD_R[0]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[0]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_4, Q => 
        \SER_CMD_WORD_R[0]_net_1\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    START_RISE : DFN1C0
      port map(D => N_START_RISE, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_8, Q => \START_RISE\);
    
    \SER_CMD_WORD_R[3]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[3]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_4, Q => 
        \SER_CMD_WORD_R[3]_net_1\);
    
    \SER_CMD_WORD_F_RNO[0]\ : NOR2B
      port map(A => \START_RISE\, B => ELK_TX_DAT(0), Y => 
        \N_SER_CMD_WORD_F[0]\);
    
    SER_OUT_RDEL : DFN1C0
      port map(D => \SER_OUT_RI\, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_12, Q => ELK_OUT_R);
    
    \SER_CMD_WORD_F[1]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[1]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_7, Q => 
        \SER_CMD_WORD_F[1]_net_1\);
    
    START_RISE_RNO : NOR2B
      port map(A => \CLK40M_GEN_DEL0\, B => CLK_40M_GL, Y => 
        N_START_RISE);
    
    \SER_CMD_WORD_R_RNO[2]\ : MX2
      port map(A => \SER_CMD_WORD_R[1]_net_1\, B => ELK_TX_DAT(5), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_R[2]\);
    
    SER_OUT_FDEL : DFN1C0
      port map(D => \SER_OUT_FI\, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_16, Q => ELK_OUT_F);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity DDR_BIDIR_LVDS_DUAL_CLK_19 is

    port( DCB_SALT_SEL_c_i : in    std_logic;
          ELK19_DAT_P      : inout std_logic := 'Z';
          ELK19_DAT_N      : inout std_logic := 'Z';
          ELK_OUT_R        : in    std_logic;
          ELK_OUT_F        : in    std_logic;
          CCC_160M_FXD     : in    std_logic;
          CCC_160M_ADJ     : in    std_logic;
          ELK_IN_DDR_R     : out   std_logic;
          ELK_IN_DDR_F     : out   std_logic
        );

end DDR_BIDIR_LVDS_DUAL_CLK_19;

architecture DEF_ARCH of DDR_BIDIR_LVDS_DUAL_CLK_19 is 

  component DDR_REG
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          QR  : out   std_logic;
          QF  : out   std_logic
        );
  end component;

  component DDR_OUT
    port( DR  : in    std_logic := 'U';
          DF  : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component BIBUF_LVDS
    port( PADP : inout   std_logic;
          PADN : inout   std_logic;
          D    : in    std_logic := 'U';
          E    : in    std_logic := 'U';
          Y    : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal DDR_BIDIR_LVDS_DUAL_CLK_19_GND, BIBUF_LVDS_0_Y, 
        DDR_OUT_0_Q, \VCC\ : std_logic;

begin 


    DDR_REG_0 : DDR_REG
      port map(D => BIBUF_LVDS_0_Y, CLK => CCC_160M_ADJ, CLR => 
        DDR_BIDIR_LVDS_DUAL_CLK_19_GND, QR => ELK_IN_DDR_R, QF
         => ELK_IN_DDR_F);
    
    DDR_OUT_0 : DDR_OUT
      port map(DR => ELK_OUT_R, DF => ELK_OUT_F, CLK => 
        CCC_160M_FXD, CLR => DDR_BIDIR_LVDS_DUAL_CLK_19_GND, Q
         => DDR_OUT_0_Q);
    
    BIBUF_LVDS_0 : BIBUF_LVDS
      port map(PADP => ELK19_DAT_P, PADN => ELK19_DAT_N, D => 
        DDR_OUT_0_Q, E => DCB_SALT_SEL_c_i, Y => BIBUF_LVDS_0_Y);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    GND_i : GND
      port map(Y => DDR_BIDIR_LVDS_DUAL_CLK_19_GND);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SYNC_DAT_SEL_19 is

    port( ELK_TX_DAT                 : out   std_logic_vector(7 downto 0);
          PATT_ELK_DAT_19            : in    std_logic_vector(7 downto 0);
          OP_MODE_c_6_0              : in    std_logic;
          OP_MODE_c_5_0              : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_15 : in    std_logic;
          CLK_40M_GL                 : in    std_logic
        );

end SYNC_DAT_SEL_19;

architecture DEF_ARCH of SYNC_DAT_SEL_19 is 

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \N_SERDAT[0]\, \N_SERDAT[1]\, \N_SERDAT[2]\, 
        \N_SERDAT[3]\, \N_SERDAT[4]\, \N_SERDAT[5]\, 
        \N_SERDAT[6]\, \N_SERDAT[7]\, \GND\, \VCC\ : std_logic;

begin 


    \SERDAT_RNO[4]\ : NOR2A
      port map(A => PATT_ELK_DAT_19(4), B => OP_MODE_c_6_0, Y => 
        \N_SERDAT[4]\);
    
    \SERDAT_RNO[0]\ : NOR2A
      port map(A => PATT_ELK_DAT_19(0), B => OP_MODE_c_5_0, Y => 
        \N_SERDAT[0]\);
    
    \SERDAT[6]\ : DFN1C0
      port map(D => \N_SERDAT[6]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_15, Q => ELK_TX_DAT(6));
    
    \SERDAT[4]\ : DFN1C0
      port map(D => \N_SERDAT[4]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_15, Q => ELK_TX_DAT(4));
    
    \SERDAT_RNO[7]\ : OR2
      port map(A => PATT_ELK_DAT_19(7), B => OP_MODE_c_6_0, Y => 
        \N_SERDAT[7]\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \SERDAT_RNO[3]\ : OR2
      port map(A => PATT_ELK_DAT_19(3), B => OP_MODE_c_5_0, Y => 
        \N_SERDAT[3]\);
    
    \SERDAT_RNO[2]\ : OR2
      port map(A => PATT_ELK_DAT_19(2), B => OP_MODE_c_5_0, Y => 
        \N_SERDAT[2]\);
    
    \SERDAT[5]\ : DFN1C0
      port map(D => \N_SERDAT[5]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_15, Q => ELK_TX_DAT(5));
    
    \SERDAT[7]\ : DFN1C0
      port map(D => \N_SERDAT[7]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_15, Q => ELK_TX_DAT(7));
    
    GND_i : GND
      port map(Y => \GND\);
    
    \SERDAT_RNO[5]\ : NOR2A
      port map(A => PATT_ELK_DAT_19(5), B => OP_MODE_c_6_0, Y => 
        \N_SERDAT[5]\);
    
    \SERDAT[0]\ : DFN1C0
      port map(D => \N_SERDAT[0]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_15, Q => ELK_TX_DAT(0));
    
    \SERDAT_RNO[6]\ : NOR2A
      port map(A => PATT_ELK_DAT_19(6), B => OP_MODE_c_6_0, Y => 
        \N_SERDAT[6]\);
    
    \SERDAT[1]\ : DFN1C0
      port map(D => \N_SERDAT[1]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_15, Q => ELK_TX_DAT(1));
    
    \SERDAT_RNO[1]\ : OR2
      port map(A => PATT_ELK_DAT_19(1), B => OP_MODE_c_5_0, Y => 
        \N_SERDAT[1]\);
    
    \SERDAT[3]\ : DFN1C0
      port map(D => \N_SERDAT[3]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_15, Q => ELK_TX_DAT(3));
    
    \SERDAT[2]\ : DFN1C0
      port map(D => \N_SERDAT[2]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_15, Q => ELK_TX_DAT(2));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity ELINK_SLAVE_15_14 is

    port( BIT_OS_SEL_0_d0            : in    std_logic;
          BIT_OS_SEL_0               : in    std_logic_vector(2 downto 1);
          BIT_OS_SEL_1               : in    std_logic_vector(2 downto 1);
          BIT_OS_SEL_2_0             : in    std_logic;
          ELK_RX_SER_WORD_19         : out   std_logic_vector(7 downto 0);
          OP_MODE_c_5_0              : in    std_logic;
          OP_MODE_c_6_0              : in    std_logic;
          PATT_ELK_DAT_19            : in    std_logic_vector(7 downto 0);
          MASTER_DCB_POR_B_i_0_i     : in    std_logic;
          ELK19_DAT_N                : inout std_logic := 'Z';
          ELK19_DAT_P                : inout std_logic := 'Z';
          DCB_SALT_SEL_c_i           : in    std_logic;
          CCC_160M_FXD               : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_10 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_16 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_12 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_8  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_0  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_7  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_4  : in    std_logic;
          CLK_40M_GL                 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_15 : in    std_logic;
          DEV_RST_B_c_0              : in    std_logic;
          CCC_160M_ADJ               : in    std_logic
        );

end ELINK_SLAVE_15_14;

architecture DEF_ARCH of ELINK_SLAVE_15_14 is 

  component SLAVE_DES320S_1_17_17
    port( ELK_RX_SER_WORD_19     : out   std_logic_vector(7 downto 0);
          BIT_OS_SEL_2_0         : in    std_logic := 'U';
          BIT_OS_SEL_1           : in    std_logic_vector(2 downto 1) := (others => 'U');
          BIT_OS_SEL_0           : in    std_logic_vector(2 downto 1) := (others => 'U');
          BIT_OS_SEL_0_d0        : in    std_logic := 'U';
          CLK_40M_GL             : in    std_logic := 'U';
          CCC_160M_FXD           : in    std_logic := 'U';
          ELK_IN_R               : in    std_logic := 'U';
          ELK_IN_F               : in    std_logic := 'U';
          MASTER_DCB_POR_B_i_0_i : in    std_logic := 'U';
          CCC_160M_ADJ           : in    std_logic := 'U'
        );
  end component;

  component SER320M_3_34_19
    port( ELK_TX_DAT                 : in    std_logic_vector(7 downto 0) := (others => 'U');
          MASTER_SALT_POR_B_i_0_i_4  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_7  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_0  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_8  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_12 : in    std_logic := 'U';
          ELK_OUT_R                  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_16 : in    std_logic := 'U';
          ELK_OUT_F                  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_10 : in    std_logic := 'U';
          CCC_160M_FXD               : in    std_logic := 'U';
          CLK_40M_GL                 : in    std_logic := 'U'
        );
  end component;

  component DDR_BIDIR_LVDS_DUAL_CLK_19
    port( DCB_SALT_SEL_c_i : in    std_logic := 'U';
          ELK19_DAT_P      : inout   std_logic;
          ELK19_DAT_N      : inout   std_logic;
          ELK_OUT_R        : in    std_logic := 'U';
          ELK_OUT_F        : in    std_logic := 'U';
          CCC_160M_FXD     : in    std_logic := 'U';
          CCC_160M_ADJ     : in    std_logic := 'U';
          ELK_IN_DDR_R     : out   std_logic;
          ELK_IN_DDR_F     : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component SYNC_DAT_SEL_19
    port( ELK_TX_DAT                 : out   std_logic_vector(7 downto 0);
          PATT_ELK_DAT_19            : in    std_logic_vector(7 downto 0) := (others => 'U');
          OP_MODE_c_6_0              : in    std_logic := 'U';
          OP_MODE_c_5_0              : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_15 : in    std_logic := 'U';
          CLK_40M_GL                 : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \ELK_IN_F\, ELK_IN_DDR_F, \ELK_IN_R\, ELK_IN_DDR_R, 
        \ELK_TX_DAT[0]\, \ELK_TX_DAT[1]\, \ELK_TX_DAT[2]\, 
        \ELK_TX_DAT[3]\, \ELK_TX_DAT[4]\, \ELK_TX_DAT[5]\, 
        \ELK_TX_DAT[6]\, \ELK_TX_DAT[7]\, ELK_OUT_R, ELK_OUT_F, 
        \GND\, \VCC\ : std_logic;

    for all : SLAVE_DES320S_1_17_17
	Use entity work.SLAVE_DES320S_1_17_17(DEF_ARCH);
    for all : SER320M_3_34_19
	Use entity work.SER320M_3_34_19(DEF_ARCH);
    for all : DDR_BIDIR_LVDS_DUAL_CLK_19
	Use entity work.DDR_BIDIR_LVDS_DUAL_CLK_19(DEF_ARCH);
    for all : SYNC_DAT_SEL_19
	Use entity work.SYNC_DAT_SEL_19(DEF_ARCH);
begin 


    U_SLAVE_1ELK : SLAVE_DES320S_1_17_17
      port map(ELK_RX_SER_WORD_19(7) => ELK_RX_SER_WORD_19(7), 
        ELK_RX_SER_WORD_19(6) => ELK_RX_SER_WORD_19(6), 
        ELK_RX_SER_WORD_19(5) => ELK_RX_SER_WORD_19(5), 
        ELK_RX_SER_WORD_19(4) => ELK_RX_SER_WORD_19(4), 
        ELK_RX_SER_WORD_19(3) => ELK_RX_SER_WORD_19(3), 
        ELK_RX_SER_WORD_19(2) => ELK_RX_SER_WORD_19(2), 
        ELK_RX_SER_WORD_19(1) => ELK_RX_SER_WORD_19(1), 
        ELK_RX_SER_WORD_19(0) => ELK_RX_SER_WORD_19(0), 
        BIT_OS_SEL_2_0 => BIT_OS_SEL_2_0, BIT_OS_SEL_1(2) => 
        BIT_OS_SEL_1(2), BIT_OS_SEL_1(1) => BIT_OS_SEL_1(1), 
        BIT_OS_SEL_0(2) => BIT_OS_SEL_0(2), BIT_OS_SEL_0(1) => 
        BIT_OS_SEL_0(1), BIT_OS_SEL_0_d0 => BIT_OS_SEL_0_d0, 
        CLK_40M_GL => CLK_40M_GL, CCC_160M_FXD => CCC_160M_FXD, 
        ELK_IN_R => \ELK_IN_R\, ELK_IN_F => \ELK_IN_F\, 
        MASTER_DCB_POR_B_i_0_i => MASTER_DCB_POR_B_i_0_i, 
        CCC_160M_ADJ => CCC_160M_ADJ);
    
    U_ELK1_CMD_TX : SER320M_3_34_19
      port map(ELK_TX_DAT(7) => \ELK_TX_DAT[7]\, ELK_TX_DAT(6)
         => \ELK_TX_DAT[6]\, ELK_TX_DAT(5) => \ELK_TX_DAT[5]\, 
        ELK_TX_DAT(4) => \ELK_TX_DAT[4]\, ELK_TX_DAT(3) => 
        \ELK_TX_DAT[3]\, ELK_TX_DAT(2) => \ELK_TX_DAT[2]\, 
        ELK_TX_DAT(1) => \ELK_TX_DAT[1]\, ELK_TX_DAT(0) => 
        \ELK_TX_DAT[0]\, MASTER_SALT_POR_B_i_0_i_4 => 
        MASTER_SALT_POR_B_i_0_i_4, MASTER_SALT_POR_B_i_0_i_7 => 
        MASTER_SALT_POR_B_i_0_i_7, MASTER_SALT_POR_B_i_0_i_0 => 
        MASTER_SALT_POR_B_i_0_i_0, MASTER_SALT_POR_B_i_0_i_8 => 
        MASTER_SALT_POR_B_i_0_i_8, MASTER_SALT_POR_B_i_0_i_12 => 
        MASTER_SALT_POR_B_i_0_i_12, ELK_OUT_R => ELK_OUT_R, 
        MASTER_SALT_POR_B_i_0_i_16 => MASTER_SALT_POR_B_i_0_i_16, 
        ELK_OUT_F => ELK_OUT_F, MASTER_SALT_POR_B_i_0_i_10 => 
        MASTER_SALT_POR_B_i_0_i_10, CCC_160M_FXD => CCC_160M_FXD, 
        CLK_40M_GL => CLK_40M_GL);
    
    U_DDR_ELK1 : DDR_BIDIR_LVDS_DUAL_CLK_19
      port map(DCB_SALT_SEL_c_i => DCB_SALT_SEL_c_i, ELK19_DAT_P
         => ELK19_DAT_P, ELK19_DAT_N => ELK19_DAT_N, ELK_OUT_R
         => ELK_OUT_R, ELK_OUT_F => ELK_OUT_F, CCC_160M_FXD => 
        CCC_160M_FXD, CCC_160M_ADJ => CCC_160M_ADJ, ELK_IN_DDR_R
         => ELK_IN_DDR_R, ELK_IN_DDR_F => ELK_IN_DDR_F);
    
    ELK_IN_F : DFN1C0
      port map(D => ELK_IN_DDR_F, CLK => CCC_160M_ADJ, CLR => 
        DEV_RST_B_c_0, Q => \ELK_IN_F\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    U_ELK1_SERDAT_SOURCE : SYNC_DAT_SEL_19
      port map(ELK_TX_DAT(7) => \ELK_TX_DAT[7]\, ELK_TX_DAT(6)
         => \ELK_TX_DAT[6]\, ELK_TX_DAT(5) => \ELK_TX_DAT[5]\, 
        ELK_TX_DAT(4) => \ELK_TX_DAT[4]\, ELK_TX_DAT(3) => 
        \ELK_TX_DAT[3]\, ELK_TX_DAT(2) => \ELK_TX_DAT[2]\, 
        ELK_TX_DAT(1) => \ELK_TX_DAT[1]\, ELK_TX_DAT(0) => 
        \ELK_TX_DAT[0]\, PATT_ELK_DAT_19(7) => PATT_ELK_DAT_19(7), 
        PATT_ELK_DAT_19(6) => PATT_ELK_DAT_19(6), 
        PATT_ELK_DAT_19(5) => PATT_ELK_DAT_19(5), 
        PATT_ELK_DAT_19(4) => PATT_ELK_DAT_19(4), 
        PATT_ELK_DAT_19(3) => PATT_ELK_DAT_19(3), 
        PATT_ELK_DAT_19(2) => PATT_ELK_DAT_19(2), 
        PATT_ELK_DAT_19(1) => PATT_ELK_DAT_19(1), 
        PATT_ELK_DAT_19(0) => PATT_ELK_DAT_19(0), OP_MODE_c_6_0
         => OP_MODE_c_6_0, OP_MODE_c_5_0 => OP_MODE_c_5_0, 
        MASTER_SALT_POR_B_i_0_i_15 => MASTER_SALT_POR_B_i_0_i_15, 
        CLK_40M_GL => CLK_40M_GL);
    
    ELK_IN_R : DFN1C0
      port map(D => ELK_IN_DDR_R, CLK => CCC_160M_ADJ, CLR => 
        DEV_RST_B_c_0, Q => \ELK_IN_R\);
    
    GND_i : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SLAVE_DES320S_1_17_7 is

    port( ELK_RX_SER_WORD_9      : out   std_logic_vector(7 downto 0);
          BIT_OS_SEL_4_0         : in    std_logic;
          BIT_OS_SEL_5           : in    std_logic_vector(2 downto 1);
          BIT_OS_SEL_3           : in    std_logic_vector(2 downto 1);
          BIT_OS_SEL_2           : in    std_logic_vector(2 downto 1);
          CLK_40M_GL             : in    std_logic;
          CCC_160M_FXD           : in    std_logic;
          ELK_IN_R               : in    std_logic;
          ELK_IN_F               : in    std_logic;
          MASTER_DCB_POR_B_i_0_i : in    std_logic;
          CCC_160M_ADJ           : in    std_logic
        );

end SLAVE_DES320S_1_17_7;

architecture DEF_ARCH of SLAVE_DES320S_1_17_7 is 

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal N_17, \ARB_BYTE[0]_net_1\, \ARB_BYTE[4]_net_1\, N_18, 
        \ARB_BYTE[1]_net_1\, \ARB_BYTE[5]_net_1\, N_19, 
        \ARB_BYTE[2]_net_1\, \ARB_BYTE[6]_net_1\, N_20, 
        \ARB_BYTE[3]_net_1\, \ARB_BYTE[7]_net_1\, N_21, 
        \ARB_BYTE[8]_net_1\, N_22, \ARB_BYTE[9]_net_1\, N_23, 
        \ARB_BYTE[10]_net_1\, N_24, \ARB_BYTE[11]_net_1\, N_31, 
        \ARB_BYTE[12]_net_1\, N_32, \ARB_BYTE[13]_net_1\, N_33, 
        N_34, N_35, N_36, N_37, N_38, N_39, N_40, N_56, 
        \ARB_BYTE[14]_net_1\, N_64, \N_RECD_SER_WORD[0]\, 
        \N_RECD_SER_WORD[1]\, \N_RECD_SER_WORD[2]\, 
        \N_RECD_SER_WORD[3]\, \N_RECD_SER_WORD[4]\, 
        \N_RECD_SER_WORD[5]\, \N_RECD_SER_WORD[6]\, 
        \N_RECD_SER_WORD[7]\, \ADJ_SER_IN_F_0DEL\, 
        \ADJ_SER_IN_R_0DEL\, \ADJ_SER_IN_F_1DEL\, 
        \ADJ_SER_IN_R_1DEL\, \Q[0]_net_1\, \ADJ_Q[0]_net_1\, 
        \Q[1]_net_1\, \ADJ_Q[1]_net_1\, \Q[2]_net_1\, 
        \ADJ_Q[2]_net_1\, \Q[3]_net_1\, \ADJ_Q[3]_net_1\, 
        \Q[4]_net_1\, \ADJ_Q[4]_net_1\, \Q[5]_net_1\, 
        \ADJ_Q[5]_net_1\, \Q[6]_net_1\, \ADJ_Q[6]_net_1\, 
        \Q[7]_net_1\, \ADJ_Q[7]_net_1\, \Q[8]_net_1\, 
        \ADJ_Q[8]_net_1\, \Q[9]_net_1\, \ADJ_Q[9]_net_1\, 
        \Q[10]_net_1\, \ADJ_Q[10]_net_1\, \Q[11]_net_1\, 
        \ADJ_Q[11]_net_1\, \Q[12]_net_1\, \ADJ_Q[12]_net_1\, 
        \Q[13]_net_1\, \ADJ_Q[13]_net_1\, \Q[14]_net_1\, 
        \ADJ_Q[14]_net_1\, \ARB_WRD_40M_FIXED[0]_net_1\, 
        \ARB_WRD_40M_FIXED[1]_net_1\, 
        \ARB_WRD_40M_FIXED[2]_net_1\, 
        \ARB_WRD_40M_FIXED[3]_net_1\, 
        \ARB_WRD_40M_FIXED[4]_net_1\, 
        \ARB_WRD_40M_FIXED[5]_net_1\, 
        \ARB_WRD_40M_FIXED[6]_net_1\, 
        \ARB_WRD_40M_FIXED[7]_net_1\, 
        \ARB_WRD_40M_FIXED[8]_net_1\, 
        \ARB_WRD_40M_FIXED[9]_net_1\, 
        \ARB_WRD_40M_FIXED[10]_net_1\, 
        \ARB_WRD_40M_FIXED[11]_net_1\, 
        \ARB_WRD_40M_FIXED[12]_net_1\, 
        \ARB_WRD_40M_FIXED[13]_net_1\, 
        \ARB_WRD_40M_FIXED[14]_net_1\, \GND\, \VCC\ : std_logic;

begin 


    \ARB_BYTE_RNI5FPV1[2]\ : MX2
      port map(A => N_19, B => N_21, S => BIT_OS_SEL_2(1), Y => 
        N_35);
    
    \RECD_SER_WORD_RNO[5]\ : MX2
      port map(A => N_38, B => N_39, S => BIT_OS_SEL_4_0, Y => 
        \N_RECD_SER_WORD[5]\);
    
    \ARB_WRD_40M_FIXED[9]\ : DFN1C0
      port map(D => \Q[9]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[9]_net_1\);
    
    \ARB_BYTE_RNI09PL[13]\ : MX2
      port map(A => \ARB_BYTE[9]_net_1\, B => 
        \ARB_BYTE[13]_net_1\, S => BIT_OS_SEL_3(2), Y => N_32);
    
    \ADJ_Q[4]\ : DFN1C0
      port map(D => \ADJ_Q[2]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[4]_net_1\);
    
    \ARB_BYTE_RNIAMS02[3]\ : MX2
      port map(A => N_20, B => N_22, S => BIT_OS_SEL_3(1), Y => 
        N_36);
    
    \ARB_BYTE_RNI5IUB1[10]\ : MX2
      port map(A => N_23, B => N_31, S => BIT_OS_SEL_3(1), Y => 
        N_39);
    
    \ARB_BYTE[6]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[6]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[6]_net_1\);
    
    ADJ_SER_IN_F_1DEL : DFN1C0
      port map(D => \ADJ_SER_IN_F_0DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_F_1DEL\);
    
    \ARB_BYTE[0]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[0]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[0]_net_1\);
    
    \Q[11]\ : DFN1C0
      port map(D => \ADJ_Q[11]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[11]_net_1\);
    
    \ADJ_Q[8]\ : DFN1C0
      port map(D => \ADJ_Q[6]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[8]_net_1\);
    
    \ARB_BYTE_RNIP4SL1[11]\ : MX2
      port map(A => N_22, B => N_24, S => BIT_OS_SEL_3(1), Y => 
        N_38);
    
    \ADJ_Q[6]\ : DFN1C0
      port map(D => \ADJ_Q[4]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[6]_net_1\);
    
    \ADJ_Q[12]\ : DFN1C0
      port map(D => \ADJ_Q[10]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[12]_net_1\);
    
    \RECD_SER_WORD_RNO_1[0]\ : MX2
      port map(A => \ARB_BYTE[0]_net_1\, B => \ARB_BYTE[4]_net_1\, 
        S => BIT_OS_SEL_2(2), Y => N_17);
    
    \Q[1]\ : DFN1C0
      port map(D => \ADJ_Q[1]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[1]_net_1\);
    
    \ARB_BYTE_RNICJMV[3]\ : MX2
      port map(A => \ARB_BYTE[3]_net_1\, B => \ARB_BYTE[7]_net_1\, 
        S => BIT_OS_SEL_2(2), Y => N_20);
    
    \ARB_BYTE_RNIPVLK[10]\ : MX2
      port map(A => \ARB_BYTE[6]_net_1\, B => 
        \ARB_BYTE[10]_net_1\, S => BIT_OS_SEL_2(2), Y => N_23);
    
    \ARB_BYTE[4]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[4]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[4]_net_1\);
    
    \ADJ_Q[2]\ : DFN1C0
      port map(D => \ADJ_Q[0]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[2]_net_1\);
    
    \RECD_SER_WORD_RNO_1[7]\ : MX2
      port map(A => \ARB_BYTE[10]_net_1\, B => 
        \ARB_BYTE[14]_net_1\, S => BIT_OS_SEL_5(2), Y => N_56);
    
    \RECD_SER_WORD[4]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[4]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_9(4));
    
    \Q[5]\ : DFN1C0
      port map(D => \ADJ_Q[5]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[5]_net_1\);
    
    \ADJ_Q[11]\ : DFN1C0
      port map(D => \ADJ_Q[9]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[11]_net_1\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \ADJ_Q[3]\ : DFN1C0
      port map(D => \ADJ_Q[1]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[3]_net_1\);
    
    \Q[10]\ : DFN1C0
      port map(D => \ADJ_Q[10]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[10]_net_1\);
    
    \ARB_WRD_40M_FIXED[6]\ : DFN1C0
      port map(D => \Q[6]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[6]_net_1\);
    
    \ARB_WRD_40M_FIXED[1]\ : DFN1C0
      port map(D => \Q[1]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[1]_net_1\);
    
    \RECD_SER_WORD[3]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[3]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_9(3));
    
    \RECD_SER_WORD[0]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[0]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_9(0));
    
    \RECD_SER_WORD_RNO[3]\ : MX2
      port map(A => N_36, B => N_37, S => BIT_OS_SEL_4_0, Y => 
        \N_RECD_SER_WORD[3]\);
    
    \Q[0]\ : DFN1C0
      port map(D => \ADJ_Q[0]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[0]_net_1\);
    
    \ARB_BYTE_RNIELMV[4]\ : MX2
      port map(A => \ARB_BYTE[4]_net_1\, B => \ARB_BYTE[8]_net_1\, 
        S => BIT_OS_SEL_2(2), Y => N_21);
    
    \RECD_SER_WORD_RNO_0[7]\ : MX2
      port map(A => N_31, B => N_56, S => BIT_OS_SEL_5(1), Y => 
        N_64);
    
    \Q[7]\ : DFN1C0
      port map(D => \ADJ_Q[7]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[7]_net_1\);
    
    \ARB_BYTE[14]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[14]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[14]_net_1\);
    
    \ARB_WRD_40M_FIXED[2]\ : DFN1C0
      port map(D => \Q[2]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[2]_net_1\);
    
    \ARB_WRD_40M_FIXED[14]\ : DFN1C0
      port map(D => \Q[14]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[14]_net_1\);
    
    \RECD_SER_WORD_RNO[2]\ : MX2
      port map(A => N_35, B => N_36, S => BIT_OS_SEL_4_0, Y => 
        \N_RECD_SER_WORD[2]\);
    
    \ARB_BYTE[2]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[2]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[2]_net_1\);
    
    \ADJ_Q[7]\ : DFN1C0
      port map(D => \ADJ_Q[5]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[7]_net_1\);
    
    \ARB_BYTE[8]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[8]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[8]_net_1\);
    
    \RECD_SER_WORD[5]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[5]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_9(5));
    
    \ARB_BYTE_RNIL0SL1[10]\ : MX2
      port map(A => N_21, B => N_23, S => BIT_OS_SEL_3(1), Y => 
        N_37);
    
    \ARB_BYTE[12]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[12]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[12]_net_1\);
    
    \RECD_SER_WORD[1]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[1]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_9(1));
    
    \ARB_BYTE_RNI9MUB1[13]\ : MX2
      port map(A => N_24, B => N_32, S => BIT_OS_SEL_3(1), Y => 
        N_40);
    
    \ARB_BYTE_RNIR1MK[11]\ : MX2
      port map(A => \ARB_BYTE[7]_net_1\, B => 
        \ARB_BYTE[11]_net_1\, S => BIT_OS_SEL_2(2), Y => N_24);
    
    \Q[3]\ : DFN1C0
      port map(D => \ADJ_Q[3]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[3]_net_1\);
    
    ADJ_SER_IN_F_0DEL : DFN1C0
      port map(D => ELK_IN_F, CLK => CCC_160M_ADJ, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_F_0DEL\);
    
    \RECD_SER_WORD_RNO[7]\ : MX2
      port map(A => N_40, B => N_64, S => BIT_OS_SEL_4_0, Y => 
        \N_RECD_SER_WORD[7]\);
    
    \RECD_SER_WORD_RNO[1]\ : MX2
      port map(A => N_34, B => N_35, S => BIT_OS_SEL_4_0, Y => 
        \N_RECD_SER_WORD[1]\);
    
    \ARB_WRD_40M_FIXED[4]\ : DFN1C0
      port map(D => \Q[4]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[4]_net_1\);
    
    \RECD_SER_WORD_RNO[0]\ : MX2
      port map(A => N_33, B => N_34, S => BIT_OS_SEL_4_0, Y => 
        \N_RECD_SER_WORD[0]\);
    
    \Q[6]\ : DFN1C0
      port map(D => \ADJ_Q[6]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[6]_net_1\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \ARB_WRD_40M_FIXED[8]\ : DFN1C0
      port map(D => \Q[8]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[8]_net_1\);
    
    \ARB_BYTE[11]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[11]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[11]_net_1\);
    
    \Q[9]\ : DFN1C0
      port map(D => \ADJ_Q[9]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[9]_net_1\);
    
    \ARB_BYTE_RNI1BPV1[1]\ : MX2
      port map(A => N_18, B => N_20, S => BIT_OS_SEL_2(1), Y => 
        N_34);
    
    \Q[14]\ : DFN1C0
      port map(D => \ADJ_Q[14]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[14]_net_1\);
    
    ADJ_SER_IN_R_0DEL : DFN1C0
      port map(D => ELK_IN_R, CLK => CCC_160M_ADJ, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_R_0DEL\);
    
    \Q[13]\ : DFN1C0
      port map(D => \ADJ_Q[13]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[13]_net_1\);
    
    \ARB_BYTE[9]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[9]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[9]_net_1\);
    
    ADJ_SER_IN_R_1DEL : DFN1C0
      port map(D => \ADJ_SER_IN_R_0DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_R_1DEL\);
    
    \ARB_BYTE[10]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[10]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[10]_net_1\);
    
    \ADJ_Q[9]\ : DFN1C0
      port map(D => \ADJ_Q[7]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[9]_net_1\);
    
    \RECD_SER_WORD[7]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[7]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_9(7));
    
    \ARB_WRD_40M_FIXED[5]\ : DFN1C0
      port map(D => \Q[5]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[5]_net_1\);
    
    \ARB_WRD_40M_FIXED[12]\ : DFN1C0
      port map(D => \Q[12]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[12]_net_1\);
    
    \ARB_WRD_40M_FIXED[11]\ : DFN1C0
      port map(D => \Q[11]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[11]_net_1\);
    
    \ARB_WRD_40M_FIXED[0]\ : DFN1C0
      port map(D => \Q[0]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[0]_net_1\);
    
    \ADJ_Q[10]\ : DFN1C0
      port map(D => \ADJ_Q[8]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[10]_net_1\);
    
    \Q[2]\ : DFN1C0
      port map(D => \ADJ_Q[2]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[2]_net_1\);
    
    \ADJ_Q[1]\ : DFN1C0
      port map(D => \ADJ_SER_IN_F_1DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[1]_net_1\);
    
    \RECD_SER_WORD[6]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[6]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_9(6));
    
    \RECD_SER_WORD[2]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[2]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_9(2));
    
    \ADJ_Q[13]\ : DFN1C0
      port map(D => \ADJ_Q[11]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[13]_net_1\);
    
    \ARB_BYTE_RNIU6PL[12]\ : MX2
      port map(A => \ARB_BYTE[8]_net_1\, B => 
        \ARB_BYTE[12]_net_1\, S => BIT_OS_SEL_3(2), Y => N_31);
    
    \Q[8]\ : DFN1C0
      port map(D => \ADJ_Q[8]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[8]_net_1\);
    
    \ARB_BYTE[5]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[5]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[5]_net_1\);
    
    \ADJ_Q[14]\ : DFN1C0
      port map(D => \ADJ_Q[12]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[14]_net_1\);
    
    \RECD_SER_WORD_RNO[4]\ : MX2
      port map(A => N_37, B => N_38, S => BIT_OS_SEL_4_0, Y => 
        \N_RECD_SER_WORD[4]\);
    
    \Q[12]\ : DFN1C0
      port map(D => \ADJ_Q[12]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[12]_net_1\);
    
    \ARB_BYTE[13]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[13]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[13]_net_1\);
    
    \ARB_BYTE_RNIGNMV[5]\ : MX2
      port map(A => \ARB_BYTE[5]_net_1\, B => \ARB_BYTE[9]_net_1\, 
        S => BIT_OS_SEL_2(2), Y => N_22);
    
    \ARB_WRD_40M_FIXED[3]\ : DFN1C0
      port map(D => \Q[3]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[3]_net_1\);
    
    \ARB_BYTE_RNI8FMV[1]\ : MX2
      port map(A => \ARB_BYTE[1]_net_1\, B => \ARB_BYTE[5]_net_1\, 
        S => BIT_OS_SEL_2(2), Y => N_18);
    
    \ARB_BYTE[7]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[7]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[7]_net_1\);
    
    \RECD_SER_WORD_RNO_0[0]\ : MX2
      port map(A => N_17, B => N_19, S => BIT_OS_SEL_2(1), Y => 
        N_33);
    
    \Q[4]\ : DFN1C0
      port map(D => \ADJ_Q[4]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[4]_net_1\);
    
    \ARB_WRD_40M_FIXED[7]\ : DFN1C0
      port map(D => \Q[7]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[7]_net_1\);
    
    \RECD_SER_WORD_RNO[6]\ : MX2
      port map(A => N_39, B => N_40, S => BIT_OS_SEL_4_0, Y => 
        \N_RECD_SER_WORD[6]\);
    
    \ARB_BYTE[3]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[3]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[3]_net_1\);
    
    \ADJ_Q[5]\ : DFN1C0
      port map(D => \ADJ_Q[3]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[5]_net_1\);
    
    \ARB_BYTE[1]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[1]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[1]_net_1\);
    
    \ARB_WRD_40M_FIXED[13]\ : DFN1C0
      port map(D => \Q[13]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[13]_net_1\);
    
    \ARB_BYTE_RNIAHMV[2]\ : MX2
      port map(A => \ARB_BYTE[2]_net_1\, B => \ARB_BYTE[6]_net_1\, 
        S => BIT_OS_SEL_2(2), Y => N_19);
    
    \ADJ_Q[0]\ : DFN1C0
      port map(D => \ADJ_SER_IN_R_1DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[0]_net_1\);
    
    \ARB_WRD_40M_FIXED[10]\ : DFN1C0
      port map(D => \Q[10]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[10]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SER320M_3_34_9 is

    port( ELK_TX_DAT                 : in    std_logic_vector(7 downto 0);
          MASTER_SALT_POR_B_i_0_i_0  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_4  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_3  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_2  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_13 : in    std_logic;
          ELK_OUT_R                  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_16 : in    std_logic;
          ELK_OUT_F                  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_12 : in    std_logic;
          CCC_160M_FXD               : in    std_logic;
          CLK_40M_GL                 : in    std_logic
        );

end SER320M_3_34_9;

architecture DEF_ARCH of SER320M_3_34_9 is 

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \N_SER_CMD_WORD_R[0]\, \START_RISE\, 
        \N_SER_CMD_WORD_F[0]\, \N_SER_CMD_WORD_R[3]\, 
        \SER_CMD_WORD_R[2]_net_1\, \N_SER_CMD_WORD_R[2]\, 
        \SER_CMD_WORD_R[1]_net_1\, \N_SER_CMD_WORD_R[1]\, 
        \SER_CMD_WORD_R[0]_net_1\, \N_SER_CMD_WORD_F[3]\, 
        \SER_CMD_WORD_F[2]_net_1\, \N_SER_CMD_WORD_F[2]\, 
        \SER_CMD_WORD_F[1]_net_1\, \N_SER_CMD_WORD_F[1]\, 
        \SER_CMD_WORD_F[0]_net_1\, N_START_RISE, 
        \CLK40M_GEN_DEL0\, \SER_OUT_FI\, \SER_OUT_RI\, 
        \SER_CMD_WORD_F[3]_net_1\, \SER_CMD_WORD_R[3]_net_1\, 
        \GND\, \VCC\ : std_logic;

begin 


    SER_OUT_FI : DFN1C0
      port map(D => \SER_CMD_WORD_F[3]_net_1\, CLK => 
        CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_12, Q => 
        \SER_OUT_FI\);
    
    \SER_CMD_WORD_F[3]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[3]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_4, Q => 
        \SER_CMD_WORD_F[3]_net_1\);
    
    \SER_CMD_WORD_R[1]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[1]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_0, Q => 
        \SER_CMD_WORD_R[1]_net_1\);
    
    \SER_CMD_WORD_R[2]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[2]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_0, Q => 
        \SER_CMD_WORD_R[2]_net_1\);
    
    \SER_CMD_WORD_R_RNO[3]\ : MX2
      port map(A => \SER_CMD_WORD_R[2]_net_1\, B => ELK_TX_DAT(7), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_R[3]\);
    
    \SER_CMD_WORD_R_RNO[0]\ : NOR2B
      port map(A => \START_RISE\, B => ELK_TX_DAT(1), Y => 
        \N_SER_CMD_WORD_R[0]\);
    
    \SER_CMD_WORD_F[0]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[0]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_3, Q => 
        \SER_CMD_WORD_F[0]_net_1\);
    
    \SER_CMD_WORD_R_RNO[1]\ : MX2
      port map(A => \SER_CMD_WORD_R[0]_net_1\, B => ELK_TX_DAT(3), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_R[1]\);
    
    \SER_CMD_WORD_F_RNO[2]\ : MX2
      port map(A => \SER_CMD_WORD_F[1]_net_1\, B => ELK_TX_DAT(4), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_F[2]\);
    
    \SER_CMD_WORD_F_RNO[3]\ : MX2
      port map(A => \SER_CMD_WORD_F[2]_net_1\, B => ELK_TX_DAT(6), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_F[3]\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    CLK40M_GEN_DEL0 : DFN1C0
      port map(D => CLK_40M_GL, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_12, Q => \CLK40M_GEN_DEL0\);
    
    SER_OUT_RI : DFN1C0
      port map(D => \SER_CMD_WORD_R[3]_net_1\, CLK => 
        CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_13, Q => 
        \SER_OUT_RI\);
    
    \SER_CMD_WORD_F[2]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[2]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_4, Q => 
        \SER_CMD_WORD_F[2]_net_1\);
    
    \SER_CMD_WORD_F_RNO[1]\ : MX2
      port map(A => \SER_CMD_WORD_F[0]_net_1\, B => ELK_TX_DAT(2), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_F[1]\);
    
    \SER_CMD_WORD_R[0]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[0]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_0, Q => 
        \SER_CMD_WORD_R[0]_net_1\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    START_RISE : DFN1C0
      port map(D => N_START_RISE, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_2, Q => \START_RISE\);
    
    \SER_CMD_WORD_R[3]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[3]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_0, Q => 
        \SER_CMD_WORD_R[3]_net_1\);
    
    \SER_CMD_WORD_F_RNO[0]\ : NOR2B
      port map(A => \START_RISE\, B => ELK_TX_DAT(0), Y => 
        \N_SER_CMD_WORD_F[0]\);
    
    SER_OUT_RDEL : DFN1C0
      port map(D => \SER_OUT_RI\, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_13, Q => ELK_OUT_R);
    
    \SER_CMD_WORD_F[1]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[1]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_4, Q => 
        \SER_CMD_WORD_F[1]_net_1\);
    
    START_RISE_RNO : NOR2B
      port map(A => \CLK40M_GEN_DEL0\, B => CLK_40M_GL, Y => 
        N_START_RISE);
    
    \SER_CMD_WORD_R_RNO[2]\ : MX2
      port map(A => \SER_CMD_WORD_R[1]_net_1\, B => ELK_TX_DAT(5), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_R[2]\);
    
    SER_OUT_FDEL : DFN1C0
      port map(D => \SER_OUT_FI\, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_16, Q => ELK_OUT_F);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity DDR_BIDIR_LVDS_DUAL_CLK_9 is

    port( DCB_SALT_SEL_c_i : in    std_logic;
          ELK9_DAT_P       : inout std_logic := 'Z';
          ELK9_DAT_N       : inout std_logic := 'Z';
          ELK_OUT_R        : in    std_logic;
          ELK_OUT_F        : in    std_logic;
          CCC_160M_FXD     : in    std_logic;
          CCC_160M_ADJ     : in    std_logic;
          ELK_IN_DDR_R     : out   std_logic;
          ELK_IN_DDR_F     : out   std_logic
        );

end DDR_BIDIR_LVDS_DUAL_CLK_9;

architecture DEF_ARCH of DDR_BIDIR_LVDS_DUAL_CLK_9 is 

  component DDR_REG
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          QR  : out   std_logic;
          QF  : out   std_logic
        );
  end component;

  component DDR_OUT
    port( DR  : in    std_logic := 'U';
          DF  : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component BIBUF_LVDS
    port( PADP : inout   std_logic;
          PADN : inout   std_logic;
          D    : in    std_logic := 'U';
          E    : in    std_logic := 'U';
          Y    : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal DDR_BIDIR_LVDS_DUAL_CLK_9_GND, BIBUF_LVDS_0_Y, 
        DDR_OUT_0_Q, \VCC\ : std_logic;

begin 


    DDR_REG_0 : DDR_REG
      port map(D => BIBUF_LVDS_0_Y, CLK => CCC_160M_ADJ, CLR => 
        DDR_BIDIR_LVDS_DUAL_CLK_9_GND, QR => ELK_IN_DDR_R, QF => 
        ELK_IN_DDR_F);
    
    DDR_OUT_0 : DDR_OUT
      port map(DR => ELK_OUT_R, DF => ELK_OUT_F, CLK => 
        CCC_160M_FXD, CLR => DDR_BIDIR_LVDS_DUAL_CLK_9_GND, Q => 
        DDR_OUT_0_Q);
    
    BIBUF_LVDS_0 : BIBUF_LVDS
      port map(PADP => ELK9_DAT_P, PADN => ELK9_DAT_N, D => 
        DDR_OUT_0_Q, E => DCB_SALT_SEL_c_i, Y => BIBUF_LVDS_0_Y);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    GND_i : GND
      port map(Y => DDR_BIDIR_LVDS_DUAL_CLK_9_GND);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SYNC_DAT_SEL_9 is

    port( ELK_TX_DAT                : out   std_logic_vector(7 downto 0);
          PATT_ELK_DAT_9            : in    std_logic_vector(7 downto 0);
          OP_MODE_c_3_0             : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_7 : in    std_logic;
          CLK_40M_GL                : in    std_logic
        );

end SYNC_DAT_SEL_9;

architecture DEF_ARCH of SYNC_DAT_SEL_9 is 

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \N_SERDAT[0]\, \N_SERDAT[1]\, \N_SERDAT[2]\, 
        \N_SERDAT[3]\, \N_SERDAT[4]\, \N_SERDAT[5]\, 
        \N_SERDAT[6]\, \N_SERDAT[7]\, \GND\, \VCC\ : std_logic;

begin 


    \SERDAT_RNO[4]\ : NOR2A
      port map(A => PATT_ELK_DAT_9(4), B => OP_MODE_c_3_0, Y => 
        \N_SERDAT[4]\);
    
    \SERDAT_RNO[0]\ : NOR2A
      port map(A => PATT_ELK_DAT_9(0), B => OP_MODE_c_3_0, Y => 
        \N_SERDAT[0]\);
    
    \SERDAT[6]\ : DFN1C0
      port map(D => \N_SERDAT[6]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_7, Q => ELK_TX_DAT(6));
    
    \SERDAT[4]\ : DFN1C0
      port map(D => \N_SERDAT[4]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_7, Q => ELK_TX_DAT(4));
    
    \SERDAT_RNO[7]\ : OR2
      port map(A => PATT_ELK_DAT_9(7), B => OP_MODE_c_3_0, Y => 
        \N_SERDAT[7]\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \SERDAT_RNO[3]\ : OR2
      port map(A => PATT_ELK_DAT_9(3), B => OP_MODE_c_3_0, Y => 
        \N_SERDAT[3]\);
    
    \SERDAT_RNO[2]\ : OR2
      port map(A => PATT_ELK_DAT_9(2), B => OP_MODE_c_3_0, Y => 
        \N_SERDAT[2]\);
    
    \SERDAT[5]\ : DFN1C0
      port map(D => \N_SERDAT[5]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_7, Q => ELK_TX_DAT(5));
    
    \SERDAT[7]\ : DFN1C0
      port map(D => \N_SERDAT[7]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_7, Q => ELK_TX_DAT(7));
    
    GND_i : GND
      port map(Y => \GND\);
    
    \SERDAT_RNO[5]\ : NOR2A
      port map(A => PATT_ELK_DAT_9(5), B => OP_MODE_c_3_0, Y => 
        \N_SERDAT[5]\);
    
    \SERDAT[0]\ : DFN1C0
      port map(D => \N_SERDAT[0]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_7, Q => ELK_TX_DAT(0));
    
    \SERDAT_RNO[6]\ : NOR2A
      port map(A => PATT_ELK_DAT_9(6), B => OP_MODE_c_3_0, Y => 
        \N_SERDAT[6]\);
    
    \SERDAT[1]\ : DFN1C0
      port map(D => \N_SERDAT[1]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_7, Q => ELK_TX_DAT(1));
    
    \SERDAT_RNO[1]\ : OR2
      port map(A => PATT_ELK_DAT_9(1), B => OP_MODE_c_3_0, Y => 
        \N_SERDAT[1]\);
    
    \SERDAT[3]\ : DFN1C0
      port map(D => \N_SERDAT[3]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_7, Q => ELK_TX_DAT(3));
    
    \SERDAT[2]\ : DFN1C0
      port map(D => \N_SERDAT[2]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_7, Q => ELK_TX_DAT(2));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity ELINK_SLAVE_15_4 is

    port( BIT_OS_SEL_2               : in    std_logic_vector(2 downto 1);
          BIT_OS_SEL_3               : in    std_logic_vector(2 downto 1);
          BIT_OS_SEL_5               : in    std_logic_vector(2 downto 1);
          BIT_OS_SEL_4_0             : in    std_logic;
          ELK_RX_SER_WORD_9          : out   std_logic_vector(7 downto 0);
          OP_MODE_c_3_0              : in    std_logic;
          PATT_ELK_DAT_9             : in    std_logic_vector(7 downto 0);
          MASTER_DCB_POR_B_i_0_i     : in    std_logic;
          ELK9_DAT_N                 : inout std_logic := 'Z';
          ELK9_DAT_P                 : inout std_logic := 'Z';
          DCB_SALT_SEL_c_i           : in    std_logic;
          CCC_160M_FXD               : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_12 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_16 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_13 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_2  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_3  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_4  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_0  : in    std_logic;
          CLK_40M_GL                 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_7  : in    std_logic;
          DEV_RST_B_c_0              : in    std_logic;
          CCC_160M_ADJ               : in    std_logic
        );

end ELINK_SLAVE_15_4;

architecture DEF_ARCH of ELINK_SLAVE_15_4 is 

  component SLAVE_DES320S_1_17_7
    port( ELK_RX_SER_WORD_9      : out   std_logic_vector(7 downto 0);
          BIT_OS_SEL_4_0         : in    std_logic := 'U';
          BIT_OS_SEL_5           : in    std_logic_vector(2 downto 1) := (others => 'U');
          BIT_OS_SEL_3           : in    std_logic_vector(2 downto 1) := (others => 'U');
          BIT_OS_SEL_2           : in    std_logic_vector(2 downto 1) := (others => 'U');
          CLK_40M_GL             : in    std_logic := 'U';
          CCC_160M_FXD           : in    std_logic := 'U';
          ELK_IN_R               : in    std_logic := 'U';
          ELK_IN_F               : in    std_logic := 'U';
          MASTER_DCB_POR_B_i_0_i : in    std_logic := 'U';
          CCC_160M_ADJ           : in    std_logic := 'U'
        );
  end component;

  component SER320M_3_34_9
    port( ELK_TX_DAT                 : in    std_logic_vector(7 downto 0) := (others => 'U');
          MASTER_SALT_POR_B_i_0_i_0  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_4  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_3  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_2  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_13 : in    std_logic := 'U';
          ELK_OUT_R                  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_16 : in    std_logic := 'U';
          ELK_OUT_F                  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_12 : in    std_logic := 'U';
          CCC_160M_FXD               : in    std_logic := 'U';
          CLK_40M_GL                 : in    std_logic := 'U'
        );
  end component;

  component DDR_BIDIR_LVDS_DUAL_CLK_9
    port( DCB_SALT_SEL_c_i : in    std_logic := 'U';
          ELK9_DAT_P       : inout   std_logic;
          ELK9_DAT_N       : inout   std_logic;
          ELK_OUT_R        : in    std_logic := 'U';
          ELK_OUT_F        : in    std_logic := 'U';
          CCC_160M_FXD     : in    std_logic := 'U';
          CCC_160M_ADJ     : in    std_logic := 'U';
          ELK_IN_DDR_R     : out   std_logic;
          ELK_IN_DDR_F     : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component SYNC_DAT_SEL_9
    port( ELK_TX_DAT                : out   std_logic_vector(7 downto 0);
          PATT_ELK_DAT_9            : in    std_logic_vector(7 downto 0) := (others => 'U');
          OP_MODE_c_3_0             : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_7 : in    std_logic := 'U';
          CLK_40M_GL                : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \ELK_IN_F\, ELK_IN_DDR_F, \ELK_IN_R\, ELK_IN_DDR_R, 
        \ELK_TX_DAT[0]\, \ELK_TX_DAT[1]\, \ELK_TX_DAT[2]\, 
        \ELK_TX_DAT[3]\, \ELK_TX_DAT[4]\, \ELK_TX_DAT[5]\, 
        \ELK_TX_DAT[6]\, \ELK_TX_DAT[7]\, ELK_OUT_R, ELK_OUT_F, 
        \GND\, \VCC\ : std_logic;

    for all : SLAVE_DES320S_1_17_7
	Use entity work.SLAVE_DES320S_1_17_7(DEF_ARCH);
    for all : SER320M_3_34_9
	Use entity work.SER320M_3_34_9(DEF_ARCH);
    for all : DDR_BIDIR_LVDS_DUAL_CLK_9
	Use entity work.DDR_BIDIR_LVDS_DUAL_CLK_9(DEF_ARCH);
    for all : SYNC_DAT_SEL_9
	Use entity work.SYNC_DAT_SEL_9(DEF_ARCH);
begin 


    U_SLAVE_1ELK : SLAVE_DES320S_1_17_7
      port map(ELK_RX_SER_WORD_9(7) => ELK_RX_SER_WORD_9(7), 
        ELK_RX_SER_WORD_9(6) => ELK_RX_SER_WORD_9(6), 
        ELK_RX_SER_WORD_9(5) => ELK_RX_SER_WORD_9(5), 
        ELK_RX_SER_WORD_9(4) => ELK_RX_SER_WORD_9(4), 
        ELK_RX_SER_WORD_9(3) => ELK_RX_SER_WORD_9(3), 
        ELK_RX_SER_WORD_9(2) => ELK_RX_SER_WORD_9(2), 
        ELK_RX_SER_WORD_9(1) => ELK_RX_SER_WORD_9(1), 
        ELK_RX_SER_WORD_9(0) => ELK_RX_SER_WORD_9(0), 
        BIT_OS_SEL_4_0 => BIT_OS_SEL_4_0, BIT_OS_SEL_5(2) => 
        BIT_OS_SEL_5(2), BIT_OS_SEL_5(1) => BIT_OS_SEL_5(1), 
        BIT_OS_SEL_3(2) => BIT_OS_SEL_3(2), BIT_OS_SEL_3(1) => 
        BIT_OS_SEL_3(1), BIT_OS_SEL_2(2) => BIT_OS_SEL_2(2), 
        BIT_OS_SEL_2(1) => BIT_OS_SEL_2(1), CLK_40M_GL => 
        CLK_40M_GL, CCC_160M_FXD => CCC_160M_FXD, ELK_IN_R => 
        \ELK_IN_R\, ELK_IN_F => \ELK_IN_F\, 
        MASTER_DCB_POR_B_i_0_i => MASTER_DCB_POR_B_i_0_i, 
        CCC_160M_ADJ => CCC_160M_ADJ);
    
    U_ELK1_CMD_TX : SER320M_3_34_9
      port map(ELK_TX_DAT(7) => \ELK_TX_DAT[7]\, ELK_TX_DAT(6)
         => \ELK_TX_DAT[6]\, ELK_TX_DAT(5) => \ELK_TX_DAT[5]\, 
        ELK_TX_DAT(4) => \ELK_TX_DAT[4]\, ELK_TX_DAT(3) => 
        \ELK_TX_DAT[3]\, ELK_TX_DAT(2) => \ELK_TX_DAT[2]\, 
        ELK_TX_DAT(1) => \ELK_TX_DAT[1]\, ELK_TX_DAT(0) => 
        \ELK_TX_DAT[0]\, MASTER_SALT_POR_B_i_0_i_0 => 
        MASTER_SALT_POR_B_i_0_i_0, MASTER_SALT_POR_B_i_0_i_4 => 
        MASTER_SALT_POR_B_i_0_i_4, MASTER_SALT_POR_B_i_0_i_3 => 
        MASTER_SALT_POR_B_i_0_i_3, MASTER_SALT_POR_B_i_0_i_2 => 
        MASTER_SALT_POR_B_i_0_i_2, MASTER_SALT_POR_B_i_0_i_13 => 
        MASTER_SALT_POR_B_i_0_i_13, ELK_OUT_R => ELK_OUT_R, 
        MASTER_SALT_POR_B_i_0_i_16 => MASTER_SALT_POR_B_i_0_i_16, 
        ELK_OUT_F => ELK_OUT_F, MASTER_SALT_POR_B_i_0_i_12 => 
        MASTER_SALT_POR_B_i_0_i_12, CCC_160M_FXD => CCC_160M_FXD, 
        CLK_40M_GL => CLK_40M_GL);
    
    U_DDR_ELK1 : DDR_BIDIR_LVDS_DUAL_CLK_9
      port map(DCB_SALT_SEL_c_i => DCB_SALT_SEL_c_i, ELK9_DAT_P
         => ELK9_DAT_P, ELK9_DAT_N => ELK9_DAT_N, ELK_OUT_R => 
        ELK_OUT_R, ELK_OUT_F => ELK_OUT_F, CCC_160M_FXD => 
        CCC_160M_FXD, CCC_160M_ADJ => CCC_160M_ADJ, ELK_IN_DDR_R
         => ELK_IN_DDR_R, ELK_IN_DDR_F => ELK_IN_DDR_F);
    
    ELK_IN_F : DFN1C0
      port map(D => ELK_IN_DDR_F, CLK => CCC_160M_ADJ, CLR => 
        DEV_RST_B_c_0, Q => \ELK_IN_F\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    U_ELK1_SERDAT_SOURCE : SYNC_DAT_SEL_9
      port map(ELK_TX_DAT(7) => \ELK_TX_DAT[7]\, ELK_TX_DAT(6)
         => \ELK_TX_DAT[6]\, ELK_TX_DAT(5) => \ELK_TX_DAT[5]\, 
        ELK_TX_DAT(4) => \ELK_TX_DAT[4]\, ELK_TX_DAT(3) => 
        \ELK_TX_DAT[3]\, ELK_TX_DAT(2) => \ELK_TX_DAT[2]\, 
        ELK_TX_DAT(1) => \ELK_TX_DAT[1]\, ELK_TX_DAT(0) => 
        \ELK_TX_DAT[0]\, PATT_ELK_DAT_9(7) => PATT_ELK_DAT_9(7), 
        PATT_ELK_DAT_9(6) => PATT_ELK_DAT_9(6), PATT_ELK_DAT_9(5)
         => PATT_ELK_DAT_9(5), PATT_ELK_DAT_9(4) => 
        PATT_ELK_DAT_9(4), PATT_ELK_DAT_9(3) => PATT_ELK_DAT_9(3), 
        PATT_ELK_DAT_9(2) => PATT_ELK_DAT_9(2), PATT_ELK_DAT_9(1)
         => PATT_ELK_DAT_9(1), PATT_ELK_DAT_9(0) => 
        PATT_ELK_DAT_9(0), OP_MODE_c_3_0 => OP_MODE_c_3_0, 
        MASTER_SALT_POR_B_i_0_i_7 => MASTER_SALT_POR_B_i_0_i_7, 
        CLK_40M_GL => CLK_40M_GL);
    
    ELK_IN_R : DFN1C0
      port map(D => ELK_IN_DDR_R, CLK => CCC_160M_ADJ, CLR => 
        DEV_RST_B_c_0, Q => \ELK_IN_R\);
    
    GND_i : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity GP_PATT_GEN_1 is

    port( TFC_ADDRB              : out   std_logic_vector(7 downto 0);
          TFC_RX_SER_WORD        : in    std_logic_vector(7 downto 0);
          TFC_STOP_ADDR          : in    std_logic_vector(7 downto 0);
          TFC_STRT_ADDR          : in    std_logic_vector(7 downto 0);
          OP_MODE_0              : in    std_logic;
          OP_MODE_c_0            : in    std_logic;
          P_MASTER_POR_B_c_24    : in    std_logic;
          P_MASTER_POR_B_c       : in    std_logic;
          P_MASTER_POR_B_c_31    : in    std_logic;
          P_MASTER_POR_B_c_30    : in    std_logic;
          P_MASTER_POR_B_c_1     : in    std_logic;
          P_MASTER_POR_B_c_5     : in    std_logic;
          P_MASTER_POR_B_c_4     : in    std_logic;
          P_MASTER_POR_B_c_28    : in    std_logic;
          DCB_SALT_SEL_c         : in    std_logic;
          P_MASTER_POR_B_c_15    : in    std_logic;
          P_MASTER_POR_B_c_16_0  : in    std_logic;
          TFC_RWB                : out   std_logic;
          P_MASTER_POR_B_c_9     : in    std_logic;
          TFC_RAM_BLKB_EN        : out   std_logic;
          P_USB_MASTER_EN_c_22_0 : in    std_logic;
          ALIGN_ACTIVE           : in    std_logic;
          P_MASTER_POR_B_c_27_1  : in    std_logic;
          CLK_40M_GL             : in    std_logic
        );

end GP_PATT_GEN_1;

architecture DEF_ARCH of GP_PATT_GEN_1 is 

  component OA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component DFN1E1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E0P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component INV
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XNOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component AO1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component OA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

    signal \GP_PG_SM_0[10]_net_1\, \GP_PG_SM_ns[0]\, 
        \DWACT_ADD_CI_0_g_array_11[0]\, 
        \DWACT_ADD_CI_0_g_array_2[0]\, 
        \DWACT_ADD_CI_0_pog_array_1_1[0]\, 
        \DWACT_ADD_CI_0_g_array_1[0]\, 
        \DWACT_ADD_CI_0_pog_array_1[0]\, \DWACT_ADD_CI_0_TMP[0]\, 
        \TFC_ADDRB[1]\, \DWACT_ADD_CI_0_g_array_12_1[0]\, 
        \TFC_ADDRB[4]\, \DWACT_ADD_CI_0_g_array_12_2[0]\, 
        \TFC_ADDRB[6]\, \DWACT_ADD_CI_0_g_array_12[0]\, 
        \TFC_ADDRB[2]\, \RX_SER_WORD_2DEL_i[1]\, 
        \RX_SER_WORD_2DEL[1]_net_1\, \RX_SER_WORD_2DEL_i[2]\, 
        \RX_SER_WORD_2DEL[2]_net_1\, \RX_SER_WORD_2DEL_i[3]\, 
        \RX_SER_WORD_2DEL[3]_net_1\, \RX_SER_WORD_2DEL_i[7]\, 
        \RX_SER_WORD_2DEL[7]_net_1\, \N_ADDR_POINTER_i_o2_0[7]\, 
        N_39, N_214_li, \GP_PG_SM[10]_net_1\, 
        \GP_PG_SM_ns_0_a2_0[5]\, \GP_PG_SM[5]_net_1\, 
        \GP_PG_SM[4]_net_1\, \GP_PG_SM_ns_i_i_a4_0[7]\, 
        \GP_PG_SM[3]_net_1\, \GP_PG_SM[2]_net_1\, 
        \GP_PG_SM_ns_i_i_a4_1[1]\, \GP_PG_SM[9]_net_1\, N_45, 
        \GP_PG_SM_ns_i_i_a4_0_1[7]\, \GP_PG_SM[8]_net_1\, N_114, 
        \GP_PG_SM_ns_i_i_a4_0[2]\, N_213_li, 
        \GP_PG_SM_ns_0_a4_1[0]\, N_315, \GP_PG_SM[1]_net_1\, 
        \GP_PG_SM_ns_0_a2_0_1[5]\, \GP_PG_SM_ns_0_a4_0[6]\, 
        \GP_PG_SM[6]_net_1\, un1_RX_SER_WORD_2DEL_NE_4, 
        \RX_SER_WORD_2DEL[5]_net_1\, \RX_SER_WORD_2DEL[4]_net_1\, 
        un1_RX_SER_WORD_2DEL_NE_1, un1_RX_SER_WORD_2DEL_NE_3, 
        un1_RX_SER_WORD_2DEL_NE_2, \RX_SER_WORD_2DEL[0]_net_1\, 
        \RX_SER_WORD_2DEL[6]_net_1\, un1_RX_SER_WORD_3DEL_NE_4, 
        \RX_SER_WORD_3DEL[5]_net_1\, \RX_SER_WORD_3DEL[4]_net_1\, 
        un1_RX_SER_WORD_3DEL_NE_1, un1_RX_SER_WORD_3DEL_NE_3, 
        \RX_SER_WORD_3DEL_i_0[2]\, \RX_SER_WORD_3DEL_i_0[3]\, 
        un1_RX_SER_WORD_3DEL_NE_2, \RX_SER_WORD_3DEL[0]_net_1\, 
        \RX_SER_WORD_3DEL_i_0[1]\, \RX_SER_WORD_3DEL[6]_net_1\, 
        \RX_SER_WORD_3DEL_i_0[7]\, un1_RX_SER_WORD_3DEL_1, 
        un1_RX_SER_WORD_2DEL_1, N_38, N_105, N_106, N_104, N_36, 
        N_102, N_103, N_101, N_34, N_382, N_383, N_381, N_30, 
        N_375, N_377, N_376, N_26, N_86, N_88, N_87, N_24, N_83, 
        N_85, N_84, N_107, N_40, \GP_PG_SM_RNO[1]_net_1\, N_73, 
        N_61, N_42, N_69, N_116, N_71, N_50, N_110, N_80, N_160_3, 
        N_28, N_89, N_374, N_373, N_32, N_378, N_380, N_379, N_76, 
        N_47, N_22, N_210_li, \GP_PG_SM[7]_net_1\, N_18, N_117, 
        N_64, \GP_PG_SM_ns_0_a2_0_1[3]\, \GP_PG_SM_ns[3]\, 
        \GP_PG_SM_ns_0_a2_0[3]\, N_25, I_34, 
        \LOC_STRT_ADDR[7]_net_1\, I_31, \LOC_STRT_ADDR[6]_net_1\, 
        I_33, \LOC_STRT_ADDR[4]_net_1\, I_29, 
        \LOC_STRT_ADDR[2]_net_1\, I_30, \LOC_STRT_ADDR[1]_net_1\, 
        \DWACT_ADD_CI_0_partial_sum[0]\, \LOC_STRT_ADDR[0]_net_1\, 
        \GP_PG_SM[0]_net_1\, \GP_PG_SM_ns[10]\, 
        \GP_PG_SM_RNITIQ71[10]_net_1\, \GP_PG_SM_ns[5]\, N_65, 
        \GP_PG_SM_ns[6]\, N_79, \GP_PG_SM_RNO[3]_net_1\, 
        \GP_PG_SM_RNO[2]_net_1\, N_74, \LOC_STRT_ADDR[3]_net_1\, 
        I_27, \LOC_STRT_ADDR[5]_net_1\, I_28, N_238, 
        \LOC_STOP_ADDR[0]_net_1\, \LOC_STOP_ADDR[1]_net_1\, 
        \LOC_STOP_ADDR[2]_net_1\, \LOC_STOP_ADDR[3]_net_1\, 
        \LOC_STOP_ADDR[4]_net_1\, \LOC_STOP_ADDR[5]_net_1\, 
        \LOC_STOP_ADDR[6]_net_1\, \LOC_STOP_ADDR[7]_net_1\, 
        \RX_SER_WORD_1DEL[0]_net_1\, \RX_SER_WORD_1DEL[1]_net_1\, 
        \RX_SER_WORD_1DEL[2]_net_1\, \RX_SER_WORD_1DEL[3]_net_1\, 
        \RX_SER_WORD_1DEL[4]_net_1\, \RX_SER_WORD_1DEL[5]_net_1\, 
        \RX_SER_WORD_1DEL[6]_net_1\, \RX_SER_WORD_1DEL[7]_net_1\, 
        \TFC_ADDRB[0]\, \TFC_ADDRB[3]\, \TFC_ADDRB[5]\, 
        \TFC_ADDRB[7]\, \DWACT_COMP0_E[1]\, \DWACT_COMP0_E[2]\, 
        \DWACT_COMP0_E[0]\, N_11, N_10, N_9, N_6, N_8, N_7, N_5, 
        N_2, N_3, N_4, \ACT_LT3_E[3]\, \ACT_LT3_E[4]\, 
        \ACT_LT3_E[5]\, \ACT_LT3_E[0]\, \ACT_LT3_E[1]\, 
        \ACT_LT3_E[2]\, \DWACT_BL_EQUAL_0_E[2]\, 
        \DWACT_BL_EQUAL_0_E[1]\, \DWACT_BL_EQUAL_0_E[0]\, \GND\, 
        \VCC\ : std_logic;

begin 

    TFC_ADDRB(7) <= \TFC_ADDRB[7]\;
    TFC_ADDRB(6) <= \TFC_ADDRB[6]\;
    TFC_ADDRB(5) <= \TFC_ADDRB[5]\;
    TFC_ADDRB(4) <= \TFC_ADDRB[4]\;
    TFC_ADDRB(3) <= \TFC_ADDRB[3]\;
    TFC_ADDRB(2) <= \TFC_ADDRB[2]\;
    TFC_ADDRB(1) <= \TFC_ADDRB[1]\;
    TFC_ADDRB(0) <= \TFC_ADDRB[0]\;

    \ADDR_POINTER_RNO_2[1]\ : OA1B
      port map(A => N_107, B => \N_ADDR_POINTER_i_o2_0[7]\, C => 
        TFC_STRT_ADDR(1), Y => N_101);
    
    un1_ADDR_POINTER_2_I_46 : AND2
      port map(A => \TFC_ADDRB[2]\, B => \TFC_ADDRB[3]\, Y => 
        \DWACT_ADD_CI_0_pog_array_1[0]\);
    
    \GP_PG.un1_ADDR_POINTER_0_I_25\ : AO1
      port map(A => \DWACT_COMP0_E[1]\, B => \DWACT_COMP0_E[2]\, 
        C => \DWACT_COMP0_E[0]\, Y => N_214_li);
    
    \GP_PG_SM_RNO_0[8]\ : NOR2B
      port map(A => \GP_PG_SM[9]_net_1\, B => N_213_li, Y => 
        \GP_PG_SM_ns_i_i_a4_0[2]\);
    
    \GP_PG_SM_RNIP30G[6]\ : NOR2
      port map(A => \GP_PG_SM[6]_net_1\, B => \GP_PG_SM[7]_net_1\, 
        Y => N_114);
    
    \ADDR_POINTER_RNO_0[4]\ : OA1B
      port map(A => N_107, B => \N_ADDR_POINTER_i_o2_0[7]\, C => 
        TFC_STRT_ADDR(4), Y => N_375);
    
    un1_ADDR_POINTER_2_I_45 : NOR2B
      port map(A => \DWACT_ADD_CI_0_g_array_1[0]\, B => 
        \TFC_ADDRB[2]\, Y => \DWACT_ADD_CI_0_g_array_12[0]\);
    
    \GP_PG_SM_RNO_1[4]\ : NOR3C
      port map(A => N_214_li, B => N_117, C => 
        \GP_PG_SM[4]_net_1\, Y => N_79);
    
    \ADDR_POINTER[2]\ : DFN1C0
      port map(D => N_34, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_30, Q => \TFC_ADDRB[2]\);
    
    \RX_SER_WORD_1DEL[7]\ : DFN1C0
      port map(D => TFC_RX_SER_WORD(7), CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_31, Q => \RX_SER_WORD_1DEL[7]_net_1\);
    
    \ADDR_POINTER_RNO_0[6]\ : OA1B
      port map(A => N_107, B => \N_ADDR_POINTER_i_o2_0[7]\, C => 
        TFC_STRT_ADDR(6), Y => N_86);
    
    \GP_PG.un1_ADDR_POINTER_0_I_21\ : OR2A
      port map(A => \TFC_ADDRB[4]\, B => \LOC_STOP_ADDR[4]_net_1\, 
        Y => N_9);
    
    \GP_PG_SM_RNO_2[2]\ : OR2B
      port map(A => N_47, B => \GP_PG_SM[2]_net_1\, Y => N_65);
    
    \RX_SER_WORD_3DEL[7]\ : DFN1P0
      port map(D => \RX_SER_WORD_2DEL_i[7]\, CLK => CLK_40M_GL, 
        PRE => P_MASTER_POR_B_c_24, Q => 
        \RX_SER_WORD_3DEL_i_0[7]\);
    
    \RX_SER_WORD_3DEL_RNI019I4[0]\ : NOR2B
      port map(A => un1_RX_SER_WORD_2DEL_1, B => 
        un1_RX_SER_WORD_3DEL_1, Y => N_210_li);
    
    \LOC_STOP_ADDR[2]\ : DFN1E1C0
      port map(D => TFC_STOP_ADDR(2), CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_1, E => \GP_PG_SM_0[10]_net_1\, Q => 
        \LOC_STOP_ADDR[2]_net_1\);
    
    un1_ADDR_POINTER_2_I_28 : XOR2
      port map(A => \TFC_ADDRB[5]\, B => 
        \DWACT_ADD_CI_0_g_array_12_1[0]\, Y => I_28);
    
    \ADDR_POINTER_RNO[5]\ : NOR3
      port map(A => N_89, B => N_374, C => N_373, Y => N_28);
    
    \LOC_STOP_ADDR[1]\ : DFN1E1C0
      port map(D => TFC_STOP_ADDR(1), CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_1, E => \GP_PG_SM_0[10]_net_1\, Q => 
        \LOC_STOP_ADDR[1]_net_1\);
    
    \GP_PG_SM_RNO[8]\ : NOR3C
      port map(A => N_315, B => \GP_PG_SM_ns_i_i_a4_0[2]\, C => 
        N_116, Y => N_80);
    
    \GP_PG_SM_RNIHRVF[3]\ : OR2
      port map(A => \GP_PG_SM[3]_net_1\, B => \GP_PG_SM[2]_net_1\, 
        Y => N_39);
    
    \RX_SER_WORD_1DEL[0]\ : DFN1C0
      port map(D => TFC_RX_SER_WORD(0), CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_30, Q => \RX_SER_WORD_1DEL[0]_net_1\);
    
    \ADDR_POINTER_RNO_0[5]\ : OA1B
      port map(A => N_107, B => \N_ADDR_POINTER_i_o2_0[7]\, C => 
        TFC_STRT_ADDR(5), Y => N_89);
    
    \GP_PG_SM_RNI6RVV[5]\ : NOR2
      port map(A => N_40, B => N_39, Y => N_110);
    
    \RX_SER_WORD_3DEL[0]\ : DFN1C0
      port map(D => \RX_SER_WORD_2DEL[0]_net_1\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_24, Q => 
        \RX_SER_WORD_3DEL[0]_net_1\);
    
    un1_ADDR_POINTER_2_I_31 : XOR2
      port map(A => \TFC_ADDRB[6]\, B => 
        \DWACT_ADD_CI_0_g_array_11[0]\, Y => I_31);
    
    \ADDR_POINTER_RNO[3]\ : NOR3
      port map(A => N_378, B => N_380, C => N_379, Y => N_32);
    
    \ADDR_POINTER[1]\ : DFN1C0
      port map(D => N_36, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_30, Q => \TFC_ADDRB[1]\);
    
    \GP_PG_SM[0]\ : DFN1C0
      port map(D => \GP_PG_SM_ns[10]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_28, Q => \GP_PG_SM[0]_net_1\);
    
    \LOC_STRT_ADDR[5]\ : DFN1E1C0
      port map(D => TFC_STRT_ADDR(5), CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_4, E => \GP_PG_SM_0[10]_net_1\, Q => 
        \LOC_STRT_ADDR[5]_net_1\);
    
    \ADDR_POINTER_RNO_2[7]\ : NOR3A
      port map(A => N_42, B => \GP_PG_SM[10]_net_1\, C => I_34, Y
         => N_84);
    
    \ADDR_POINTER_RNO_1[0]\ : NOR3A
      port map(A => N_39, B => N_214_li, C => 
        \LOC_STRT_ADDR[0]_net_1\, Y => N_106);
    
    \RX_SER_WORD_2DEL_RNIE4KR1[4]\ : OR3
      port map(A => \RX_SER_WORD_2DEL[5]_net_1\, B => 
        \RX_SER_WORD_2DEL[4]_net_1\, C => 
        un1_RX_SER_WORD_2DEL_NE_1, Y => un1_RX_SER_WORD_2DEL_NE_4);
    
    \GP_PG_SM_RNO_0[3]\ : NOR3C
      port map(A => OP_MODE_0, B => \GP_PG_SM[8]_net_1\, C => 
        N_114, Y => \GP_PG_SM_ns_i_i_a4_0_1[7]\);
    
    \GP_PG.un1_ADDR_POINTER_0_I_17\ : OR2A
      port map(A => \LOC_STOP_ADDR[4]_net_1\, B => \TFC_ADDRB[4]\, 
        Y => N_5);
    
    \ADDR_POINTER_RNO_2[0]\ : OA1B
      port map(A => N_107, B => \N_ADDR_POINTER_i_o2_0[7]\, C => 
        TFC_STRT_ADDR(0), Y => N_104);
    
    R_BLKB : DFN1E0P0
      port map(D => N_160_3, CLK => CLK_40M_GL, PRE => 
        P_MASTER_POR_B_c_9, E => N_238, Q => TFC_RAM_BLKB_EN);
    
    \LOC_STRT_ADDR[0]\ : DFN1E1C0
      port map(D => TFC_STRT_ADDR(0), CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_4, E => \GP_PG_SM_0[10]_net_1\, Q => 
        \LOC_STRT_ADDR[0]_net_1\);
    
    \GP_PG_SM_RNO[7]\ : OA1
      port map(A => \GP_PG_SM_ns_0_a2_0[3]\, B => 
        \GP_PG_SM_ns_0_a2_0_1[3]\, C => N_25, Y => 
        \GP_PG_SM_ns[3]\);
    
    \RX_SER_WORD_3DEL_RNO[2]\ : INV
      port map(A => \RX_SER_WORD_2DEL[2]_net_1\, Y => 
        \RX_SER_WORD_2DEL_i[2]\);
    
    \GP_PG_SM_RNO_1[5]\ : NOR3C
      port map(A => N_214_li, B => N_117, C => 
        \GP_PG_SM_ns_0_a2_0[5]\, Y => N_18);
    
    \RX_SER_WORD_1DEL[4]\ : DFN1C0
      port map(D => TFC_RX_SER_WORD(4), CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_31, Q => \RX_SER_WORD_1DEL[4]_net_1\);
    
    \ADDR_POINTER[6]\ : DFN1C0
      port map(D => N_26, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_30, Q => \TFC_ADDRB[6]\);
    
    \GP_PG.un1_ADDR_POINTER_0_I_7\ : NOR2A
      port map(A => \LOC_STOP_ADDR[5]_net_1\, B => \TFC_ADDRB[5]\, 
        Y => \ACT_LT3_E[0]\);
    
    \RX_SER_WORD_1DEL[2]\ : DFN1C0
      port map(D => TFC_RX_SER_WORD(2), CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_31, Q => \RX_SER_WORD_1DEL[2]_net_1\);
    
    \RX_SER_WORD_3DEL[4]\ : DFN1C0
      port map(D => \RX_SER_WORD_2DEL[4]_net_1\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_24, Q => 
        \RX_SER_WORD_3DEL[4]_net_1\);
    
    R_BLKB_RNO : OR3A
      port map(A => OP_MODE_c_0, B => \GP_PG_SM[1]_net_1\, C => 
        N_45, Y => N_160_3);
    
    \ADDR_POINTER_RNO_1[6]\ : NOR3A
      port map(A => N_39, B => N_214_li, C => 
        \LOC_STRT_ADDR[6]_net_1\, Y => N_88);
    
    \RX_SER_WORD_3DEL[2]\ : DFN1P0
      port map(D => \RX_SER_WORD_2DEL_i[2]\, CLK => CLK_40M_GL, 
        PRE => P_MASTER_POR_B_c_24, Q => 
        \RX_SER_WORD_3DEL_i_0[2]\);
    
    \GP_PG.un1_ADDR_POINTER_0_I_13\ : AOI1A
      port map(A => \ACT_LT3_E[3]\, B => \ACT_LT3_E[4]\, C => 
        \ACT_LT3_E[5]\, Y => \DWACT_COMP0_E[0]\);
    
    \GP_PG_SM_RNO[9]\ : NOR3C
      port map(A => \GP_PG_SM_ns_i_i_a4_1[1]\, B => N_315, C => 
        N_116, Y => N_69);
    
    \GP_PG_SM_RNISG4E6[5]\ : NOR3A
      port map(A => N_40, B => N_39, C => N_214_li, Y => N_107);
    
    \GP_PG.un1_ADDR_POINTER_0_I_1\ : XNOR2
      port map(A => \TFC_ADDRB[7]\, B => \LOC_STOP_ADDR[7]_net_1\, 
        Y => \DWACT_BL_EQUAL_0_E[2]\);
    
    \ADDR_POINTER_RNO_0[7]\ : OA1B
      port map(A => N_107, B => \N_ADDR_POINTER_i_o2_0[7]\, C => 
        TFC_STRT_ADDR(7), Y => N_83);
    
    \GP_PG.un1_ADDR_POINTER_0_I_4\ : AND3
      port map(A => \DWACT_BL_EQUAL_0_E[2]\, B => 
        \DWACT_BL_EQUAL_0_E[1]\, C => \DWACT_BL_EQUAL_0_E[0]\, Y
         => \DWACT_COMP0_E[1]\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    un1_ADDR_POINTER_2_I_34 : XOR2
      port map(A => \TFC_ADDRB[7]\, B => 
        \DWACT_ADD_CI_0_g_array_12_2[0]\, Y => I_34);
    
    LOC_DIR_MODE_RNIJUPO : AO1C
      port map(A => N_213_li, B => ALIGN_ACTIVE, C => 
        P_USB_MASTER_EN_c_22_0, Y => N_45);
    
    \GP_PG_SM_RNIDNVF[1]\ : OR2
      port map(A => \GP_PG_SM[1]_net_1\, B => \GP_PG_SM[0]_net_1\, 
        Y => N_61);
    
    \GP_PG.un1_ADDR_POINTER_0_I_24\ : OA1
      port map(A => N_11, B => N_10, C => N_9, Y => 
        \DWACT_COMP0_E[2]\);
    
    un1_ADDR_POINTER_2_I_33 : XOR2
      port map(A => \TFC_ADDRB[4]\, B => 
        \DWACT_ADD_CI_0_g_array_2[0]\, Y => I_33);
    
    \GP_PG_SM[6]\ : DFN1C0
      port map(D => N_22, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_28, Q => \GP_PG_SM[6]_net_1\);
    
    \RX_SER_WORD_2DEL_RNI94QT[6]\ : OR2A
      port map(A => \RX_SER_WORD_2DEL[7]_net_1\, B => 
        \RX_SER_WORD_2DEL[6]_net_1\, Y => 
        un1_RX_SER_WORD_2DEL_NE_1);
    
    \GP_PG_SM_RNO_1[2]\ : AOI1B
      port map(A => \GP_PG_SM[6]_net_1\, B => OP_MODE_0, C => 
        N_65, Y => N_74);
    
    \LOC_STOP_ADDR[4]\ : DFN1E1C0
      port map(D => TFC_STOP_ADDR(4), CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_1, E => \GP_PG_SM_0[10]_net_1\, Q => 
        \LOC_STOP_ADDR[4]_net_1\);
    
    \LOC_STOP_ADDR[5]\ : DFN1E1C0
      port map(D => TFC_STOP_ADDR(5), CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_1, E => \GP_PG_SM_0[10]_net_1\, Q => 
        \LOC_STOP_ADDR[5]_net_1\);
    
    \ADDR_POINTER_RNO_0[0]\ : NOR3A
      port map(A => N_42, B => \GP_PG_SM[10]_net_1\, C => 
        \DWACT_ADD_CI_0_partial_sum[0]\, Y => N_105);
    
    un1_ADDR_POINTER_2_I_36 : NOR2B
      port map(A => \DWACT_ADD_CI_0_TMP[0]\, B => \TFC_ADDRB[1]\, 
        Y => \DWACT_ADD_CI_0_g_array_1[0]\);
    
    \GP_PG.un1_ADDR_POINTER_0_I_12\ : AND2A
      port map(A => \LOC_STOP_ADDR[7]_net_1\, B => \TFC_ADDRB[7]\, 
        Y => \ACT_LT3_E[5]\);
    
    un1_ADDR_POINTER_2_I_29 : XOR2
      port map(A => \TFC_ADDRB[2]\, B => 
        \DWACT_ADD_CI_0_g_array_1[0]\, Y => I_29);
    
    \GP_PG_SM[5]\ : DFN1C0
      port map(D => \GP_PG_SM_ns[5]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_28, Q => \GP_PG_SM[5]_net_1\);
    
    un1_ADDR_POINTER_2_I_35 : NOR2B
      port map(A => \DWACT_ADD_CI_0_g_array_1[0]\, B => 
        \DWACT_ADD_CI_0_pog_array_1[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_2[0]\);
    
    \GP_PG_SM_RNIT7081[9]\ : NOR3A
      port map(A => N_315, B => \GP_PG_SM[1]_net_1\, C => 
        \GP_PG_SM[9]_net_1\, Y => \GP_PG_SM_ns_0_a4_1[0]\);
    
    \ADDR_POINTER_RNO[4]\ : NOR3
      port map(A => N_375, B => N_377, C => N_376, Y => N_30);
    
    \ADDR_POINTER[0]\ : DFN1C0
      port map(D => N_38, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_30, Q => \TFC_ADDRB[0]\);
    
    \RX_SER_WORD_3DEL_RNIISGD[4]\ : OR3
      port map(A => \RX_SER_WORD_3DEL[5]_net_1\, B => 
        \RX_SER_WORD_3DEL[4]_net_1\, C => 
        un1_RX_SER_WORD_3DEL_NE_1, Y => un1_RX_SER_WORD_3DEL_NE_4);
    
    \GP_PG_SM_RNICMV71[5]\ : NOR2A
      port map(A => N_117, B => N_40, Y => N_25);
    
    \GP_PG_SM_RNO_0[9]\ : NOR3A
      port map(A => OP_MODE_c_0, B => \GP_PG_SM[9]_net_1\, C => 
        N_45, Y => \GP_PG_SM_ns_i_i_a4_1[1]\);
    
    \GP_PG_SM_RNO[2]\ : AOI1
      port map(A => N_64, B => \GP_PG_SM[0]_net_1\, C => N_74, Y
         => \GP_PG_SM_RNO[2]_net_1\);
    
    \ADDR_POINTER_RNO[0]\ : NOR3
      port map(A => N_105, B => N_106, C => N_104, Y => N_38);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \GP_PG_SM_RNIU8V56[10]\ : OA1A
      port map(A => N_39, B => N_214_li, C => 
        \GP_PG_SM[10]_net_1\, Y => \N_ADDR_POINTER_i_o2_0[7]\);
    
    \ADDR_POINTER_RNO_0[2]\ : NOR3A
      port map(A => N_42, B => \GP_PG_SM[10]_net_1\, C => I_29, Y
         => N_382);
    
    \GP_PG_SM[7]\ : DFN1C0
      port map(D => \GP_PG_SM_ns[3]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_28, Q => \GP_PG_SM[7]_net_1\);
    
    \RX_SER_WORD_2DEL_RNICO7N3[0]\ : OR3
      port map(A => un1_RX_SER_WORD_2DEL_NE_3, B => 
        un1_RX_SER_WORD_2DEL_NE_2, C => un1_RX_SER_WORD_2DEL_NE_4, 
        Y => un1_RX_SER_WORD_2DEL_1);
    
    \GP_PG_SM_RNO_2[5]\ : NOR2A
      port map(A => \GP_PG_SM[5]_net_1\, B => \GP_PG_SM[4]_net_1\, 
        Y => \GP_PG_SM_ns_0_a2_0[5]\);
    
    \GP_PG_SM[1]\ : DFN1C0
      port map(D => \GP_PG_SM_RNO[1]_net_1\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_28, Q => \GP_PG_SM[1]_net_1\);
    
    \GP_PG.un1_ADDR_POINTER_0_I_19\ : OA1A
      port map(A => \TFC_ADDRB[3]\, B => \LOC_STOP_ADDR[3]_net_1\, 
        C => N_3, Y => N_7);
    
    un1_ADDR_POINTER_2_I_1 : AND2
      port map(A => \TFC_ADDRB[0]\, B => 
        \GP_PG_SM_RNITIQ71[10]_net_1\, Y => 
        \DWACT_ADD_CI_0_TMP[0]\);
    
    \GP_PG_SM_RNO_1[3]\ : NOR3B
      port map(A => \GP_PG_SM_ns_i_i_a4_0[7]\, B => N_47, C => 
        N_61, Y => N_76);
    
    \GP_PG_SM_RNO_2[3]\ : NOR2A
      port map(A => \GP_PG_SM[3]_net_1\, B => \GP_PG_SM[2]_net_1\, 
        Y => \GP_PG_SM_ns_i_i_a4_0[7]\);
    
    \GP_PG_SM_RNO[4]\ : AO1
      port map(A => \GP_PG_SM_ns_0_a4_0[6]\, B => N_117, C => 
        N_79, Y => \GP_PG_SM_ns[6]\);
    
    \GP_PG_SM_RNISG4E6_0[5]\ : OR2
      port map(A => N_110, B => N_214_li, Y => N_42);
    
    LOC_DIR_MODE : DFN1E1C0
      port map(D => DCB_SALT_SEL_c, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_15, E => \GP_PG_SM[10]_net_1\, Q => 
        N_213_li);
    
    \ADDR_POINTER_RNO_2[3]\ : NOR3A
      port map(A => N_42, B => \GP_PG_SM[10]_net_1\, C => I_27, Y
         => N_379);
    
    un1_ADDR_POINTER_2_I_27 : XOR2
      port map(A => \TFC_ADDRB[3]\, B => 
        \DWACT_ADD_CI_0_g_array_12[0]\, Y => I_27);
    
    \ADDR_POINTER_RNO_1[7]\ : NOR3A
      port map(A => N_39, B => N_214_li, C => 
        \LOC_STRT_ADDR[7]_net_1\, Y => N_85);
    
    \RX_SER_WORD_3DEL_RNO[1]\ : INV
      port map(A => \RX_SER_WORD_2DEL[1]_net_1\, Y => 
        \RX_SER_WORD_2DEL_i[1]\);
    
    \GP_PG_SM[10]\ : DFN1P0
      port map(D => \GP_PG_SM_ns[0]\, CLK => CLK_40M_GL, PRE => 
        P_MASTER_POR_B_c_27_1, Q => \GP_PG_SM[10]_net_1\);
    
    un1_ADDR_POINTER_2_I_49 : AND2
      port map(A => \TFC_ADDRB[4]\, B => \TFC_ADDRB[5]\, Y => 
        \DWACT_ADD_CI_0_pog_array_1_1[0]\);
    
    \ADDR_POINTER[4]\ : DFN1C0
      port map(D => N_30, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_30, Q => \TFC_ADDRB[4]\);
    
    \GP_PG.un1_ADDR_POINTER_0_I_20\ : AO1C
      port map(A => \TFC_ADDRB[2]\, B => \LOC_STOP_ADDR[2]_net_1\, 
        C => N_2, Y => N_8);
    
    \GP_PG_SM_ns_i_i_o2[7]\ : OR2
      port map(A => N_214_li, B => OP_MODE_c_0, Y => N_47);
    
    \GP_PG.un1_ADDR_POINTER_0_I_15\ : OR2A
      port map(A => \TFC_ADDRB[2]\, B => \LOC_STOP_ADDR[2]_net_1\, 
        Y => N_3);
    
    \GP_PG_SM[4]\ : DFN1C0
      port map(D => \GP_PG_SM_ns[6]\, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_28, Q => \GP_PG_SM[4]_net_1\);
    
    \GP_PG_SM_RNO_0[2]\ : OR3C
      port map(A => OP_MODE_c_0, B => \GP_PG_SM[2]_net_1\, C => 
        N_214_li, Y => N_64);
    
    \RX_SER_WORD_2DEL[6]\ : DFN1C0
      port map(D => \RX_SER_WORD_1DEL[6]_net_1\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c, Q => 
        \RX_SER_WORD_2DEL[6]_net_1\);
    
    \GP_PG.un1_ADDR_POINTER_0_I_11\ : OR2A
      port map(A => \LOC_STOP_ADDR[7]_net_1\, B => \TFC_ADDRB[7]\, 
        Y => \ACT_LT3_E[4]\);
    
    \ADDR_POINTER_RNO_1[2]\ : NOR3A
      port map(A => N_39, B => N_214_li, C => 
        \LOC_STRT_ADDR[2]_net_1\, Y => N_383);
    
    \GP_PG_SM_RNO_0[4]\ : NOR2A
      port map(A => \GP_PG_SM[6]_net_1\, B => OP_MODE_0, Y => 
        \GP_PG_SM_ns_0_a4_0[6]\);
    
    \GP_PG_SM_RNI0RDP3[0]\ : AO1A
      port map(A => OP_MODE_c_0, B => \GP_PG_SM[0]_net_1\, C => 
        N_71, Y => \GP_PG_SM_ns[0]\);
    
    \GP_PG_SM_RNIJIVF1[1]\ : NOR2A
      port map(A => N_110, B => N_61, Y => N_116);
    
    \ADDR_POINTER_RNO[2]\ : NOR3
      port map(A => N_382, B => N_383, C => N_381, Y => N_34);
    
    \LOC_STOP_ADDR[7]\ : DFN1E1C0
      port map(D => TFC_STOP_ADDR(7), CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_1, E => \GP_PG_SM_0[10]_net_1\, Q => 
        \LOC_STOP_ADDR[7]_net_1\);
    
    \ADDR_POINTER_RNO[1]\ : NOR3
      port map(A => N_102, B => N_103, C => N_101, Y => N_36);
    
    \RX_SER_WORD_3DEL_RNI38O6[2]\ : OR2
      port map(A => \RX_SER_WORD_3DEL_i_0[2]\, B => 
        \RX_SER_WORD_3DEL_i_0[3]\, Y => un1_RX_SER_WORD_3DEL_NE_3);
    
    \GP_PG_SM_RNITIQ71[10]\ : OR2A
      port map(A => N_110, B => \GP_PG_SM[10]_net_1\, Y => 
        \GP_PG_SM_RNITIQ71[10]_net_1\);
    
    \GP_PG_SM_0[10]\ : DFN1P0
      port map(D => \GP_PG_SM_ns[0]\, CLK => CLK_40M_GL, PRE => 
        P_MASTER_POR_B_c_27_1, Q => \GP_PG_SM_0[10]_net_1\);
    
    \RX_SER_WORD_2DEL_RNI1SPT[2]\ : OR2B
      port map(A => \RX_SER_WORD_2DEL[2]_net_1\, B => 
        \RX_SER_WORD_2DEL[3]_net_1\, Y => 
        un1_RX_SER_WORD_2DEL_NE_3);
    
    \LOC_STRT_ADDR[2]\ : DFN1E1C0
      port map(D => TFC_STRT_ADDR(2), CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_4, E => \GP_PG_SM_0[10]_net_1\, Q => 
        \LOC_STRT_ADDR[2]_net_1\);
    
    \RX_SER_WORD_2DEL[5]\ : DFN1C0
      port map(D => \RX_SER_WORD_1DEL[5]_net_1\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c, Q => 
        \RX_SER_WORD_2DEL[5]_net_1\);
    
    \ADDR_POINTER_RNO_0[1]\ : NOR3A
      port map(A => N_42, B => \GP_PG_SM[10]_net_1\, C => I_30, Y
         => N_102);
    
    \RX_SER_WORD_2DEL[3]\ : DFN1C0
      port map(D => \RX_SER_WORD_1DEL[3]_net_1\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c, Q => 
        \RX_SER_WORD_2DEL[3]_net_1\);
    
    \GP_PG_SM_RNO[6]\ : NOR3C
      port map(A => N_210_li, B => \GP_PG_SM[7]_net_1\, C => 
        N_116, Y => N_22);
    
    \GP_PG_SM_RNIBU3D3[0]\ : NOR3C
      port map(A => N_50, B => \GP_PG_SM_ns_0_a4_1[0]\, C => 
        N_110, Y => N_71);
    
    \ADDR_POINTER_RNO_1[5]\ : NOR3A
      port map(A => N_39, B => N_214_li, C => 
        \LOC_STRT_ADDR[5]_net_1\, Y => N_374);
    
    \GP_PG_SM_RNI8R351[0]\ : AO1C
      port map(A => \GP_PG_SM[0]_net_1\, B => N_45, C => 
        OP_MODE_c_0, Y => N_50);
    
    \LOC_STRT_ADDR[3]\ : DFN1E1C0
      port map(D => TFC_STRT_ADDR(3), CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_4, E => \GP_PG_SM_0[10]_net_1\, Q => 
        \LOC_STRT_ADDR[3]_net_1\);
    
    \RX_SER_WORD_3DEL_RNIK81R[0]\ : OR3
      port map(A => un1_RX_SER_WORD_3DEL_NE_3, B => 
        un1_RX_SER_WORD_3DEL_NE_2, C => un1_RX_SER_WORD_3DEL_NE_4, 
        Y => un1_RX_SER_WORD_3DEL_1);
    
    \LOC_STRT_ADDR[1]\ : DFN1E1C0
      port map(D => TFC_STRT_ADDR(1), CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_4, E => \GP_PG_SM_0[10]_net_1\, Q => 
        \LOC_STRT_ADDR[1]_net_1\);
    
    \LOC_STRT_ADDR[7]\ : DFN1E1C0
      port map(D => TFC_STRT_ADDR(7), CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_5, E => \GP_PG_SM[10]_net_1\, Q => 
        \LOC_STRT_ADDR[7]_net_1\);
    
    \GP_PG_SM[8]\ : DFN1C0
      port map(D => N_80, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_28, Q => \GP_PG_SM[8]_net_1\);
    
    \GP_PG.un1_ADDR_POINTER_0_I_9\ : AND2A
      port map(A => \LOC_STOP_ADDR[6]_net_1\, B => \TFC_ADDRB[6]\, 
        Y => \ACT_LT3_E[2]\);
    
    \GP_PG.un1_ADDR_POINTER_0_I_3\ : XNOR2
      port map(A => \TFC_ADDRB[5]\, B => \LOC_STOP_ADDR[5]_net_1\, 
        Y => \DWACT_BL_EQUAL_0_E[0]\);
    
    \ADDR_POINTER_RNO_1[1]\ : NOR3A
      port map(A => N_39, B => N_214_li, C => 
        \LOC_STRT_ADDR[1]_net_1\, Y => N_103);
    
    \ADDR_POINTER_RNO_2[2]\ : OA1B
      port map(A => N_107, B => \N_ADDR_POINTER_i_o2_0[7]\, C => 
        TFC_STRT_ADDR(2), Y => N_381);
    
    \GP_PG_SM[3]\ : DFN1C0
      port map(D => \GP_PG_SM_RNO[3]_net_1\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_28, Q => \GP_PG_SM[3]_net_1\);
    
    \RX_SER_WORD_3DEL_RNO[7]\ : INV
      port map(A => \RX_SER_WORD_2DEL[7]_net_1\, Y => 
        \RX_SER_WORD_2DEL_i[7]\);
    
    \ADDR_POINTER[3]\ : DFN1C0
      port map(D => N_32, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_30, Q => \TFC_ADDRB[3]\);
    
    \RX_SER_WORD_2DEL[1]\ : DFN1C0
      port map(D => \RX_SER_WORD_1DEL[1]_net_1\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c, Q => 
        \RX_SER_WORD_2DEL[1]_net_1\);
    
    \GP_PG_SM_RNO_0[5]\ : NOR3B
      port map(A => \GP_PG_SM[8]_net_1\, B => N_114, C => 
        OP_MODE_0, Y => \GP_PG_SM_ns_0_a2_0_1[5]\);
    
    \GP_PG.un1_ADDR_POINTER_0_I_23\ : OA1A
      port map(A => N_6, B => N_8, C => N_7, Y => N_11);
    
    \RX_SER_WORD_3DEL_RNIBGO6[6]\ : OR2
      port map(A => \RX_SER_WORD_3DEL[6]_net_1\, B => 
        \RX_SER_WORD_3DEL_i_0[7]\, Y => un1_RX_SER_WORD_3DEL_NE_1);
    
    \GP_PG.un1_ADDR_POINTER_0_I_2\ : XNOR2
      port map(A => \TFC_ADDRB[6]\, B => \LOC_STOP_ADDR[6]_net_1\, 
        Y => \DWACT_BL_EQUAL_0_E[1]\);
    
    \GP_PG_SM_RNI770O[8]\ : NOR2A
      port map(A => N_114, B => \GP_PG_SM[8]_net_1\, Y => N_315);
    
    \GP_PG.un1_ADDR_POINTER_0_I_14\ : OR2A
      port map(A => \LOC_STOP_ADDR[1]_net_1\, B => \TFC_ADDRB[1]\, 
        Y => N_2);
    
    \ADDR_POINTER_RNO_2[6]\ : NOR3A
      port map(A => N_42, B => \GP_PG_SM[10]_net_1\, C => I_31, Y
         => N_87);
    
    \RX_SER_WORD_3DEL_RNO[3]\ : INV
      port map(A => \RX_SER_WORD_2DEL[3]_net_1\, Y => 
        \RX_SER_WORD_2DEL_i[3]\);
    
    \ADDR_POINTER_RNO[7]\ : NOR3
      port map(A => N_83, B => N_85, C => N_84, Y => N_24);
    
    \GP_PG.un1_ADDR_POINTER_0_I_8\ : OR2A
      port map(A => \LOC_STOP_ADDR[6]_net_1\, B => \TFC_ADDRB[6]\, 
        Y => \ACT_LT3_E[1]\);
    
    \ADDR_POINTER[7]\ : DFN1C0
      port map(D => N_24, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_30, Q => \TFC_ADDRB[7]\);
    
    \LOC_STOP_ADDR[3]\ : DFN1E1C0
      port map(D => TFC_STOP_ADDR(3), CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_1, E => \GP_PG_SM_0[10]_net_1\, Q => 
        \LOC_STOP_ADDR[3]_net_1\);
    
    \RX_SER_WORD_1DEL[6]\ : DFN1C0
      port map(D => TFC_RX_SER_WORD(6), CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_31, Q => \RX_SER_WORD_1DEL[6]_net_1\);
    
    \RX_SER_WORD_2DEL[7]\ : DFN1C0
      port map(D => \RX_SER_WORD_1DEL[7]_net_1\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c, Q => 
        \RX_SER_WORD_2DEL[7]_net_1\);
    
    \GP_PG_SM_RNO_1[7]\ : NOR3B
      port map(A => \GP_PG_SM[9]_net_1\, B => N_315, C => 
        N_213_li, Y => \GP_PG_SM_ns_0_a2_0_1[3]\);
    
    un1_ADDR_POINTER_2_I_24 : XOR2
      port map(A => \TFC_ADDRB[0]\, B => 
        \GP_PG_SM_RNITIQ71[10]_net_1\, Y => 
        \DWACT_ADD_CI_0_partial_sum[0]\);
    
    \RX_SER_WORD_3DEL[6]\ : DFN1C0
      port map(D => \RX_SER_WORD_2DEL[6]_net_1\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_24, Q => 
        \RX_SER_WORD_3DEL[6]_net_1\);
    
    \GP_PG_SM_RNO[0]\ : AO1
      port map(A => \GP_PG_SM[0]_net_1\, B => OP_MODE_c_0, C => 
        \GP_PG_SM[1]_net_1\, Y => \GP_PG_SM_ns[10]\);
    
    \GP_PG_SM[9]\ : DFN1C0
      port map(D => N_69, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_28, Q => \GP_PG_SM[9]_net_1\);
    
    \ADDR_POINTER_RNO_2[5]\ : NOR3A
      port map(A => N_42, B => \GP_PG_SM[10]_net_1\, C => I_28, Y
         => N_373);
    
    un1_ADDR_POINTER_2_I_41 : NOR2B
      port map(A => \DWACT_ADD_CI_0_g_array_2[0]\, B => 
        \DWACT_ADD_CI_0_pog_array_1_1[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_11[0]\);
    
    \ADDR_POINTER_RNO_1[4]\ : NOR3A
      port map(A => N_39, B => N_214_li, C => 
        \LOC_STRT_ADDR[4]_net_1\, Y => N_377);
    
    \GP_PG.un1_ADDR_POINTER_0_I_22\ : AO1C
      port map(A => \TFC_ADDRB[3]\, B => \LOC_STOP_ADDR[3]_net_1\, 
        C => N_5, Y => N_10);
    
    \RX_SER_WORD_2DEL[0]\ : DFN1C0
      port map(D => \RX_SER_WORD_1DEL[0]_net_1\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c, Q => 
        \RX_SER_WORD_2DEL[0]_net_1\);
    
    \LOC_STOP_ADDR[0]\ : DFN1E1C0
      port map(D => TFC_STOP_ADDR(0), CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_1, E => \GP_PG_SM_0[10]_net_1\, Q => 
        \LOC_STOP_ADDR[0]_net_1\);
    
    \RX_SER_WORD_1DEL[5]\ : DFN1C0
      port map(D => TFC_RX_SER_WORD(5), CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_31, Q => \RX_SER_WORD_1DEL[5]_net_1\);
    
    \GP_PG.un1_ADDR_POINTER_0_I_18\ : AO1C
      port map(A => \LOC_STOP_ADDR[1]_net_1\, B => \TFC_ADDRB[1]\, 
        C => N_4, Y => N_6);
    
    \RX_SER_WORD_1DEL[3]\ : DFN1C0
      port map(D => TFC_RX_SER_WORD(3), CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_31, Q => \RX_SER_WORD_1DEL[3]_net_1\);
    
    \GP_PG_SM[2]\ : DFN1C0
      port map(D => \GP_PG_SM_RNO[2]_net_1\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_28, Q => \GP_PG_SM[2]_net_1\);
    
    un1_ADDR_POINTER_2_I_30 : XOR2
      port map(A => \TFC_ADDRB[1]\, B => \DWACT_ADD_CI_0_TMP[0]\, 
        Y => I_30);
    
    \RX_SER_WORD_3DEL[5]\ : DFN1C0
      port map(D => \RX_SER_WORD_2DEL[5]_net_1\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_24, Q => 
        \RX_SER_WORD_3DEL[5]_net_1\);
    
    \RX_SER_WORD_2DEL_RNITNPT[0]\ : OR2A
      port map(A => \RX_SER_WORD_2DEL[1]_net_1\, B => 
        \RX_SER_WORD_2DEL[0]_net_1\, Y => 
        un1_RX_SER_WORD_2DEL_NE_2);
    
    \GP_PG_SM_RNO[5]\ : AO1
      port map(A => \GP_PG_SM_ns_0_a2_0_1[5]\, B => N_25, C => 
        N_18, Y => \GP_PG_SM_ns[5]\);
    
    \RX_SER_WORD_3DEL[3]\ : DFN1P0
      port map(D => \RX_SER_WORD_2DEL_i[3]\, CLK => CLK_40M_GL, 
        PRE => P_MASTER_POR_B_c_24, Q => 
        \RX_SER_WORD_3DEL_i_0[3]\);
    
    \GP_PG_SM_RNINMVN[0]\ : NOR2
      port map(A => \GP_PG_SM[0]_net_1\, B => N_39, Y => N_117);
    
    \GP_PG_SM_RNO[3]\ : AO1
      port map(A => \GP_PG_SM_ns_i_i_a4_0_1[7]\, B => N_116, C
         => N_76, Y => \GP_PG_SM_RNO[3]_net_1\);
    
    \GP_PG_SM_RNILVVF[5]\ : OR2
      port map(A => \GP_PG_SM[5]_net_1\, B => \GP_PG_SM[4]_net_1\, 
        Y => N_40);
    
    \GP_PG_SM_RNO_0[7]\ : NOR2A
      port map(A => \GP_PG_SM[7]_net_1\, B => N_210_li, Y => 
        \GP_PG_SM_ns_0_a2_0[3]\);
    
    \LOC_STRT_ADDR[4]\ : DFN1E1C0
      port map(D => TFC_STRT_ADDR(4), CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_4, E => \GP_PG_SM_0[10]_net_1\, Q => 
        \LOC_STRT_ADDR[4]_net_1\);
    
    \GP_PG_SM_RNO[1]\ : NOR3
      port map(A => N_73, B => N_61, C => N_42, Y => 
        \GP_PG_SM_RNO[1]_net_1\);
    
    \ADDR_POINTER[5]\ : DFN1C0
      port map(D => N_28, CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_30, Q => \TFC_ADDRB[5]\);
    
    R_RWB : DFN1E1P0
      port map(D => N_213_li, CLK => CLK_40M_GL, PRE => 
        P_MASTER_POR_B_c_16_0, E => \GP_PG_SM[10]_net_1\, Q => 
        TFC_RWB);
    
    R_BLKB_RNO_0 : NOR2
      port map(A => \GP_PG_SM[1]_net_1\, B => 
        \GP_PG_SM[10]_net_1\, Y => N_238);
    
    \ADDR_POINTER_RNO_1[3]\ : NOR3A
      port map(A => N_39, B => N_214_li, C => 
        \LOC_STRT_ADDR[3]_net_1\, Y => N_380);
    
    \RX_SER_WORD_3DEL_RNIV3O6[0]\ : OR2
      port map(A => \RX_SER_WORD_3DEL[0]_net_1\, B => 
        \RX_SER_WORD_3DEL_i_0[1]\, Y => un1_RX_SER_WORD_3DEL_NE_2);
    
    \ADDR_POINTER_RNO_2[4]\ : NOR3A
      port map(A => N_42, B => \GP_PG_SM[10]_net_1\, C => I_33, Y
         => N_376);
    
    \ADDR_POINTER_RNO[6]\ : NOR3
      port map(A => N_86, B => N_88, C => N_87, Y => N_26);
    
    \RX_SER_WORD_2DEL[4]\ : DFN1C0
      port map(D => \RX_SER_WORD_1DEL[4]_net_1\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c, Q => 
        \RX_SER_WORD_2DEL[4]_net_1\);
    
    \LOC_STRT_ADDR[6]\ : DFN1E1C0
      port map(D => TFC_STRT_ADDR(6), CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_5, E => \GP_PG_SM_0[10]_net_1\, Q => 
        \LOC_STRT_ADDR[6]_net_1\);
    
    un1_ADDR_POINTER_2_I_44 : NOR2B
      port map(A => \DWACT_ADD_CI_0_g_array_11[0]\, B => 
        \TFC_ADDRB[6]\, Y => \DWACT_ADD_CI_0_g_array_12_2[0]\);
    
    \RX_SER_WORD_2DEL[2]\ : DFN1C0
      port map(D => \RX_SER_WORD_1DEL[2]_net_1\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c, Q => 
        \RX_SER_WORD_2DEL[2]_net_1\);
    
    \GP_PG_SM_RNO_0[1]\ : NOR2B
      port map(A => N_39, B => OP_MODE_c_0, Y => N_73);
    
    \LOC_STOP_ADDR[6]\ : DFN1E1C0
      port map(D => TFC_STOP_ADDR(6), CLK => CLK_40M_GL, CLR => 
        P_MASTER_POR_B_c_1, E => \GP_PG_SM_0[10]_net_1\, Q => 
        \LOC_STOP_ADDR[6]_net_1\);
    
    \GP_PG.un1_ADDR_POINTER_0_I_10\ : AOI1A
      port map(A => \ACT_LT3_E[0]\, B => \ACT_LT3_E[1]\, C => 
        \ACT_LT3_E[2]\, Y => \ACT_LT3_E[3]\);
    
    \RX_SER_WORD_1DEL[1]\ : DFN1C0
      port map(D => TFC_RX_SER_WORD(1), CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_30, Q => \RX_SER_WORD_1DEL[1]_net_1\);
    
    un1_ADDR_POINTER_2_I_43 : NOR2B
      port map(A => \DWACT_ADD_CI_0_g_array_2[0]\, B => 
        \TFC_ADDRB[4]\, Y => \DWACT_ADD_CI_0_g_array_12_1[0]\);
    
    \GP_PG.un1_ADDR_POINTER_0_I_16\ : NOR2A
      port map(A => \LOC_STOP_ADDR[0]_net_1\, B => \TFC_ADDRB[0]\, 
        Y => N_4);
    
    \RX_SER_WORD_3DEL[1]\ : DFN1P0
      port map(D => \RX_SER_WORD_2DEL_i[1]\, CLK => CLK_40M_GL, 
        PRE => P_MASTER_POR_B_c_24, Q => 
        \RX_SER_WORD_3DEL_i_0[1]\);
    
    \ADDR_POINTER_RNO_0[3]\ : OA1B
      port map(A => N_107, B => \N_ADDR_POINTER_i_o2_0[7]\, C => 
        TFC_STRT_ADDR(3), Y => N_378);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SLAVE_DES320S_1_17_6 is

    port( ELK_RX_SER_WORD_8      : out   std_logic_vector(7 downto 0);
          BIT_OS_SEL_5           : in    std_logic_vector(1 downto 0);
          BIT_OS_SEL_6_0         : in    std_logic;
          BIT_OS_SEL_3           : in    std_logic_vector(2 downto 1);
          BIT_OS_SEL_4_0         : in    std_logic;
          CLK_40M_GL             : in    std_logic;
          CCC_160M_FXD           : in    std_logic;
          ELK_IN_R               : in    std_logic;
          ELK_IN_F               : in    std_logic;
          MASTER_DCB_POR_B_i_0_i : in    std_logic;
          CCC_160M_ADJ           : in    std_logic
        );

end SLAVE_DES320S_1_17_6;

architecture DEF_ARCH of SLAVE_DES320S_1_17_6 is 

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal N_17, \ARB_BYTE[0]_net_1\, \ARB_BYTE[4]_net_1\, N_18, 
        \ARB_BYTE[1]_net_1\, \ARB_BYTE[5]_net_1\, N_19, 
        \ARB_BYTE[2]_net_1\, \ARB_BYTE[6]_net_1\, N_20, 
        \ARB_BYTE[3]_net_1\, \ARB_BYTE[7]_net_1\, N_21, 
        \ARB_BYTE[8]_net_1\, N_22, \ARB_BYTE[9]_net_1\, N_23, 
        \ARB_BYTE[10]_net_1\, N_24, \ARB_BYTE[11]_net_1\, N_31, 
        \ARB_BYTE[12]_net_1\, N_32, \ARB_BYTE[13]_net_1\, N_33, 
        N_34, N_35, N_36, N_37, N_38, N_39, N_40, N_56, 
        \ARB_BYTE[14]_net_1\, N_64, \N_RECD_SER_WORD[0]\, 
        \N_RECD_SER_WORD[1]\, \N_RECD_SER_WORD[2]\, 
        \N_RECD_SER_WORD[3]\, \N_RECD_SER_WORD[4]\, 
        \N_RECD_SER_WORD[5]\, \N_RECD_SER_WORD[6]\, 
        \N_RECD_SER_WORD[7]\, \ADJ_SER_IN_F_0DEL\, 
        \ADJ_SER_IN_R_0DEL\, \ADJ_SER_IN_F_1DEL\, 
        \ADJ_SER_IN_R_1DEL\, \Q[0]_net_1\, \ADJ_Q[0]_net_1\, 
        \Q[1]_net_1\, \ADJ_Q[1]_net_1\, \Q[2]_net_1\, 
        \ADJ_Q[2]_net_1\, \Q[3]_net_1\, \ADJ_Q[3]_net_1\, 
        \Q[4]_net_1\, \ADJ_Q[4]_net_1\, \Q[5]_net_1\, 
        \ADJ_Q[5]_net_1\, \Q[6]_net_1\, \ADJ_Q[6]_net_1\, 
        \Q[7]_net_1\, \ADJ_Q[7]_net_1\, \Q[8]_net_1\, 
        \ADJ_Q[8]_net_1\, \Q[9]_net_1\, \ADJ_Q[9]_net_1\, 
        \Q[10]_net_1\, \ADJ_Q[10]_net_1\, \Q[11]_net_1\, 
        \ADJ_Q[11]_net_1\, \Q[12]_net_1\, \ADJ_Q[12]_net_1\, 
        \Q[13]_net_1\, \ADJ_Q[13]_net_1\, \Q[14]_net_1\, 
        \ADJ_Q[14]_net_1\, \ARB_WRD_40M_FIXED[0]_net_1\, 
        \ARB_WRD_40M_FIXED[1]_net_1\, 
        \ARB_WRD_40M_FIXED[2]_net_1\, 
        \ARB_WRD_40M_FIXED[3]_net_1\, 
        \ARB_WRD_40M_FIXED[4]_net_1\, 
        \ARB_WRD_40M_FIXED[5]_net_1\, 
        \ARB_WRD_40M_FIXED[6]_net_1\, 
        \ARB_WRD_40M_FIXED[7]_net_1\, 
        \ARB_WRD_40M_FIXED[8]_net_1\, 
        \ARB_WRD_40M_FIXED[9]_net_1\, 
        \ARB_WRD_40M_FIXED[10]_net_1\, 
        \ARB_WRD_40M_FIXED[11]_net_1\, 
        \ARB_WRD_40M_FIXED[12]_net_1\, 
        \ARB_WRD_40M_FIXED[13]_net_1\, 
        \ARB_WRD_40M_FIXED[14]_net_1\, \GND\, \VCC\ : std_logic;

begin 


    \RECD_SER_WORD_RNO[5]\ : MX2
      port map(A => N_38, B => N_39, S => BIT_OS_SEL_5(0), Y => 
        \N_RECD_SER_WORD[5]\);
    
    \ARB_WRD_40M_FIXED[9]\ : DFN1C0
      port map(D => \Q[9]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[9]_net_1\);
    
    \ADJ_Q[4]\ : DFN1C0
      port map(D => \ADJ_Q[2]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[4]_net_1\);
    
    \ARB_BYTE_RNIJLQT[10]\ : MX2
      port map(A => N_21, B => N_23, S => BIT_OS_SEL_3(1), Y => 
        N_37);
    
    \ARB_BYTE[6]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[6]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[6]_net_1\);
    
    ADJ_SER_IN_F_1DEL : DFN1C0
      port map(D => \ADJ_SER_IN_F_0DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_F_1DEL\);
    
    \ARB_BYTE[0]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[0]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[0]_net_1\);
    
    \ARB_BYTE_RNITGAC[12]\ : MX2
      port map(A => \ARB_BYTE[8]_net_1\, B => 
        \ARB_BYTE[12]_net_1\, S => BIT_OS_SEL_4_0, Y => N_31);
    
    \Q[11]\ : DFN1C0
      port map(D => \ADJ_Q[11]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[11]_net_1\);
    
    \ADJ_Q[8]\ : DFN1C0
      port map(D => \ADJ_Q[6]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[8]_net_1\);
    
    \ARB_BYTE_RNI7Q3H[1]\ : MX2
      port map(A => \ARB_BYTE[1]_net_1\, B => \ARB_BYTE[5]_net_1\, 
        S => BIT_OS_SEL_3(2), Y => N_18);
    
    \ADJ_Q[6]\ : DFN1C0
      port map(D => \ADJ_Q[4]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[6]_net_1\);
    
    \ADJ_Q[12]\ : DFN1C0
      port map(D => \ADJ_Q[10]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[12]_net_1\);
    
    \RECD_SER_WORD_RNO_1[0]\ : MX2
      port map(A => \ARB_BYTE[0]_net_1\, B => \ARB_BYTE[4]_net_1\, 
        S => BIT_OS_SEL_3(2), Y => N_17);
    
    \Q[1]\ : DFN1C0
      port map(D => \ADJ_Q[1]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[1]_net_1\);
    
    \ARB_BYTE[4]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[4]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[4]_net_1\);
    
    \ADJ_Q[2]\ : DFN1C0
      port map(D => \ADJ_Q[0]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[2]_net_1\);
    
    \RECD_SER_WORD_RNO_1[7]\ : MX2
      port map(A => \ARB_BYTE[10]_net_1\, B => 
        \ARB_BYTE[14]_net_1\, S => BIT_OS_SEL_6_0, Y => N_56);
    
    \RECD_SER_WORD[4]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[4]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_8(4));
    
    \Q[5]\ : DFN1C0
      port map(D => \ADJ_Q[5]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[5]_net_1\);
    
    \ARB_BYTE_RNI7A1P[13]\ : MX2
      port map(A => N_24, B => N_32, S => BIT_OS_SEL_3(1), Y => 
        N_40);
    
    \ADJ_Q[11]\ : DFN1C0
      port map(D => \ADJ_Q[9]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[11]_net_1\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \ADJ_Q[3]\ : DFN1C0
      port map(D => \ADJ_Q[1]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[3]_net_1\);
    
    \Q[10]\ : DFN1C0
      port map(D => \ADJ_Q[10]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[10]_net_1\);
    
    \ARB_WRD_40M_FIXED[6]\ : DFN1C0
      port map(D => \Q[6]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[6]_net_1\);
    
    \ARB_WRD_40M_FIXED[1]\ : DFN1C0
      port map(D => \Q[1]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[1]_net_1\);
    
    \RECD_SER_WORD[3]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[3]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_8(3));
    
    \RECD_SER_WORD[0]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[0]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_8(0));
    
    \RECD_SER_WORD_RNO[3]\ : MX2
      port map(A => N_36, B => N_37, S => BIT_OS_SEL_5(0), Y => 
        \N_RECD_SER_WORD[3]\);
    
    \Q[0]\ : DFN1C0
      port map(D => \ADJ_Q[0]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[0]_net_1\);
    
    \RECD_SER_WORD_RNO_0[7]\ : MX2
      port map(A => N_31, B => N_56, S => BIT_OS_SEL_5(1), Y => 
        N_64);
    
    \Q[7]\ : DFN1C0
      port map(D => \ADJ_Q[7]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[7]_net_1\);
    
    \ARB_BYTE[14]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[14]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[14]_net_1\);
    
    \ARB_WRD_40M_FIXED[2]\ : DFN1C0
      port map(D => \Q[2]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[2]_net_1\);
    
    \ARB_WRD_40M_FIXED[14]\ : DFN1C0
      port map(D => \Q[14]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[14]_net_1\);
    
    \RECD_SER_WORD_RNO[2]\ : MX2
      port map(A => N_35, B => N_36, S => BIT_OS_SEL_5(0), Y => 
        \N_RECD_SER_WORD[2]\);
    
    \ARB_BYTE_RNI04N31[1]\ : MX2
      port map(A => N_18, B => N_20, S => BIT_OS_SEL_3(1), Y => 
        N_34);
    
    \ARB_BYTE[2]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[2]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[2]_net_1\);
    
    \ADJ_Q[7]\ : DFN1C0
      port map(D => \ADJ_Q[5]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[7]_net_1\);
    
    \ARB_BYTE[8]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[8]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[8]_net_1\);
    
    \RECD_SER_WORD[5]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[5]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_8(5));
    
    \ARB_BYTE_RNINPQT[11]\ : MX2
      port map(A => N_22, B => N_24, S => BIT_OS_SEL_3(1), Y => 
        N_38);
    
    \ARB_BYTE[12]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[12]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[12]_net_1\);
    
    \RECD_SER_WORD[1]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[1]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_8(1));
    
    \ARB_BYTE_RNI8CN31[3]\ : MX2
      port map(A => N_20, B => N_22, S => BIT_OS_SEL_3(1), Y => 
        N_36);
    
    \Q[3]\ : DFN1C0
      port map(D => \ADJ_Q[3]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[3]_net_1\);
    
    \ARB_BYTE_RNIBU3H[3]\ : MX2
      port map(A => \ARB_BYTE[3]_net_1\, B => \ARB_BYTE[7]_net_1\, 
        S => BIT_OS_SEL_3(2), Y => N_20);
    
    ADJ_SER_IN_F_0DEL : DFN1C0
      port map(D => ELK_IN_F, CLK => CCC_160M_ADJ, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_F_0DEL\);
    
    \RECD_SER_WORD_RNO[7]\ : MX2
      port map(A => N_40, B => N_64, S => BIT_OS_SEL_5(0), Y => 
        \N_RECD_SER_WORD[7]\);
    
    \RECD_SER_WORD_RNO[1]\ : MX2
      port map(A => N_34, B => N_35, S => BIT_OS_SEL_5(0), Y => 
        \N_RECD_SER_WORD[1]\);
    
    \ARB_WRD_40M_FIXED[4]\ : DFN1C0
      port map(D => \Q[4]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[4]_net_1\);
    
    \RECD_SER_WORD_RNO[0]\ : MX2
      port map(A => N_33, B => N_34, S => BIT_OS_SEL_5(0), Y => 
        \N_RECD_SER_WORD[0]\);
    
    \Q[6]\ : DFN1C0
      port map(D => \ADJ_Q[6]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[6]_net_1\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \ARB_WRD_40M_FIXED[8]\ : DFN1C0
      port map(D => \Q[8]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[8]_net_1\);
    
    \ARB_BYTE[11]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[11]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[11]_net_1\);
    
    \Q[9]\ : DFN1C0
      port map(D => \ADJ_Q[9]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[9]_net_1\);
    
    \ARB_BYTE_RNIO97B[10]\ : MX2
      port map(A => \ARB_BYTE[6]_net_1\, B => 
        \ARB_BYTE[10]_net_1\, S => BIT_OS_SEL_3(2), Y => N_23);
    
    \Q[14]\ : DFN1C0
      port map(D => \ADJ_Q[14]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[14]_net_1\);
    
    ADJ_SER_IN_R_0DEL : DFN1C0
      port map(D => ELK_IN_R, CLK => CCC_160M_ADJ, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_R_0DEL\);
    
    \Q[13]\ : DFN1C0
      port map(D => \ADJ_Q[13]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[13]_net_1\);
    
    \ARB_BYTE[9]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[9]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[9]_net_1\);
    
    ADJ_SER_IN_R_1DEL : DFN1C0
      port map(D => \ADJ_SER_IN_R_0DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_R_1DEL\);
    
    \ARB_BYTE[10]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[10]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[10]_net_1\);
    
    \ADJ_Q[9]\ : DFN1C0
      port map(D => \ADJ_Q[7]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[9]_net_1\);
    
    \RECD_SER_WORD[7]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[7]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_8(7));
    
    \ARB_WRD_40M_FIXED[5]\ : DFN1C0
      port map(D => \Q[5]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[5]_net_1\);
    
    \ARB_WRD_40M_FIXED[12]\ : DFN1C0
      port map(D => \Q[12]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[12]_net_1\);
    
    \ARB_BYTE_RNID04H[4]\ : MX2
      port map(A => \ARB_BYTE[4]_net_1\, B => \ARB_BYTE[8]_net_1\, 
        S => BIT_OS_SEL_3(2), Y => N_21);
    
    \ARB_BYTE_RNI361P[10]\ : MX2
      port map(A => N_23, B => N_31, S => BIT_OS_SEL_3(1), Y => 
        N_39);
    
    \ARB_WRD_40M_FIXED[11]\ : DFN1C0
      port map(D => \Q[11]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[11]_net_1\);
    
    \ARB_WRD_40M_FIXED[0]\ : DFN1C0
      port map(D => \Q[0]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[0]_net_1\);
    
    \ADJ_Q[10]\ : DFN1C0
      port map(D => \ADJ_Q[8]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[10]_net_1\);
    
    \Q[2]\ : DFN1C0
      port map(D => \ADJ_Q[2]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[2]_net_1\);
    
    \ADJ_Q[1]\ : DFN1C0
      port map(D => \ADJ_SER_IN_F_1DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[1]_net_1\);
    
    \RECD_SER_WORD[6]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[6]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_8(6));
    
    \RECD_SER_WORD[2]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[2]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_8(2));
    
    \ADJ_Q[13]\ : DFN1C0
      port map(D => \ADJ_Q[11]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[13]_net_1\);
    
    \Q[8]\ : DFN1C0
      port map(D => \ADJ_Q[8]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[8]_net_1\);
    
    \ARB_BYTE_RNIQB7B[11]\ : MX2
      port map(A => \ARB_BYTE[7]_net_1\, B => 
        \ARB_BYTE[11]_net_1\, S => BIT_OS_SEL_3(2), Y => N_24);
    
    \ARB_BYTE[5]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[5]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[5]_net_1\);
    
    \ADJ_Q[14]\ : DFN1C0
      port map(D => \ADJ_Q[12]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[14]_net_1\);
    
    \RECD_SER_WORD_RNO[4]\ : MX2
      port map(A => N_37, B => N_38, S => BIT_OS_SEL_5(0), Y => 
        \N_RECD_SER_WORD[4]\);
    
    \Q[12]\ : DFN1C0
      port map(D => \ADJ_Q[12]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[12]_net_1\);
    
    \ARB_BYTE_RNI9S3H[2]\ : MX2
      port map(A => \ARB_BYTE[2]_net_1\, B => \ARB_BYTE[6]_net_1\, 
        S => BIT_OS_SEL_3(2), Y => N_19);
    
    \ARB_BYTE[13]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[13]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[13]_net_1\);
    
    \ARB_BYTE_RNIF24H[5]\ : MX2
      port map(A => \ARB_BYTE[5]_net_1\, B => \ARB_BYTE[9]_net_1\, 
        S => BIT_OS_SEL_3(2), Y => N_22);
    
    \ARB_WRD_40M_FIXED[3]\ : DFN1C0
      port map(D => \Q[3]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[3]_net_1\);
    
    \ARB_BYTE[7]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[7]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[7]_net_1\);
    
    \RECD_SER_WORD_RNO_0[0]\ : MX2
      port map(A => N_17, B => N_19, S => BIT_OS_SEL_3(1), Y => 
        N_33);
    
    \Q[4]\ : DFN1C0
      port map(D => \ADJ_Q[4]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[4]_net_1\);
    
    \ARB_WRD_40M_FIXED[7]\ : DFN1C0
      port map(D => \Q[7]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[7]_net_1\);
    
    \RECD_SER_WORD_RNO[6]\ : MX2
      port map(A => N_39, B => N_40, S => BIT_OS_SEL_5(0), Y => 
        \N_RECD_SER_WORD[6]\);
    
    \ARB_BYTE[3]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[3]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[3]_net_1\);
    
    \ARB_BYTE_RNIVIAC[13]\ : MX2
      port map(A => \ARB_BYTE[9]_net_1\, B => 
        \ARB_BYTE[13]_net_1\, S => BIT_OS_SEL_4_0, Y => N_32);
    
    \ADJ_Q[5]\ : DFN1C0
      port map(D => \ADJ_Q[3]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[5]_net_1\);
    
    \ARB_BYTE[1]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[1]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[1]_net_1\);
    
    \ARB_WRD_40M_FIXED[13]\ : DFN1C0
      port map(D => \Q[13]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[13]_net_1\);
    
    \ARB_BYTE_RNI48N31[2]\ : MX2
      port map(A => N_19, B => N_21, S => BIT_OS_SEL_3(1), Y => 
        N_35);
    
    \ADJ_Q[0]\ : DFN1C0
      port map(D => \ADJ_SER_IN_R_1DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[0]_net_1\);
    
    \ARB_WRD_40M_FIXED[10]\ : DFN1C0
      port map(D => \Q[10]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[10]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SER320M_3_34_8 is

    port( ELK_TX_DAT                 : in    std_logic_vector(7 downto 0);
          MASTER_SALT_POR_B_i_0_i_15 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i    : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_3  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_2  : in    std_logic;
          ELK_OUT_R                  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_5  : in    std_logic;
          ELK_OUT_F                  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_12 : in    std_logic;
          CCC_160M_FXD               : in    std_logic;
          CLK_40M_GL                 : in    std_logic
        );

end SER320M_3_34_8;

architecture DEF_ARCH of SER320M_3_34_8 is 

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \N_SER_CMD_WORD_R[0]\, \START_RISE\, 
        \N_SER_CMD_WORD_F[0]\, \N_SER_CMD_WORD_R[3]\, 
        \SER_CMD_WORD_R[2]_net_1\, \N_SER_CMD_WORD_R[2]\, 
        \SER_CMD_WORD_R[1]_net_1\, \N_SER_CMD_WORD_R[1]\, 
        \SER_CMD_WORD_R[0]_net_1\, \N_SER_CMD_WORD_F[3]\, 
        \SER_CMD_WORD_F[2]_net_1\, \N_SER_CMD_WORD_F[2]\, 
        \SER_CMD_WORD_F[1]_net_1\, \N_SER_CMD_WORD_F[1]\, 
        \SER_CMD_WORD_F[0]_net_1\, N_START_RISE, 
        \CLK40M_GEN_DEL0\, \SER_OUT_FI\, \SER_OUT_RI\, 
        \SER_CMD_WORD_F[3]_net_1\, \SER_CMD_WORD_R[3]_net_1\, 
        \GND\, \VCC\ : std_logic;

begin 


    SER_OUT_FI : DFN1C0
      port map(D => \SER_CMD_WORD_F[3]_net_1\, CLK => 
        CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_3, Q => 
        \SER_OUT_FI\);
    
    \SER_CMD_WORD_F[3]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[3]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i, Q => 
        \SER_CMD_WORD_F[3]_net_1\);
    
    \SER_CMD_WORD_R[1]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[1]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_15, Q => 
        \SER_CMD_WORD_R[1]_net_1\);
    
    \SER_CMD_WORD_R[2]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[2]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_15, Q => 
        \SER_CMD_WORD_R[2]_net_1\);
    
    \SER_CMD_WORD_R_RNO[3]\ : MX2
      port map(A => \SER_CMD_WORD_R[2]_net_1\, B => ELK_TX_DAT(7), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_R[3]\);
    
    \SER_CMD_WORD_R_RNO[0]\ : NOR2B
      port map(A => \START_RISE\, B => ELK_TX_DAT(1), Y => 
        \N_SER_CMD_WORD_R[0]\);
    
    \SER_CMD_WORD_F[0]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[0]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i, Q => 
        \SER_CMD_WORD_F[0]_net_1\);
    
    \SER_CMD_WORD_R_RNO[1]\ : MX2
      port map(A => \SER_CMD_WORD_R[0]_net_1\, B => ELK_TX_DAT(3), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_R[1]\);
    
    \SER_CMD_WORD_F_RNO[2]\ : MX2
      port map(A => \SER_CMD_WORD_F[1]_net_1\, B => ELK_TX_DAT(4), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_F[2]\);
    
    \SER_CMD_WORD_F_RNO[3]\ : MX2
      port map(A => \SER_CMD_WORD_F[2]_net_1\, B => ELK_TX_DAT(6), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_F[3]\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    CLK40M_GEN_DEL0 : DFN1C0
      port map(D => CLK_40M_GL, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_12, Q => \CLK40M_GEN_DEL0\);
    
    SER_OUT_RI : DFN1C0
      port map(D => \SER_CMD_WORD_R[3]_net_1\, CLK => 
        CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_3, Q => 
        \SER_OUT_RI\);
    
    \SER_CMD_WORD_F[2]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[2]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i, Q => 
        \SER_CMD_WORD_F[2]_net_1\);
    
    \SER_CMD_WORD_F_RNO[1]\ : MX2
      port map(A => \SER_CMD_WORD_F[0]_net_1\, B => ELK_TX_DAT(2), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_F[1]\);
    
    \SER_CMD_WORD_R[0]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[0]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_15, Q => 
        \SER_CMD_WORD_R[0]_net_1\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    START_RISE : DFN1C0
      port map(D => N_START_RISE, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_12, Q => \START_RISE\);
    
    \SER_CMD_WORD_R[3]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[3]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_15, Q => 
        \SER_CMD_WORD_R[3]_net_1\);
    
    \SER_CMD_WORD_F_RNO[0]\ : NOR2B
      port map(A => \START_RISE\, B => ELK_TX_DAT(0), Y => 
        \N_SER_CMD_WORD_F[0]\);
    
    SER_OUT_RDEL : DFN1C0
      port map(D => \SER_OUT_RI\, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_2, Q => ELK_OUT_R);
    
    \SER_CMD_WORD_F[1]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[1]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i, Q => 
        \SER_CMD_WORD_F[1]_net_1\);
    
    START_RISE_RNO : NOR2B
      port map(A => \CLK40M_GEN_DEL0\, B => CLK_40M_GL, Y => 
        N_START_RISE);
    
    \SER_CMD_WORD_R_RNO[2]\ : MX2
      port map(A => \SER_CMD_WORD_R[1]_net_1\, B => ELK_TX_DAT(5), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_R[2]\);
    
    SER_OUT_FDEL : DFN1C0
      port map(D => \SER_OUT_FI\, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_5, Q => ELK_OUT_F);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity DDR_BIDIR_LVDS_DUAL_CLK_8 is

    port( DCB_SALT_SEL_c_i : in    std_logic;
          ELK8_DAT_P       : inout std_logic := 'Z';
          ELK8_DAT_N       : inout std_logic := 'Z';
          ELK_OUT_R        : in    std_logic;
          ELK_OUT_F        : in    std_logic;
          CCC_160M_FXD     : in    std_logic;
          CCC_160M_ADJ     : in    std_logic;
          ELK_IN_DDR_R     : out   std_logic;
          ELK_IN_DDR_F     : out   std_logic
        );

end DDR_BIDIR_LVDS_DUAL_CLK_8;

architecture DEF_ARCH of DDR_BIDIR_LVDS_DUAL_CLK_8 is 

  component DDR_REG
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          QR  : out   std_logic;
          QF  : out   std_logic
        );
  end component;

  component DDR_OUT
    port( DR  : in    std_logic := 'U';
          DF  : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component BIBUF_LVDS
    port( PADP : inout   std_logic;
          PADN : inout   std_logic;
          D    : in    std_logic := 'U';
          E    : in    std_logic := 'U';
          Y    : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal DDR_BIDIR_LVDS_DUAL_CLK_8_GND, BIBUF_LVDS_0_Y, 
        DDR_OUT_0_Q, \VCC\ : std_logic;

begin 


    DDR_REG_0 : DDR_REG
      port map(D => BIBUF_LVDS_0_Y, CLK => CCC_160M_ADJ, CLR => 
        DDR_BIDIR_LVDS_DUAL_CLK_8_GND, QR => ELK_IN_DDR_R, QF => 
        ELK_IN_DDR_F);
    
    DDR_OUT_0 : DDR_OUT
      port map(DR => ELK_OUT_R, DF => ELK_OUT_F, CLK => 
        CCC_160M_FXD, CLR => DDR_BIDIR_LVDS_DUAL_CLK_8_GND, Q => 
        DDR_OUT_0_Q);
    
    BIBUF_LVDS_0 : BIBUF_LVDS
      port map(PADP => ELK8_DAT_P, PADN => ELK8_DAT_N, D => 
        DDR_OUT_0_Q, E => DCB_SALT_SEL_c_i, Y => BIBUF_LVDS_0_Y);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    GND_i : GND
      port map(Y => DDR_BIDIR_LVDS_DUAL_CLK_8_GND);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SYNC_DAT_SEL_8 is

    port( ELK_TX_DAT                : out   std_logic_vector(7 downto 0);
          PATT_ELK_DAT_8            : in    std_logic_vector(7 downto 0);
          OP_MODE_c_0_0             : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_5 : in    std_logic;
          CLK_40M_GL                : in    std_logic
        );

end SYNC_DAT_SEL_8;

architecture DEF_ARCH of SYNC_DAT_SEL_8 is 

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \N_SERDAT[0]\, \N_SERDAT[1]\, \N_SERDAT[2]\, 
        \N_SERDAT[3]\, \N_SERDAT[4]\, \N_SERDAT[5]\, 
        \N_SERDAT[6]\, \N_SERDAT[7]\, \GND\, \VCC\ : std_logic;

begin 


    \SERDAT_RNO[4]\ : NOR2A
      port map(A => PATT_ELK_DAT_8(4), B => OP_MODE_c_0_0, Y => 
        \N_SERDAT[4]\);
    
    \SERDAT_RNO[0]\ : NOR2A
      port map(A => PATT_ELK_DAT_8(0), B => OP_MODE_c_0_0, Y => 
        \N_SERDAT[0]\);
    
    \SERDAT[6]\ : DFN1C0
      port map(D => \N_SERDAT[6]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_5, Q => ELK_TX_DAT(6));
    
    \SERDAT[4]\ : DFN1C0
      port map(D => \N_SERDAT[4]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_5, Q => ELK_TX_DAT(4));
    
    \SERDAT_RNO[7]\ : OR2
      port map(A => PATT_ELK_DAT_8(7), B => OP_MODE_c_0_0, Y => 
        \N_SERDAT[7]\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \SERDAT_RNO[3]\ : OR2
      port map(A => PATT_ELK_DAT_8(3), B => OP_MODE_c_0_0, Y => 
        \N_SERDAT[3]\);
    
    \SERDAT_RNO[2]\ : OR2
      port map(A => PATT_ELK_DAT_8(2), B => OP_MODE_c_0_0, Y => 
        \N_SERDAT[2]\);
    
    \SERDAT[5]\ : DFN1C0
      port map(D => \N_SERDAT[5]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_5, Q => ELK_TX_DAT(5));
    
    \SERDAT[7]\ : DFN1C0
      port map(D => \N_SERDAT[7]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_5, Q => ELK_TX_DAT(7));
    
    GND_i : GND
      port map(Y => \GND\);
    
    \SERDAT_RNO[5]\ : NOR2A
      port map(A => PATT_ELK_DAT_8(5), B => OP_MODE_c_0_0, Y => 
        \N_SERDAT[5]\);
    
    \SERDAT[0]\ : DFN1C0
      port map(D => \N_SERDAT[0]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_5, Q => ELK_TX_DAT(0));
    
    \SERDAT_RNO[6]\ : NOR2A
      port map(A => PATT_ELK_DAT_8(6), B => OP_MODE_c_0_0, Y => 
        \N_SERDAT[6]\);
    
    \SERDAT[1]\ : DFN1C0
      port map(D => \N_SERDAT[1]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_5, Q => ELK_TX_DAT(1));
    
    \SERDAT_RNO[1]\ : OR2
      port map(A => PATT_ELK_DAT_8(1), B => OP_MODE_c_0_0, Y => 
        \N_SERDAT[1]\);
    
    \SERDAT[3]\ : DFN1C0
      port map(D => \N_SERDAT[3]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_5, Q => ELK_TX_DAT(3));
    
    \SERDAT[2]\ : DFN1C0
      port map(D => \N_SERDAT[2]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_5, Q => ELK_TX_DAT(2));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity ELINK_SLAVE_15_3 is

    port( BIT_OS_SEL_4_0             : in    std_logic;
          BIT_OS_SEL_3               : in    std_logic_vector(2 downto 1);
          BIT_OS_SEL_6_0             : in    std_logic;
          BIT_OS_SEL_5               : in    std_logic_vector(1 downto 0);
          ELK_RX_SER_WORD_8          : out   std_logic_vector(7 downto 0);
          OP_MODE_c_0_0              : in    std_logic;
          PATT_ELK_DAT_8             : in    std_logic_vector(7 downto 0);
          MASTER_DCB_POR_B_i_0_i     : in    std_logic;
          ELK8_DAT_N                 : inout std_logic := 'Z';
          ELK8_DAT_P                 : inout std_logic := 'Z';
          DCB_SALT_SEL_c_i           : in    std_logic;
          CCC_160M_FXD               : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_12 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_2  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_3  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i    : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_15 : in    std_logic;
          CLK_40M_GL                 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_5  : in    std_logic;
          DEV_RST_B_c_1              : in    std_logic;
          DEV_RST_B_c_0              : in    std_logic;
          CCC_160M_ADJ               : in    std_logic
        );

end ELINK_SLAVE_15_3;

architecture DEF_ARCH of ELINK_SLAVE_15_3 is 

  component SLAVE_DES320S_1_17_6
    port( ELK_RX_SER_WORD_8      : out   std_logic_vector(7 downto 0);
          BIT_OS_SEL_5           : in    std_logic_vector(1 downto 0) := (others => 'U');
          BIT_OS_SEL_6_0         : in    std_logic := 'U';
          BIT_OS_SEL_3           : in    std_logic_vector(2 downto 1) := (others => 'U');
          BIT_OS_SEL_4_0         : in    std_logic := 'U';
          CLK_40M_GL             : in    std_logic := 'U';
          CCC_160M_FXD           : in    std_logic := 'U';
          ELK_IN_R               : in    std_logic := 'U';
          ELK_IN_F               : in    std_logic := 'U';
          MASTER_DCB_POR_B_i_0_i : in    std_logic := 'U';
          CCC_160M_ADJ           : in    std_logic := 'U'
        );
  end component;

  component SER320M_3_34_8
    port( ELK_TX_DAT                 : in    std_logic_vector(7 downto 0) := (others => 'U');
          MASTER_SALT_POR_B_i_0_i_15 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i    : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_3  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_2  : in    std_logic := 'U';
          ELK_OUT_R                  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_5  : in    std_logic := 'U';
          ELK_OUT_F                  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_12 : in    std_logic := 'U';
          CCC_160M_FXD               : in    std_logic := 'U';
          CLK_40M_GL                 : in    std_logic := 'U'
        );
  end component;

  component DDR_BIDIR_LVDS_DUAL_CLK_8
    port( DCB_SALT_SEL_c_i : in    std_logic := 'U';
          ELK8_DAT_P       : inout   std_logic;
          ELK8_DAT_N       : inout   std_logic;
          ELK_OUT_R        : in    std_logic := 'U';
          ELK_OUT_F        : in    std_logic := 'U';
          CCC_160M_FXD     : in    std_logic := 'U';
          CCC_160M_ADJ     : in    std_logic := 'U';
          ELK_IN_DDR_R     : out   std_logic;
          ELK_IN_DDR_F     : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component SYNC_DAT_SEL_8
    port( ELK_TX_DAT                : out   std_logic_vector(7 downto 0);
          PATT_ELK_DAT_8            : in    std_logic_vector(7 downto 0) := (others => 'U');
          OP_MODE_c_0_0             : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_5 : in    std_logic := 'U';
          CLK_40M_GL                : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \ELK_IN_F\, ELK_IN_DDR_F, \ELK_IN_R\, ELK_IN_DDR_R, 
        \ELK_TX_DAT[0]\, \ELK_TX_DAT[1]\, \ELK_TX_DAT[2]\, 
        \ELK_TX_DAT[3]\, \ELK_TX_DAT[4]\, \ELK_TX_DAT[5]\, 
        \ELK_TX_DAT[6]\, \ELK_TX_DAT[7]\, ELK_OUT_R, ELK_OUT_F, 
        \GND\, \VCC\ : std_logic;

    for all : SLAVE_DES320S_1_17_6
	Use entity work.SLAVE_DES320S_1_17_6(DEF_ARCH);
    for all : SER320M_3_34_8
	Use entity work.SER320M_3_34_8(DEF_ARCH);
    for all : DDR_BIDIR_LVDS_DUAL_CLK_8
	Use entity work.DDR_BIDIR_LVDS_DUAL_CLK_8(DEF_ARCH);
    for all : SYNC_DAT_SEL_8
	Use entity work.SYNC_DAT_SEL_8(DEF_ARCH);
begin 


    U_SLAVE_1ELK : SLAVE_DES320S_1_17_6
      port map(ELK_RX_SER_WORD_8(7) => ELK_RX_SER_WORD_8(7), 
        ELK_RX_SER_WORD_8(6) => ELK_RX_SER_WORD_8(6), 
        ELK_RX_SER_WORD_8(5) => ELK_RX_SER_WORD_8(5), 
        ELK_RX_SER_WORD_8(4) => ELK_RX_SER_WORD_8(4), 
        ELK_RX_SER_WORD_8(3) => ELK_RX_SER_WORD_8(3), 
        ELK_RX_SER_WORD_8(2) => ELK_RX_SER_WORD_8(2), 
        ELK_RX_SER_WORD_8(1) => ELK_RX_SER_WORD_8(1), 
        ELK_RX_SER_WORD_8(0) => ELK_RX_SER_WORD_8(0), 
        BIT_OS_SEL_5(1) => BIT_OS_SEL_5(1), BIT_OS_SEL_5(0) => 
        BIT_OS_SEL_5(0), BIT_OS_SEL_6_0 => BIT_OS_SEL_6_0, 
        BIT_OS_SEL_3(2) => BIT_OS_SEL_3(2), BIT_OS_SEL_3(1) => 
        BIT_OS_SEL_3(1), BIT_OS_SEL_4_0 => BIT_OS_SEL_4_0, 
        CLK_40M_GL => CLK_40M_GL, CCC_160M_FXD => CCC_160M_FXD, 
        ELK_IN_R => \ELK_IN_R\, ELK_IN_F => \ELK_IN_F\, 
        MASTER_DCB_POR_B_i_0_i => MASTER_DCB_POR_B_i_0_i, 
        CCC_160M_ADJ => CCC_160M_ADJ);
    
    U_ELK1_CMD_TX : SER320M_3_34_8
      port map(ELK_TX_DAT(7) => \ELK_TX_DAT[7]\, ELK_TX_DAT(6)
         => \ELK_TX_DAT[6]\, ELK_TX_DAT(5) => \ELK_TX_DAT[5]\, 
        ELK_TX_DAT(4) => \ELK_TX_DAT[4]\, ELK_TX_DAT(3) => 
        \ELK_TX_DAT[3]\, ELK_TX_DAT(2) => \ELK_TX_DAT[2]\, 
        ELK_TX_DAT(1) => \ELK_TX_DAT[1]\, ELK_TX_DAT(0) => 
        \ELK_TX_DAT[0]\, MASTER_SALT_POR_B_i_0_i_15 => 
        MASTER_SALT_POR_B_i_0_i_15, MASTER_SALT_POR_B_i_0_i => 
        MASTER_SALT_POR_B_i_0_i, MASTER_SALT_POR_B_i_0_i_3 => 
        MASTER_SALT_POR_B_i_0_i_3, MASTER_SALT_POR_B_i_0_i_2 => 
        MASTER_SALT_POR_B_i_0_i_2, ELK_OUT_R => ELK_OUT_R, 
        MASTER_SALT_POR_B_i_0_i_5 => MASTER_SALT_POR_B_i_0_i_5, 
        ELK_OUT_F => ELK_OUT_F, MASTER_SALT_POR_B_i_0_i_12 => 
        MASTER_SALT_POR_B_i_0_i_12, CCC_160M_FXD => CCC_160M_FXD, 
        CLK_40M_GL => CLK_40M_GL);
    
    U_DDR_ELK1 : DDR_BIDIR_LVDS_DUAL_CLK_8
      port map(DCB_SALT_SEL_c_i => DCB_SALT_SEL_c_i, ELK8_DAT_P
         => ELK8_DAT_P, ELK8_DAT_N => ELK8_DAT_N, ELK_OUT_R => 
        ELK_OUT_R, ELK_OUT_F => ELK_OUT_F, CCC_160M_FXD => 
        CCC_160M_FXD, CCC_160M_ADJ => CCC_160M_ADJ, ELK_IN_DDR_R
         => ELK_IN_DDR_R, ELK_IN_DDR_F => ELK_IN_DDR_F);
    
    ELK_IN_F : DFN1C0
      port map(D => ELK_IN_DDR_F, CLK => CCC_160M_ADJ, CLR => 
        DEV_RST_B_c_0, Q => \ELK_IN_F\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    U_ELK1_SERDAT_SOURCE : SYNC_DAT_SEL_8
      port map(ELK_TX_DAT(7) => \ELK_TX_DAT[7]\, ELK_TX_DAT(6)
         => \ELK_TX_DAT[6]\, ELK_TX_DAT(5) => \ELK_TX_DAT[5]\, 
        ELK_TX_DAT(4) => \ELK_TX_DAT[4]\, ELK_TX_DAT(3) => 
        \ELK_TX_DAT[3]\, ELK_TX_DAT(2) => \ELK_TX_DAT[2]\, 
        ELK_TX_DAT(1) => \ELK_TX_DAT[1]\, ELK_TX_DAT(0) => 
        \ELK_TX_DAT[0]\, PATT_ELK_DAT_8(7) => PATT_ELK_DAT_8(7), 
        PATT_ELK_DAT_8(6) => PATT_ELK_DAT_8(6), PATT_ELK_DAT_8(5)
         => PATT_ELK_DAT_8(5), PATT_ELK_DAT_8(4) => 
        PATT_ELK_DAT_8(4), PATT_ELK_DAT_8(3) => PATT_ELK_DAT_8(3), 
        PATT_ELK_DAT_8(2) => PATT_ELK_DAT_8(2), PATT_ELK_DAT_8(1)
         => PATT_ELK_DAT_8(1), PATT_ELK_DAT_8(0) => 
        PATT_ELK_DAT_8(0), OP_MODE_c_0_0 => OP_MODE_c_0_0, 
        MASTER_SALT_POR_B_i_0_i_5 => MASTER_SALT_POR_B_i_0_i_5, 
        CLK_40M_GL => CLK_40M_GL);
    
    ELK_IN_R : DFN1C0
      port map(D => ELK_IN_DDR_R, CLK => CCC_160M_ADJ, CLR => 
        DEV_RST_B_c_1, Q => \ELK_IN_R\);
    
    GND_i : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SLAVE_DES320S_1_17_15 is

    port( ELK_RX_SER_WORD_17     : out   std_logic_vector(7 downto 0);
          BIT_OS_SEL_3_0         : in    std_logic;
          BIT_OS_SEL_2           : in    std_logic_vector(2 downto 0);
          BIT_OS_SEL_1_0         : in    std_logic;
          BIT_OS_SEL_0_0         : in    std_logic;
          CLK_40M_GL             : in    std_logic;
          CCC_160M_FXD           : in    std_logic;
          ELK_IN_R               : in    std_logic;
          ELK_IN_F               : in    std_logic;
          MASTER_DCB_POR_B_i_0_i : in    std_logic;
          CCC_160M_ADJ           : in    std_logic
        );

end SLAVE_DES320S_1_17_15;

architecture DEF_ARCH of SLAVE_DES320S_1_17_15 is 

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal N_17, \ARB_BYTE[0]_net_1\, \ARB_BYTE[4]_net_1\, N_18, 
        \ARB_BYTE[1]_net_1\, \ARB_BYTE[5]_net_1\, N_19, 
        \ARB_BYTE[2]_net_1\, \ARB_BYTE[6]_net_1\, N_20, 
        \ARB_BYTE[3]_net_1\, \ARB_BYTE[7]_net_1\, N_21, 
        \ARB_BYTE[8]_net_1\, N_22, \ARB_BYTE[9]_net_1\, N_23, 
        \ARB_BYTE[10]_net_1\, N_24, \ARB_BYTE[11]_net_1\, N_31, 
        \ARB_BYTE[12]_net_1\, N_32, \ARB_BYTE[13]_net_1\, N_33, 
        N_34, N_35, N_36, N_37, N_38, N_39, N_40, N_56, 
        \ARB_BYTE[14]_net_1\, N_64, \N_RECD_SER_WORD[0]\, 
        \N_RECD_SER_WORD[1]\, \N_RECD_SER_WORD[2]\, 
        \N_RECD_SER_WORD[3]\, \N_RECD_SER_WORD[4]\, 
        \N_RECD_SER_WORD[5]\, \N_RECD_SER_WORD[6]\, 
        \N_RECD_SER_WORD[7]\, \ADJ_SER_IN_F_0DEL\, 
        \ADJ_SER_IN_R_0DEL\, \ADJ_SER_IN_F_1DEL\, 
        \ADJ_SER_IN_R_1DEL\, \Q[0]_net_1\, \ADJ_Q[0]_net_1\, 
        \Q[1]_net_1\, \ADJ_Q[1]_net_1\, \Q[2]_net_1\, 
        \ADJ_Q[2]_net_1\, \Q[3]_net_1\, \ADJ_Q[3]_net_1\, 
        \Q[4]_net_1\, \ADJ_Q[4]_net_1\, \Q[5]_net_1\, 
        \ADJ_Q[5]_net_1\, \Q[6]_net_1\, \ADJ_Q[6]_net_1\, 
        \Q[7]_net_1\, \ADJ_Q[7]_net_1\, \Q[8]_net_1\, 
        \ADJ_Q[8]_net_1\, \Q[9]_net_1\, \ADJ_Q[9]_net_1\, 
        \Q[10]_net_1\, \ADJ_Q[10]_net_1\, \Q[11]_net_1\, 
        \ADJ_Q[11]_net_1\, \Q[12]_net_1\, \ADJ_Q[12]_net_1\, 
        \Q[13]_net_1\, \ADJ_Q[13]_net_1\, \Q[14]_net_1\, 
        \ADJ_Q[14]_net_1\, \ARB_WRD_40M_FIXED[0]_net_1\, 
        \ARB_WRD_40M_FIXED[1]_net_1\, 
        \ARB_WRD_40M_FIXED[2]_net_1\, 
        \ARB_WRD_40M_FIXED[3]_net_1\, 
        \ARB_WRD_40M_FIXED[4]_net_1\, 
        \ARB_WRD_40M_FIXED[5]_net_1\, 
        \ARB_WRD_40M_FIXED[6]_net_1\, 
        \ARB_WRD_40M_FIXED[7]_net_1\, 
        \ARB_WRD_40M_FIXED[8]_net_1\, 
        \ARB_WRD_40M_FIXED[9]_net_1\, 
        \ARB_WRD_40M_FIXED[10]_net_1\, 
        \ARB_WRD_40M_FIXED[11]_net_1\, 
        \ARB_WRD_40M_FIXED[12]_net_1\, 
        \ARB_WRD_40M_FIXED[13]_net_1\, 
        \ARB_WRD_40M_FIXED[14]_net_1\, \GND\, \VCC\ : std_logic;

begin 


    \RECD_SER_WORD_RNO[5]\ : MX2
      port map(A => N_38, B => N_39, S => BIT_OS_SEL_3_0, Y => 
        \N_RECD_SER_WORD[5]\);
    
    \ARB_WRD_40M_FIXED[9]\ : DFN1C0
      port map(D => \Q[9]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[9]_net_1\);
    
    \ADJ_Q[4]\ : DFN1C0
      port map(D => \ADJ_Q[2]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[4]_net_1\);
    
    \ARB_BYTE[6]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[6]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[6]_net_1\);
    
    ADJ_SER_IN_F_1DEL : DFN1C0
      port map(D => \ADJ_SER_IN_F_0DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_F_1DEL\);
    
    \ARB_BYTE[0]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[0]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[0]_net_1\);
    
    \Q[11]\ : DFN1C0
      port map(D => \ADJ_Q[11]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[11]_net_1\);
    
    \ADJ_Q[8]\ : DFN1C0
      port map(D => \ADJ_Q[6]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[8]_net_1\);
    
    \ADJ_Q[6]\ : DFN1C0
      port map(D => \ADJ_Q[4]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[6]_net_1\);
    
    \ADJ_Q[12]\ : DFN1C0
      port map(D => \ADJ_Q[10]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[12]_net_1\);
    
    \RECD_SER_WORD_RNO_1[0]\ : MX2
      port map(A => \ARB_BYTE[0]_net_1\, B => \ARB_BYTE[4]_net_1\, 
        S => BIT_OS_SEL_0_0, Y => N_17);
    
    \Q[1]\ : DFN1C0
      port map(D => \ADJ_Q[1]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[1]_net_1\);
    
    \ARB_BYTE[4]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[4]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[4]_net_1\);
    
    \ADJ_Q[2]\ : DFN1C0
      port map(D => \ADJ_Q[0]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[2]_net_1\);
    
    \RECD_SER_WORD_RNO_1[7]\ : MX2
      port map(A => \ARB_BYTE[10]_net_1\, B => 
        \ARB_BYTE[14]_net_1\, S => BIT_OS_SEL_2(2), Y => N_56);
    
    \RECD_SER_WORD[4]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[4]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_17(4));
    
    \Q[5]\ : DFN1C0
      port map(D => \ADJ_Q[5]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[5]_net_1\);
    
    \ADJ_Q[11]\ : DFN1C0
      port map(D => \ADJ_Q[9]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[11]_net_1\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \ARB_BYTE_RNIQKMA2[6]\ : MX2
      port map(A => N_23, B => N_31, S => BIT_OS_SEL_1_0, Y => 
        N_39);
    
    \ADJ_Q[3]\ : DFN1C0
      port map(D => \ADJ_Q[1]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[3]_net_1\);
    
    \Q[10]\ : DFN1C0
      port map(D => \ADJ_Q[10]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[10]_net_1\);
    
    \ARB_WRD_40M_FIXED[6]\ : DFN1C0
      port map(D => \Q[6]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[6]_net_1\);
    
    \ARB_WRD_40M_FIXED[1]\ : DFN1C0
      port map(D => \Q[1]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[1]_net_1\);
    
    \ARB_BYTE_RNIRRMT[13]\ : MX2
      port map(A => \ARB_BYTE[9]_net_1\, B => 
        \ARB_BYTE[13]_net_1\, S => BIT_OS_SEL_0_0, Y => N_32);
    
    \RECD_SER_WORD[3]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[3]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_17(3));
    
    \RECD_SER_WORD[0]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[0]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_17(0));
    
    \RECD_SER_WORD_RNO[3]\ : MX2
      port map(A => N_36, B => N_37, S => BIT_OS_SEL_3_0, Y => 
        \N_RECD_SER_WORD[3]\);
    
    \Q[0]\ : DFN1C0
      port map(D => \ADJ_Q[0]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[0]_net_1\);
    
    \ARB_BYTE_RNI0UA02[3]\ : MX2
      port map(A => N_20, B => N_22, S => BIT_OS_SEL_1_0, Y => 
        N_36);
    
    \ARB_BYTE_RNIFRG52[5]\ : MX2
      port map(A => N_22, B => N_24, S => BIT_OS_SEL_1_0, Y => 
        N_38);
    
    \RECD_SER_WORD_RNO_0[7]\ : MX2
      port map(A => N_31, B => N_56, S => BIT_OS_SEL_2(1), Y => 
        N_64);
    
    \Q[7]\ : DFN1C0
      port map(D => \ADJ_Q[7]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[7]_net_1\);
    
    \ARB_BYTE[14]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[14]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[14]_net_1\);
    
    \ARB_WRD_40M_FIXED[2]\ : DFN1C0
      port map(D => \Q[2]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[2]_net_1\);
    
    \ARB_WRD_40M_FIXED[14]\ : DFN1C0
      port map(D => \Q[14]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[14]_net_1\);
    
    \RECD_SER_WORD_RNO[2]\ : MX2
      port map(A => N_35, B => N_36, S => BIT_OS_SEL_3_0, Y => 
        \N_RECD_SER_WORD[2]\);
    
    \ARB_BYTE_RNI6OGO[2]\ : MX2
      port map(A => \ARB_BYTE[2]_net_1\, B => \ARB_BYTE[6]_net_1\, 
        S => BIT_OS_SEL_0_0, Y => N_19);
    
    \ARB_BYTE[2]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[2]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[2]_net_1\);
    
    \ARB_BYTE_RNIPPMT[12]\ : MX2
      port map(A => \ARB_BYTE[8]_net_1\, B => 
        \ARB_BYTE[12]_net_1\, S => BIT_OS_SEL_0_0, Y => N_31);
    
    \ADJ_Q[7]\ : DFN1C0
      port map(D => \ADJ_Q[5]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[7]_net_1\);
    
    \ARB_BYTE[8]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[8]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[8]_net_1\);
    
    \RECD_SER_WORD[5]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[5]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_17(5));
    
    \ARB_BYTE[12]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[12]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[12]_net_1\);
    
    \ARB_BYTE_RNIUOMA2[13]\ : MX2
      port map(A => N_24, B => N_32, S => BIT_OS_SEL_1_0, Y => 
        N_40);
    
    \RECD_SER_WORD[1]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[1]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_17(1));
    
    \Q[3]\ : DFN1C0
      port map(D => \ADJ_Q[3]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[3]_net_1\);
    
    ADJ_SER_IN_F_0DEL : DFN1C0
      port map(D => ELK_IN_F, CLK => CCC_160M_ADJ, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_F_0DEL\);
    
    \RECD_SER_WORD_RNO[7]\ : MX2
      port map(A => N_40, B => N_64, S => BIT_OS_SEL_3_0, Y => 
        \N_RECD_SER_WORD[7]\);
    
    \RECD_SER_WORD_RNO[1]\ : MX2
      port map(A => N_34, B => N_35, S => BIT_OS_SEL_2(0), Y => 
        \N_RECD_SER_WORD[1]\);
    
    \ARB_WRD_40M_FIXED[4]\ : DFN1C0
      port map(D => \Q[4]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[4]_net_1\);
    
    \ARB_BYTE_RNI4MGO[1]\ : MX2
      port map(A => \ARB_BYTE[1]_net_1\, B => \ARB_BYTE[5]_net_1\, 
        S => BIT_OS_SEL_0_0, Y => N_18);
    
    \RECD_SER_WORD_RNO[0]\ : MX2
      port map(A => N_33, B => N_34, S => BIT_OS_SEL_2(0), Y => 
        \N_RECD_SER_WORD[0]\);
    
    \Q[6]\ : DFN1C0
      port map(D => \ADJ_Q[6]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[6]_net_1\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \ARB_WRD_40M_FIXED[8]\ : DFN1C0
      port map(D => \Q[8]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[8]_net_1\);
    
    \ARB_BYTE[11]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[11]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[11]_net_1\);
    
    \Q[9]\ : DFN1C0
      port map(D => \ADJ_Q[9]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[9]_net_1\);
    
    \ARB_BYTE_RNISPA02[2]\ : MX2
      port map(A => N_19, B => N_21, S => BIT_OS_SEL_1_0, Y => 
        N_35);
    
    \Q[14]\ : DFN1C0
      port map(D => \ADJ_Q[14]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[14]_net_1\);
    
    ADJ_SER_IN_R_0DEL : DFN1C0
      port map(D => ELK_IN_R, CLK => CCC_160M_ADJ, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_R_0DEL\);
    
    \Q[13]\ : DFN1C0
      port map(D => \ADJ_Q[13]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[13]_net_1\);
    
    \ARB_BYTE[9]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[9]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[9]_net_1\);
    
    ADJ_SER_IN_R_1DEL : DFN1C0
      port map(D => \ADJ_SER_IN_R_0DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_R_1DEL\);
    
    \ARB_BYTE[10]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[10]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[10]_net_1\);
    
    \ADJ_Q[9]\ : DFN1C0
      port map(D => \ADJ_Q[7]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[9]_net_1\);
    
    \RECD_SER_WORD[7]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[7]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_17(7));
    
    \ARB_WRD_40M_FIXED[5]\ : DFN1C0
      port map(D => \Q[5]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[5]_net_1\);
    
    \ARB_WRD_40M_FIXED[12]\ : DFN1C0
      port map(D => \Q[12]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[12]_net_1\);
    
    \ARB_BYTE_RNICUGO[5]\ : MX2
      port map(A => \ARB_BYTE[5]_net_1\, B => \ARB_BYTE[9]_net_1\, 
        S => BIT_OS_SEL_0_0, Y => N_22);
    
    \ARB_BYTE_RNIASGO[4]\ : MX2
      port map(A => \ARB_BYTE[4]_net_1\, B => \ARB_BYTE[8]_net_1\, 
        S => BIT_OS_SEL_0_0, Y => N_21);
    
    \ARB_WRD_40M_FIXED[11]\ : DFN1C0
      port map(D => \Q[11]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[11]_net_1\);
    
    \ARB_WRD_40M_FIXED[0]\ : DFN1C0
      port map(D => \Q[0]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[0]_net_1\);
    
    \ADJ_Q[10]\ : DFN1C0
      port map(D => \ADJ_Q[8]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[10]_net_1\);
    
    \Q[2]\ : DFN1C0
      port map(D => \ADJ_Q[2]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[2]_net_1\);
    
    \ADJ_Q[1]\ : DFN1C0
      port map(D => \ADJ_SER_IN_F_1DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[1]_net_1\);
    
    \RECD_SER_WORD[6]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[6]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_17(6));
    
    \RECD_SER_WORD[2]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[2]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_17(2));
    
    \ADJ_Q[13]\ : DFN1C0
      port map(D => \ADJ_Q[11]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[13]_net_1\);
    
    \Q[8]\ : DFN1C0
      port map(D => \ADJ_Q[8]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[8]_net_1\);
    
    \ARB_BYTE[5]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[5]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[5]_net_1\);
    
    \ADJ_Q[14]\ : DFN1C0
      port map(D => \ADJ_Q[12]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[14]_net_1\);
    
    \RECD_SER_WORD_RNO[4]\ : MX2
      port map(A => N_37, B => N_38, S => BIT_OS_SEL_3_0, Y => 
        \N_RECD_SER_WORD[4]\);
    
    \Q[12]\ : DFN1C0
      port map(D => \ADJ_Q[12]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[12]_net_1\);
    
    \ARB_BYTE[13]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[13]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[13]_net_1\);
    
    \ARB_WRD_40M_FIXED[3]\ : DFN1C0
      port map(D => \Q[3]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[3]_net_1\);
    
    \ARB_BYTE[7]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[7]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[7]_net_1\);
    
    \RECD_SER_WORD_RNO_0[0]\ : MX2
      port map(A => N_17, B => N_19, S => BIT_OS_SEL_1_0, Y => 
        N_33);
    
    \Q[4]\ : DFN1C0
      port map(D => \ADJ_Q[4]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[4]_net_1\);
    
    \ARB_WRD_40M_FIXED[7]\ : DFN1C0
      port map(D => \Q[7]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[7]_net_1\);
    
    \ARB_BYTE_RNIOLA02[1]\ : MX2
      port map(A => N_18, B => N_20, S => BIT_OS_SEL_1_0, Y => 
        N_34);
    
    \ARB_BYTE_RNIBNG52[4]\ : MX2
      port map(A => N_21, B => N_23, S => BIT_OS_SEL_1_0, Y => 
        N_37);
    
    \RECD_SER_WORD_RNO[6]\ : MX2
      port map(A => N_39, B => N_40, S => BIT_OS_SEL_3_0, Y => 
        \N_RECD_SER_WORD[6]\);
    
    \ARB_BYTE[3]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[3]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[3]_net_1\);
    
    \ARB_BYTE_RNI8QGO[3]\ : MX2
      port map(A => \ARB_BYTE[3]_net_1\, B => \ARB_BYTE[7]_net_1\, 
        S => BIT_OS_SEL_0_0, Y => N_20);
    
    \ADJ_Q[5]\ : DFN1C0
      port map(D => \ADJ_Q[3]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[5]_net_1\);
    
    \ARB_BYTE_RNILLMT[6]\ : MX2
      port map(A => \ARB_BYTE[6]_net_1\, B => 
        \ARB_BYTE[10]_net_1\, S => BIT_OS_SEL_0_0, Y => N_23);
    
    \ARB_BYTE[1]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[1]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[1]_net_1\);
    
    \ARB_WRD_40M_FIXED[13]\ : DFN1C0
      port map(D => \Q[13]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[13]_net_1\);
    
    \ARB_BYTE_RNINNMT[11]\ : MX2
      port map(A => \ARB_BYTE[7]_net_1\, B => 
        \ARB_BYTE[11]_net_1\, S => BIT_OS_SEL_0_0, Y => N_24);
    
    \ADJ_Q[0]\ : DFN1C0
      port map(D => \ADJ_SER_IN_R_1DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[0]_net_1\);
    
    \ARB_WRD_40M_FIXED[10]\ : DFN1C0
      port map(D => \Q[10]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[10]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SER320M_3_34_17 is

    port( ELK_TX_DAT                 : in    std_logic_vector(7 downto 0);
          MASTER_SALT_POR_B_i_0_i_14 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_17 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_0  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_8  : in    std_logic;
          ELK_OUT_R                  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_12 : in    std_logic;
          ELK_OUT_F                  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_9  : in    std_logic;
          CCC_160M_FXD               : in    std_logic;
          CLK_40M_GL                 : in    std_logic
        );

end SER320M_3_34_17;

architecture DEF_ARCH of SER320M_3_34_17 is 

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \N_SER_CMD_WORD_R[0]\, \START_RISE\, 
        \N_SER_CMD_WORD_F[0]\, \N_SER_CMD_WORD_R[3]\, 
        \SER_CMD_WORD_R[2]_net_1\, \N_SER_CMD_WORD_R[2]\, 
        \SER_CMD_WORD_R[1]_net_1\, \N_SER_CMD_WORD_R[1]\, 
        \SER_CMD_WORD_R[0]_net_1\, \N_SER_CMD_WORD_F[3]\, 
        \SER_CMD_WORD_F[2]_net_1\, \N_SER_CMD_WORD_F[2]\, 
        \SER_CMD_WORD_F[1]_net_1\, \N_SER_CMD_WORD_F[1]\, 
        \SER_CMD_WORD_F[0]_net_1\, N_START_RISE, 
        \CLK40M_GEN_DEL0\, \SER_OUT_FI\, \SER_OUT_RI\, 
        \SER_CMD_WORD_F[3]_net_1\, \SER_CMD_WORD_R[3]_net_1\, 
        \GND\, \VCC\ : std_logic;

begin 


    SER_OUT_FI : DFN1C0
      port map(D => \SER_CMD_WORD_F[3]_net_1\, CLK => 
        CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_0, Q => 
        \SER_OUT_FI\);
    
    \SER_CMD_WORD_F[3]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[3]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_17, Q => 
        \SER_CMD_WORD_F[3]_net_1\);
    
    \SER_CMD_WORD_R[1]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[1]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_14, Q => 
        \SER_CMD_WORD_R[1]_net_1\);
    
    \SER_CMD_WORD_R[2]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[2]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_14, Q => 
        \SER_CMD_WORD_R[2]_net_1\);
    
    \SER_CMD_WORD_R_RNO[3]\ : MX2
      port map(A => \SER_CMD_WORD_R[2]_net_1\, B => ELK_TX_DAT(7), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_R[3]\);
    
    \SER_CMD_WORD_R_RNO[0]\ : NOR2B
      port map(A => \START_RISE\, B => ELK_TX_DAT(1), Y => 
        \N_SER_CMD_WORD_R[0]\);
    
    \SER_CMD_WORD_F[0]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[0]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_17, Q => 
        \SER_CMD_WORD_F[0]_net_1\);
    
    \SER_CMD_WORD_R_RNO[1]\ : MX2
      port map(A => \SER_CMD_WORD_R[0]_net_1\, B => ELK_TX_DAT(3), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_R[1]\);
    
    \SER_CMD_WORD_F_RNO[2]\ : MX2
      port map(A => \SER_CMD_WORD_F[1]_net_1\, B => ELK_TX_DAT(4), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_F[2]\);
    
    \SER_CMD_WORD_F_RNO[3]\ : MX2
      port map(A => \SER_CMD_WORD_F[2]_net_1\, B => ELK_TX_DAT(6), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_F[3]\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    CLK40M_GEN_DEL0 : DFN1C0
      port map(D => CLK_40M_GL, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_9, Q => \CLK40M_GEN_DEL0\);
    
    SER_OUT_RI : DFN1C0
      port map(D => \SER_CMD_WORD_R[3]_net_1\, CLK => 
        CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_0, Q => 
        \SER_OUT_RI\);
    
    \SER_CMD_WORD_F[2]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[2]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_17, Q => 
        \SER_CMD_WORD_F[2]_net_1\);
    
    \SER_CMD_WORD_F_RNO[1]\ : MX2
      port map(A => \SER_CMD_WORD_F[0]_net_1\, B => ELK_TX_DAT(2), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_F[1]\);
    
    \SER_CMD_WORD_R[0]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[0]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_14, Q => 
        \SER_CMD_WORD_R[0]_net_1\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    START_RISE : DFN1C0
      port map(D => N_START_RISE, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_8, Q => \START_RISE\);
    
    \SER_CMD_WORD_R[3]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[3]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_14, Q => 
        \SER_CMD_WORD_R[3]_net_1\);
    
    \SER_CMD_WORD_F_RNO[0]\ : NOR2B
      port map(A => \START_RISE\, B => ELK_TX_DAT(0), Y => 
        \N_SER_CMD_WORD_F[0]\);
    
    SER_OUT_RDEL : DFN1C0
      port map(D => \SER_OUT_RI\, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_8, Q => ELK_OUT_R);
    
    \SER_CMD_WORD_F[1]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[1]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_17, Q => 
        \SER_CMD_WORD_F[1]_net_1\);
    
    START_RISE_RNO : NOR2B
      port map(A => \CLK40M_GEN_DEL0\, B => CLK_40M_GL, Y => 
        N_START_RISE);
    
    \SER_CMD_WORD_R_RNO[2]\ : MX2
      port map(A => \SER_CMD_WORD_R[1]_net_1\, B => ELK_TX_DAT(5), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_R[2]\);
    
    SER_OUT_FDEL : DFN1C0
      port map(D => \SER_OUT_FI\, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_12, Q => ELK_OUT_F);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity DDR_BIDIR_LVDS_DUAL_CLK_17 is

    port( DCB_SALT_SEL_c_i : in    std_logic;
          ELK17_DAT_P      : inout std_logic := 'Z';
          ELK17_DAT_N      : inout std_logic := 'Z';
          ELK_OUT_R        : in    std_logic;
          ELK_OUT_F        : in    std_logic;
          CCC_160M_FXD     : in    std_logic;
          CCC_160M_ADJ     : in    std_logic;
          ELK_IN_DDR_R     : out   std_logic;
          ELK_IN_DDR_F     : out   std_logic
        );

end DDR_BIDIR_LVDS_DUAL_CLK_17;

architecture DEF_ARCH of DDR_BIDIR_LVDS_DUAL_CLK_17 is 

  component DDR_REG
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          QR  : out   std_logic;
          QF  : out   std_logic
        );
  end component;

  component DDR_OUT
    port( DR  : in    std_logic := 'U';
          DF  : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component BIBUF_LVDS
    port( PADP : inout   std_logic;
          PADN : inout   std_logic;
          D    : in    std_logic := 'U';
          E    : in    std_logic := 'U';
          Y    : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal DDR_BIDIR_LVDS_DUAL_CLK_17_GND, BIBUF_LVDS_0_Y, 
        DDR_OUT_0_Q, \VCC\ : std_logic;

begin 


    DDR_REG_0 : DDR_REG
      port map(D => BIBUF_LVDS_0_Y, CLK => CCC_160M_ADJ, CLR => 
        DDR_BIDIR_LVDS_DUAL_CLK_17_GND, QR => ELK_IN_DDR_R, QF
         => ELK_IN_DDR_F);
    
    DDR_OUT_0 : DDR_OUT
      port map(DR => ELK_OUT_R, DF => ELK_OUT_F, CLK => 
        CCC_160M_FXD, CLR => DDR_BIDIR_LVDS_DUAL_CLK_17_GND, Q
         => DDR_OUT_0_Q);
    
    BIBUF_LVDS_0 : BIBUF_LVDS
      port map(PADP => ELK17_DAT_P, PADN => ELK17_DAT_N, D => 
        DDR_OUT_0_Q, E => DCB_SALT_SEL_c_i, Y => BIBUF_LVDS_0_Y);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    GND_i : GND
      port map(Y => DDR_BIDIR_LVDS_DUAL_CLK_17_GND);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SYNC_DAT_SEL_17 is

    port( ELK_TX_DAT                 : out   std_logic_vector(7 downto 0);
          PATT_ELK_DAT_17            : in    std_logic_vector(7 downto 0);
          OP_MODE_c_6_0              : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_12 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_11 : in    std_logic;
          CLK_40M_GL                 : in    std_logic
        );

end SYNC_DAT_SEL_17;

architecture DEF_ARCH of SYNC_DAT_SEL_17 is 

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \N_SERDAT[0]\, \N_SERDAT[1]\, \N_SERDAT[2]\, 
        \N_SERDAT[3]\, \N_SERDAT[4]\, \N_SERDAT[5]\, 
        \N_SERDAT[6]\, \N_SERDAT[7]\, \GND\, \VCC\ : std_logic;

begin 


    \SERDAT_RNO[4]\ : NOR2A
      port map(A => PATT_ELK_DAT_17(4), B => OP_MODE_c_6_0, Y => 
        \N_SERDAT[4]\);
    
    \SERDAT_RNO[0]\ : NOR2A
      port map(A => PATT_ELK_DAT_17(0), B => OP_MODE_c_6_0, Y => 
        \N_SERDAT[0]\);
    
    \SERDAT[6]\ : DFN1C0
      port map(D => \N_SERDAT[6]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_11, Q => ELK_TX_DAT(6));
    
    \SERDAT[4]\ : DFN1C0
      port map(D => \N_SERDAT[4]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_11, Q => ELK_TX_DAT(4));
    
    \SERDAT_RNO[7]\ : OR2
      port map(A => PATT_ELK_DAT_17(7), B => OP_MODE_c_6_0, Y => 
        \N_SERDAT[7]\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \SERDAT_RNO[3]\ : OR2
      port map(A => PATT_ELK_DAT_17(3), B => OP_MODE_c_6_0, Y => 
        \N_SERDAT[3]\);
    
    \SERDAT_RNO[2]\ : OR2
      port map(A => PATT_ELK_DAT_17(2), B => OP_MODE_c_6_0, Y => 
        \N_SERDAT[2]\);
    
    \SERDAT[5]\ : DFN1C0
      port map(D => \N_SERDAT[5]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_11, Q => ELK_TX_DAT(5));
    
    \SERDAT[7]\ : DFN1C0
      port map(D => \N_SERDAT[7]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_12, Q => ELK_TX_DAT(7));
    
    GND_i : GND
      port map(Y => \GND\);
    
    \SERDAT_RNO[5]\ : NOR2A
      port map(A => PATT_ELK_DAT_17(5), B => OP_MODE_c_6_0, Y => 
        \N_SERDAT[5]\);
    
    \SERDAT[0]\ : DFN1C0
      port map(D => \N_SERDAT[0]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_11, Q => ELK_TX_DAT(0));
    
    \SERDAT_RNO[6]\ : NOR2A
      port map(A => PATT_ELK_DAT_17(6), B => OP_MODE_c_6_0, Y => 
        \N_SERDAT[6]\);
    
    \SERDAT[1]\ : DFN1C0
      port map(D => \N_SERDAT[1]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_11, Q => ELK_TX_DAT(1));
    
    \SERDAT_RNO[1]\ : OR2
      port map(A => PATT_ELK_DAT_17(1), B => OP_MODE_c_6_0, Y => 
        \N_SERDAT[1]\);
    
    \SERDAT[3]\ : DFN1C0
      port map(D => \N_SERDAT[3]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_11, Q => ELK_TX_DAT(3));
    
    \SERDAT[2]\ : DFN1C0
      port map(D => \N_SERDAT[2]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_11, Q => ELK_TX_DAT(2));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity ELINK_SLAVE_15_12 is

    port( BIT_OS_SEL_0_0             : in    std_logic;
          BIT_OS_SEL_1_0             : in    std_logic;
          BIT_OS_SEL_2               : in    std_logic_vector(2 downto 0);
          BIT_OS_SEL_3_0             : in    std_logic;
          ELK_RX_SER_WORD_17         : out   std_logic_vector(7 downto 0);
          OP_MODE_c_6_0              : in    std_logic;
          PATT_ELK_DAT_17            : in    std_logic_vector(7 downto 0);
          MASTER_DCB_POR_B_i_0_i     : in    std_logic;
          ELK17_DAT_N                : inout std_logic := 'Z';
          ELK17_DAT_P                : inout std_logic := 'Z';
          DCB_SALT_SEL_c_i           : in    std_logic;
          CCC_160M_FXD               : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_9  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_8  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_0  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_17 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_14 : in    std_logic;
          CLK_40M_GL                 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_11 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_12 : in    std_logic;
          DEV_RST_B_c_1              : in    std_logic;
          CCC_160M_ADJ               : in    std_logic
        );

end ELINK_SLAVE_15_12;

architecture DEF_ARCH of ELINK_SLAVE_15_12 is 

  component SLAVE_DES320S_1_17_15
    port( ELK_RX_SER_WORD_17     : out   std_logic_vector(7 downto 0);
          BIT_OS_SEL_3_0         : in    std_logic := 'U';
          BIT_OS_SEL_2           : in    std_logic_vector(2 downto 0) := (others => 'U');
          BIT_OS_SEL_1_0         : in    std_logic := 'U';
          BIT_OS_SEL_0_0         : in    std_logic := 'U';
          CLK_40M_GL             : in    std_logic := 'U';
          CCC_160M_FXD           : in    std_logic := 'U';
          ELK_IN_R               : in    std_logic := 'U';
          ELK_IN_F               : in    std_logic := 'U';
          MASTER_DCB_POR_B_i_0_i : in    std_logic := 'U';
          CCC_160M_ADJ           : in    std_logic := 'U'
        );
  end component;

  component SER320M_3_34_17
    port( ELK_TX_DAT                 : in    std_logic_vector(7 downto 0) := (others => 'U');
          MASTER_SALT_POR_B_i_0_i_14 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_17 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_0  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_8  : in    std_logic := 'U';
          ELK_OUT_R                  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_12 : in    std_logic := 'U';
          ELK_OUT_F                  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_9  : in    std_logic := 'U';
          CCC_160M_FXD               : in    std_logic := 'U';
          CLK_40M_GL                 : in    std_logic := 'U'
        );
  end component;

  component DDR_BIDIR_LVDS_DUAL_CLK_17
    port( DCB_SALT_SEL_c_i : in    std_logic := 'U';
          ELK17_DAT_P      : inout   std_logic;
          ELK17_DAT_N      : inout   std_logic;
          ELK_OUT_R        : in    std_logic := 'U';
          ELK_OUT_F        : in    std_logic := 'U';
          CCC_160M_FXD     : in    std_logic := 'U';
          CCC_160M_ADJ     : in    std_logic := 'U';
          ELK_IN_DDR_R     : out   std_logic;
          ELK_IN_DDR_F     : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component SYNC_DAT_SEL_17
    port( ELK_TX_DAT                 : out   std_logic_vector(7 downto 0);
          PATT_ELK_DAT_17            : in    std_logic_vector(7 downto 0) := (others => 'U');
          OP_MODE_c_6_0              : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_12 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_11 : in    std_logic := 'U';
          CLK_40M_GL                 : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \ELK_IN_F\, ELK_IN_DDR_F, \ELK_IN_R\, ELK_IN_DDR_R, 
        \ELK_TX_DAT[0]\, \ELK_TX_DAT[1]\, \ELK_TX_DAT[2]\, 
        \ELK_TX_DAT[3]\, \ELK_TX_DAT[4]\, \ELK_TX_DAT[5]\, 
        \ELK_TX_DAT[6]\, \ELK_TX_DAT[7]\, ELK_OUT_R, ELK_OUT_F, 
        \GND\, \VCC\ : std_logic;

    for all : SLAVE_DES320S_1_17_15
	Use entity work.SLAVE_DES320S_1_17_15(DEF_ARCH);
    for all : SER320M_3_34_17
	Use entity work.SER320M_3_34_17(DEF_ARCH);
    for all : DDR_BIDIR_LVDS_DUAL_CLK_17
	Use entity work.DDR_BIDIR_LVDS_DUAL_CLK_17(DEF_ARCH);
    for all : SYNC_DAT_SEL_17
	Use entity work.SYNC_DAT_SEL_17(DEF_ARCH);
begin 


    U_SLAVE_1ELK : SLAVE_DES320S_1_17_15
      port map(ELK_RX_SER_WORD_17(7) => ELK_RX_SER_WORD_17(7), 
        ELK_RX_SER_WORD_17(6) => ELK_RX_SER_WORD_17(6), 
        ELK_RX_SER_WORD_17(5) => ELK_RX_SER_WORD_17(5), 
        ELK_RX_SER_WORD_17(4) => ELK_RX_SER_WORD_17(4), 
        ELK_RX_SER_WORD_17(3) => ELK_RX_SER_WORD_17(3), 
        ELK_RX_SER_WORD_17(2) => ELK_RX_SER_WORD_17(2), 
        ELK_RX_SER_WORD_17(1) => ELK_RX_SER_WORD_17(1), 
        ELK_RX_SER_WORD_17(0) => ELK_RX_SER_WORD_17(0), 
        BIT_OS_SEL_3_0 => BIT_OS_SEL_3_0, BIT_OS_SEL_2(2) => 
        BIT_OS_SEL_2(2), BIT_OS_SEL_2(1) => BIT_OS_SEL_2(1), 
        BIT_OS_SEL_2(0) => BIT_OS_SEL_2(0), BIT_OS_SEL_1_0 => 
        BIT_OS_SEL_1_0, BIT_OS_SEL_0_0 => BIT_OS_SEL_0_0, 
        CLK_40M_GL => CLK_40M_GL, CCC_160M_FXD => CCC_160M_FXD, 
        ELK_IN_R => \ELK_IN_R\, ELK_IN_F => \ELK_IN_F\, 
        MASTER_DCB_POR_B_i_0_i => MASTER_DCB_POR_B_i_0_i, 
        CCC_160M_ADJ => CCC_160M_ADJ);
    
    U_ELK1_CMD_TX : SER320M_3_34_17
      port map(ELK_TX_DAT(7) => \ELK_TX_DAT[7]\, ELK_TX_DAT(6)
         => \ELK_TX_DAT[6]\, ELK_TX_DAT(5) => \ELK_TX_DAT[5]\, 
        ELK_TX_DAT(4) => \ELK_TX_DAT[4]\, ELK_TX_DAT(3) => 
        \ELK_TX_DAT[3]\, ELK_TX_DAT(2) => \ELK_TX_DAT[2]\, 
        ELK_TX_DAT(1) => \ELK_TX_DAT[1]\, ELK_TX_DAT(0) => 
        \ELK_TX_DAT[0]\, MASTER_SALT_POR_B_i_0_i_14 => 
        MASTER_SALT_POR_B_i_0_i_14, MASTER_SALT_POR_B_i_0_i_17
         => MASTER_SALT_POR_B_i_0_i_17, MASTER_SALT_POR_B_i_0_i_0
         => MASTER_SALT_POR_B_i_0_i_0, MASTER_SALT_POR_B_i_0_i_8
         => MASTER_SALT_POR_B_i_0_i_8, ELK_OUT_R => ELK_OUT_R, 
        MASTER_SALT_POR_B_i_0_i_12 => MASTER_SALT_POR_B_i_0_i_12, 
        ELK_OUT_F => ELK_OUT_F, MASTER_SALT_POR_B_i_0_i_9 => 
        MASTER_SALT_POR_B_i_0_i_9, CCC_160M_FXD => CCC_160M_FXD, 
        CLK_40M_GL => CLK_40M_GL);
    
    U_DDR_ELK1 : DDR_BIDIR_LVDS_DUAL_CLK_17
      port map(DCB_SALT_SEL_c_i => DCB_SALT_SEL_c_i, ELK17_DAT_P
         => ELK17_DAT_P, ELK17_DAT_N => ELK17_DAT_N, ELK_OUT_R
         => ELK_OUT_R, ELK_OUT_F => ELK_OUT_F, CCC_160M_FXD => 
        CCC_160M_FXD, CCC_160M_ADJ => CCC_160M_ADJ, ELK_IN_DDR_R
         => ELK_IN_DDR_R, ELK_IN_DDR_F => ELK_IN_DDR_F);
    
    ELK_IN_F : DFN1C0
      port map(D => ELK_IN_DDR_F, CLK => CCC_160M_ADJ, CLR => 
        DEV_RST_B_c_1, Q => \ELK_IN_F\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    U_ELK1_SERDAT_SOURCE : SYNC_DAT_SEL_17
      port map(ELK_TX_DAT(7) => \ELK_TX_DAT[7]\, ELK_TX_DAT(6)
         => \ELK_TX_DAT[6]\, ELK_TX_DAT(5) => \ELK_TX_DAT[5]\, 
        ELK_TX_DAT(4) => \ELK_TX_DAT[4]\, ELK_TX_DAT(3) => 
        \ELK_TX_DAT[3]\, ELK_TX_DAT(2) => \ELK_TX_DAT[2]\, 
        ELK_TX_DAT(1) => \ELK_TX_DAT[1]\, ELK_TX_DAT(0) => 
        \ELK_TX_DAT[0]\, PATT_ELK_DAT_17(7) => PATT_ELK_DAT_17(7), 
        PATT_ELK_DAT_17(6) => PATT_ELK_DAT_17(6), 
        PATT_ELK_DAT_17(5) => PATT_ELK_DAT_17(5), 
        PATT_ELK_DAT_17(4) => PATT_ELK_DAT_17(4), 
        PATT_ELK_DAT_17(3) => PATT_ELK_DAT_17(3), 
        PATT_ELK_DAT_17(2) => PATT_ELK_DAT_17(2), 
        PATT_ELK_DAT_17(1) => PATT_ELK_DAT_17(1), 
        PATT_ELK_DAT_17(0) => PATT_ELK_DAT_17(0), OP_MODE_c_6_0
         => OP_MODE_c_6_0, MASTER_SALT_POR_B_i_0_i_12 => 
        MASTER_SALT_POR_B_i_0_i_12, MASTER_SALT_POR_B_i_0_i_11
         => MASTER_SALT_POR_B_i_0_i_11, CLK_40M_GL => CLK_40M_GL);
    
    ELK_IN_R : DFN1C0
      port map(D => ELK_IN_DDR_R, CLK => CCC_160M_ADJ, CLR => 
        DEV_RST_B_c_1, Q => \ELK_IN_R\);
    
    GND_i : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SLAVE_DES320S_1_17_13 is

    port( ELK_RX_SER_WORD_15     : out   std_logic_vector(7 downto 0);
          BIT_OS_SEL_3           : in    std_logic_vector(1 downto 0);
          BIT_OS_SEL_4_0         : in    std_logic;
          BIT_OS_SEL_2           : in    std_logic_vector(2 downto 1);
          BIT_OS_SEL_1_0         : in    std_logic;
          CLK_40M_GL             : in    std_logic;
          CCC_160M_FXD           : in    std_logic;
          ELK_IN_R               : in    std_logic;
          ELK_IN_F               : in    std_logic;
          MASTER_DCB_POR_B_i_0_i : in    std_logic;
          CCC_160M_ADJ           : in    std_logic
        );

end SLAVE_DES320S_1_17_13;

architecture DEF_ARCH of SLAVE_DES320S_1_17_13 is 

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal N_17, \ARB_BYTE[0]_net_1\, \ARB_BYTE[4]_net_1\, N_18, 
        \ARB_BYTE[1]_net_1\, \ARB_BYTE[5]_net_1\, N_19, 
        \ARB_BYTE[2]_net_1\, \ARB_BYTE[6]_net_1\, N_20, 
        \ARB_BYTE[3]_net_1\, \ARB_BYTE[7]_net_1\, N_21, 
        \ARB_BYTE[8]_net_1\, N_22, \ARB_BYTE[9]_net_1\, N_23, 
        \ARB_BYTE[10]_net_1\, N_24, \ARB_BYTE[11]_net_1\, N_31, 
        \ARB_BYTE[12]_net_1\, N_32, \ARB_BYTE[13]_net_1\, N_33, 
        N_34, N_35, N_36, N_37, N_38, N_39, N_40, N_56, 
        \ARB_BYTE[14]_net_1\, N_64, \N_RECD_SER_WORD[0]\, 
        \N_RECD_SER_WORD[1]\, \N_RECD_SER_WORD[2]\, 
        \N_RECD_SER_WORD[3]\, \N_RECD_SER_WORD[4]\, 
        \N_RECD_SER_WORD[5]\, \N_RECD_SER_WORD[6]\, 
        \N_RECD_SER_WORD[7]\, \ADJ_SER_IN_F_0DEL\, 
        \ADJ_SER_IN_R_0DEL\, \ADJ_SER_IN_F_1DEL\, 
        \ADJ_SER_IN_R_1DEL\, \Q[0]_net_1\, \ADJ_Q[0]_net_1\, 
        \Q[1]_net_1\, \ADJ_Q[1]_net_1\, \Q[2]_net_1\, 
        \ADJ_Q[2]_net_1\, \Q[3]_net_1\, \ADJ_Q[3]_net_1\, 
        \Q[4]_net_1\, \ADJ_Q[4]_net_1\, \Q[5]_net_1\, 
        \ADJ_Q[5]_net_1\, \Q[6]_net_1\, \ADJ_Q[6]_net_1\, 
        \Q[7]_net_1\, \ADJ_Q[7]_net_1\, \Q[8]_net_1\, 
        \ADJ_Q[8]_net_1\, \Q[9]_net_1\, \ADJ_Q[9]_net_1\, 
        \Q[10]_net_1\, \ADJ_Q[10]_net_1\, \Q[11]_net_1\, 
        \ADJ_Q[11]_net_1\, \Q[12]_net_1\, \ADJ_Q[12]_net_1\, 
        \Q[13]_net_1\, \ADJ_Q[13]_net_1\, \Q[14]_net_1\, 
        \ADJ_Q[14]_net_1\, \ARB_WRD_40M_FIXED[0]_net_1\, 
        \ARB_WRD_40M_FIXED[1]_net_1\, 
        \ARB_WRD_40M_FIXED[2]_net_1\, 
        \ARB_WRD_40M_FIXED[3]_net_1\, 
        \ARB_WRD_40M_FIXED[4]_net_1\, 
        \ARB_WRD_40M_FIXED[5]_net_1\, 
        \ARB_WRD_40M_FIXED[6]_net_1\, 
        \ARB_WRD_40M_FIXED[7]_net_1\, 
        \ARB_WRD_40M_FIXED[8]_net_1\, 
        \ARB_WRD_40M_FIXED[9]_net_1\, 
        \ARB_WRD_40M_FIXED[10]_net_1\, 
        \ARB_WRD_40M_FIXED[11]_net_1\, 
        \ARB_WRD_40M_FIXED[12]_net_1\, 
        \ARB_WRD_40M_FIXED[13]_net_1\, 
        \ARB_WRD_40M_FIXED[14]_net_1\, \GND\, \VCC\ : std_logic;

begin 


    \RECD_SER_WORD_RNO[5]\ : MX2
      port map(A => N_38, B => N_39, S => BIT_OS_SEL_3(0), Y => 
        \N_RECD_SER_WORD[5]\);
    
    \ARB_WRD_40M_FIXED[9]\ : DFN1C0
      port map(D => \Q[9]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[9]_net_1\);
    
    \ADJ_Q[4]\ : DFN1C0
      port map(D => \ADJ_Q[2]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[4]_net_1\);
    
    \ARB_BYTE_RNI198Q[1]\ : MX2
      port map(A => \ARB_BYTE[1]_net_1\, B => \ARB_BYTE[5]_net_1\, 
        S => BIT_OS_SEL_1_0, Y => N_18);
    
    \ARB_BYTE[6]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[6]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[6]_net_1\);
    
    ADJ_SER_IN_F_1DEL : DFN1C0
      port map(D => \ADJ_SER_IN_F_0DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_F_1DEL\);
    
    \ARB_BYTE[0]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[0]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[0]_net_1\);
    
    \Q[11]\ : DFN1C0
      port map(D => \ADJ_Q[11]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[11]_net_1\);
    
    \ADJ_Q[8]\ : DFN1C0
      port map(D => \ADJ_Q[6]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[8]_net_1\);
    
    \ADJ_Q[6]\ : DFN1C0
      port map(D => \ADJ_Q[4]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[6]_net_1\);
    
    \ADJ_Q[12]\ : DFN1C0
      port map(D => \ADJ_Q[10]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[12]_net_1\);
    
    \RECD_SER_WORD_RNO_1[0]\ : MX2
      port map(A => \ARB_BYTE[0]_net_1\, B => \ARB_BYTE[4]_net_1\, 
        S => BIT_OS_SEL_1_0, Y => N_17);
    
    \Q[1]\ : DFN1C0
      port map(D => \ADJ_Q[1]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[1]_net_1\);
    
    \ARB_BYTE_RNIJUSK1[1]\ : MX2
      port map(A => N_18, B => N_20, S => BIT_OS_SEL_2(1), Y => 
        N_34);
    
    \ARB_BYTE_RNIQ0S41[13]\ : MX2
      port map(A => N_24, B => N_32, S => BIT_OS_SEL_2(1), Y => 
        N_40);
    
    \ARB_BYTE_RNIA2BK1[11]\ : MX2
      port map(A => N_22, B => N_24, S => BIT_OS_SEL_2(1), Y => 
        N_38);
    
    \ARB_BYTE[4]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[4]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[4]_net_1\);
    
    \ADJ_Q[2]\ : DFN1C0
      port map(D => \ADJ_Q[0]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[2]_net_1\);
    
    \RECD_SER_WORD_RNO_1[7]\ : MX2
      port map(A => \ARB_BYTE[10]_net_1\, B => 
        \ARB_BYTE[14]_net_1\, S => BIT_OS_SEL_4_0, Y => N_56);
    
    \RECD_SER_WORD[4]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[4]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_15(4));
    
    \Q[5]\ : DFN1C0
      port map(D => \ADJ_Q[5]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[5]_net_1\);
    
    \ADJ_Q[11]\ : DFN1C0
      port map(D => \ADJ_Q[9]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[11]_net_1\);
    
    \ARB_BYTE_RNI5D8Q[3]\ : MX2
      port map(A => \ARB_BYTE[3]_net_1\, B => \ARB_BYTE[7]_net_1\, 
        S => BIT_OS_SEL_1_0, Y => N_20);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \ADJ_Q[3]\ : DFN1C0
      port map(D => \ADJ_Q[1]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[3]_net_1\);
    
    \Q[10]\ : DFN1C0
      port map(D => \ADJ_Q[10]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[10]_net_1\);
    
    \ARB_WRD_40M_FIXED[6]\ : DFN1C0
      port map(D => \Q[6]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[6]_net_1\);
    
    \ARB_BYTE_RNII6MP[10]\ : MX2
      port map(A => \ARB_BYTE[6]_net_1\, B => 
        \ARB_BYTE[10]_net_1\, S => BIT_OS_SEL_1_0, Y => N_23);
    
    \ARB_WRD_40M_FIXED[1]\ : DFN1C0
      port map(D => \Q[1]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[1]_net_1\);
    
    \RECD_SER_WORD[3]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[3]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_15(3));
    
    \RECD_SER_WORD[0]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[0]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_15(0));
    
    \RECD_SER_WORD_RNO[3]\ : MX2
      port map(A => N_36, B => N_37, S => BIT_OS_SEL_3(0), Y => 
        \N_RECD_SER_WORD[3]\);
    
    \Q[0]\ : DFN1C0
      port map(D => \ADJ_Q[0]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[0]_net_1\);
    
    \RECD_SER_WORD_RNO_0[7]\ : MX2
      port map(A => N_31, B => N_56, S => BIT_OS_SEL_3(1), Y => 
        N_64);
    
    \Q[7]\ : DFN1C0
      port map(D => \ADJ_Q[7]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[7]_net_1\);
    
    \ARB_BYTE[14]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[14]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[14]_net_1\);
    
    \ARB_WRD_40M_FIXED[2]\ : DFN1C0
      port map(D => \Q[2]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[2]_net_1\);
    
    \ARB_WRD_40M_FIXED[14]\ : DFN1C0
      port map(D => \Q[14]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[14]_net_1\);
    
    \RECD_SER_WORD_RNO[2]\ : MX2
      port map(A => N_35, B => N_36, S => BIT_OS_SEL_3(0), Y => 
        \N_RECD_SER_WORD[2]\);
    
    \ARB_BYTE[2]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[2]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[2]_net_1\);
    
    \ADJ_Q[7]\ : DFN1C0
      port map(D => \ADJ_Q[5]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[7]_net_1\);
    
    \ARB_BYTE_RNIK8MP[11]\ : MX2
      port map(A => \ARB_BYTE[7]_net_1\, B => 
        \ARB_BYTE[11]_net_1\, S => BIT_OS_SEL_1_0, Y => N_24);
    
    \ARB_BYTE[8]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[8]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[8]_net_1\);
    
    \RECD_SER_WORD[5]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[5]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_15(5));
    
    \ARB_BYTE[12]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[12]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[12]_net_1\);
    
    \RECD_SER_WORD[1]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[1]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_15(1));
    
    \ARB_BYTE_RNI6UAK1[10]\ : MX2
      port map(A => N_21, B => N_23, S => BIT_OS_SEL_2(1), Y => 
        N_37);
    
    \Q[3]\ : DFN1C0
      port map(D => \ADJ_Q[3]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[3]_net_1\);
    
    \ARB_BYTE_RNINDPA[12]\ : MX2
      port map(A => \ARB_BYTE[8]_net_1\, B => 
        \ARB_BYTE[12]_net_1\, S => BIT_OS_SEL_2(2), Y => N_31);
    
    ADJ_SER_IN_F_0DEL : DFN1C0
      port map(D => ELK_IN_F, CLK => CCC_160M_ADJ, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_F_0DEL\);
    
    \RECD_SER_WORD_RNO[7]\ : MX2
      port map(A => N_40, B => N_64, S => BIT_OS_SEL_3(0), Y => 
        \N_RECD_SER_WORD[7]\);
    
    \RECD_SER_WORD_RNO[1]\ : MX2
      port map(A => N_34, B => N_35, S => BIT_OS_SEL_3(0), Y => 
        \N_RECD_SER_WORD[1]\);
    
    \ARB_WRD_40M_FIXED[4]\ : DFN1C0
      port map(D => \Q[4]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[4]_net_1\);
    
    \RECD_SER_WORD_RNO[0]\ : MX2
      port map(A => N_33, B => N_34, S => BIT_OS_SEL_3(0), Y => 
        \N_RECD_SER_WORD[0]\);
    
    \Q[6]\ : DFN1C0
      port map(D => \ADJ_Q[6]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[6]_net_1\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \ARB_WRD_40M_FIXED[8]\ : DFN1C0
      port map(D => \Q[8]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[8]_net_1\);
    
    \ARB_BYTE_RNI7F8Q[4]\ : MX2
      port map(A => \ARB_BYTE[4]_net_1\, B => \ARB_BYTE[8]_net_1\, 
        S => BIT_OS_SEL_1_0, Y => N_21);
    
    \ARB_BYTE[11]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[11]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[11]_net_1\);
    
    \Q[9]\ : DFN1C0
      port map(D => \ADJ_Q[9]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[9]_net_1\);
    
    \Q[14]\ : DFN1C0
      port map(D => \ADJ_Q[14]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[14]_net_1\);
    
    ADJ_SER_IN_R_0DEL : DFN1C0
      port map(D => ELK_IN_R, CLK => CCC_160M_ADJ, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_R_0DEL\);
    
    \Q[13]\ : DFN1C0
      port map(D => \ADJ_Q[13]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[13]_net_1\);
    
    \ARB_BYTE[9]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[9]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[9]_net_1\);
    
    ADJ_SER_IN_R_1DEL : DFN1C0
      port map(D => \ADJ_SER_IN_R_0DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_R_1DEL\);
    
    \ARB_BYTE[10]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[10]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[10]_net_1\);
    
    \ADJ_Q[9]\ : DFN1C0
      port map(D => \ADJ_Q[7]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[9]_net_1\);
    
    \RECD_SER_WORD[7]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[7]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_15(7));
    
    \ARB_WRD_40M_FIXED[5]\ : DFN1C0
      port map(D => \Q[5]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[5]_net_1\);
    
    \ARB_WRD_40M_FIXED[12]\ : DFN1C0
      port map(D => \Q[12]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[12]_net_1\);
    
    \ARB_BYTE_RNIMSR41[10]\ : MX2
      port map(A => N_23, B => N_31, S => BIT_OS_SEL_2(1), Y => 
        N_39);
    
    \ARB_WRD_40M_FIXED[11]\ : DFN1C0
      port map(D => \Q[11]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[11]_net_1\);
    
    \ARB_WRD_40M_FIXED[0]\ : DFN1C0
      port map(D => \Q[0]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[0]_net_1\);
    
    \ADJ_Q[10]\ : DFN1C0
      port map(D => \ADJ_Q[8]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[10]_net_1\);
    
    \Q[2]\ : DFN1C0
      port map(D => \ADJ_Q[2]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[2]_net_1\);
    
    \ARB_BYTE_RNIPFPA[13]\ : MX2
      port map(A => \ARB_BYTE[9]_net_1\, B => 
        \ARB_BYTE[13]_net_1\, S => BIT_OS_SEL_2(2), Y => N_32);
    
    \ARB_BYTE_RNI9H8Q[5]\ : MX2
      port map(A => \ARB_BYTE[5]_net_1\, B => \ARB_BYTE[9]_net_1\, 
        S => BIT_OS_SEL_1_0, Y => N_22);
    
    \ADJ_Q[1]\ : DFN1C0
      port map(D => \ADJ_SER_IN_F_1DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[1]_net_1\);
    
    \RECD_SER_WORD[6]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[6]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_15(6));
    
    \ARB_BYTE_RNI3B8Q[2]\ : MX2
      port map(A => \ARB_BYTE[2]_net_1\, B => \ARB_BYTE[6]_net_1\, 
        S => BIT_OS_SEL_1_0, Y => N_19);
    
    \RECD_SER_WORD[2]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[2]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_15(2));
    
    \ADJ_Q[13]\ : DFN1C0
      port map(D => \ADJ_Q[11]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[13]_net_1\);
    
    \ARB_BYTE_RNIR6TK1[3]\ : MX2
      port map(A => N_20, B => N_22, S => BIT_OS_SEL_2(1), Y => 
        N_36);
    
    \Q[8]\ : DFN1C0
      port map(D => \ADJ_Q[8]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[8]_net_1\);
    
    \ARB_BYTE[5]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[5]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[5]_net_1\);
    
    \ADJ_Q[14]\ : DFN1C0
      port map(D => \ADJ_Q[12]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[14]_net_1\);
    
    \RECD_SER_WORD_RNO[4]\ : MX2
      port map(A => N_37, B => N_38, S => BIT_OS_SEL_3(0), Y => 
        \N_RECD_SER_WORD[4]\);
    
    \Q[12]\ : DFN1C0
      port map(D => \ADJ_Q[12]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[12]_net_1\);
    
    \ARB_BYTE[13]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[13]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[13]_net_1\);
    
    \ARB_WRD_40M_FIXED[3]\ : DFN1C0
      port map(D => \Q[3]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[3]_net_1\);
    
    \ARB_BYTE[7]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[7]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[7]_net_1\);
    
    \RECD_SER_WORD_RNO_0[0]\ : MX2
      port map(A => N_17, B => N_19, S => BIT_OS_SEL_2(1), Y => 
        N_33);
    
    \Q[4]\ : DFN1C0
      port map(D => \ADJ_Q[4]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[4]_net_1\);
    
    \ARB_WRD_40M_FIXED[7]\ : DFN1C0
      port map(D => \Q[7]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[7]_net_1\);
    
    \RECD_SER_WORD_RNO[6]\ : MX2
      port map(A => N_39, B => N_40, S => BIT_OS_SEL_3(0), Y => 
        \N_RECD_SER_WORD[6]\);
    
    \ARB_BYTE[3]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[3]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[3]_net_1\);
    
    \ADJ_Q[5]\ : DFN1C0
      port map(D => \ADJ_Q[3]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[5]_net_1\);
    
    \ARB_BYTE[1]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[1]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[1]_net_1\);
    
    \ARB_BYTE_RNIN2TK1[2]\ : MX2
      port map(A => N_19, B => N_21, S => BIT_OS_SEL_2(1), Y => 
        N_35);
    
    \ARB_WRD_40M_FIXED[13]\ : DFN1C0
      port map(D => \Q[13]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[13]_net_1\);
    
    \ADJ_Q[0]\ : DFN1C0
      port map(D => \ADJ_SER_IN_R_1DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[0]_net_1\);
    
    \ARB_WRD_40M_FIXED[10]\ : DFN1C0
      port map(D => \Q[10]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[10]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SER320M_3_34_15 is

    port( ELK_TX_DAT                : in    std_logic_vector(7 downto 0);
          MASTER_SALT_POR_B_i_0_i_6 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_1 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_9 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_5 : in    std_logic;
          ELK_OUT_R                 : out   std_logic;
          ELK_OUT_F                 : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_8 : in    std_logic;
          CCC_160M_FXD              : in    std_logic;
          CLK_40M_GL                : in    std_logic
        );

end SER320M_3_34_15;

architecture DEF_ARCH of SER320M_3_34_15 is 

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \N_SER_CMD_WORD_R[0]\, \START_RISE\, 
        \N_SER_CMD_WORD_F[0]\, \N_SER_CMD_WORD_R[3]\, 
        \SER_CMD_WORD_R[2]_net_1\, \N_SER_CMD_WORD_R[2]\, 
        \SER_CMD_WORD_R[1]_net_1\, \N_SER_CMD_WORD_R[1]\, 
        \SER_CMD_WORD_R[0]_net_1\, \N_SER_CMD_WORD_F[3]\, 
        \SER_CMD_WORD_F[2]_net_1\, \N_SER_CMD_WORD_F[2]\, 
        \SER_CMD_WORD_F[1]_net_1\, \N_SER_CMD_WORD_F[1]\, 
        \SER_CMD_WORD_F[0]_net_1\, N_START_RISE, 
        \CLK40M_GEN_DEL0\, \SER_OUT_FI\, \SER_OUT_RI\, 
        \SER_CMD_WORD_F[3]_net_1\, \SER_CMD_WORD_R[3]_net_1\, 
        \GND\, \VCC\ : std_logic;

begin 


    SER_OUT_FI : DFN1C0
      port map(D => \SER_CMD_WORD_F[3]_net_1\, CLK => 
        CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_1, Q => 
        \SER_OUT_FI\);
    
    \SER_CMD_WORD_F[3]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[3]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_9, Q => 
        \SER_CMD_WORD_F[3]_net_1\);
    
    \SER_CMD_WORD_R[1]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[1]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_6, Q => 
        \SER_CMD_WORD_R[1]_net_1\);
    
    \SER_CMD_WORD_R[2]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[2]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_6, Q => 
        \SER_CMD_WORD_R[2]_net_1\);
    
    \SER_CMD_WORD_R_RNO[3]\ : MX2
      port map(A => \SER_CMD_WORD_R[2]_net_1\, B => ELK_TX_DAT(7), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_R[3]\);
    
    \SER_CMD_WORD_R_RNO[0]\ : NOR2B
      port map(A => \START_RISE\, B => ELK_TX_DAT(1), Y => 
        \N_SER_CMD_WORD_R[0]\);
    
    \SER_CMD_WORD_F[0]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[0]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_9, Q => 
        \SER_CMD_WORD_F[0]_net_1\);
    
    \SER_CMD_WORD_R_RNO[1]\ : MX2
      port map(A => \SER_CMD_WORD_R[0]_net_1\, B => ELK_TX_DAT(3), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_R[1]\);
    
    \SER_CMD_WORD_F_RNO[2]\ : MX2
      port map(A => \SER_CMD_WORD_F[1]_net_1\, B => ELK_TX_DAT(4), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_F[2]\);
    
    \SER_CMD_WORD_F_RNO[3]\ : MX2
      port map(A => \SER_CMD_WORD_F[2]_net_1\, B => ELK_TX_DAT(6), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_F[3]\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    CLK40M_GEN_DEL0 : DFN1C0
      port map(D => CLK_40M_GL, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_8, Q => \CLK40M_GEN_DEL0\);
    
    SER_OUT_RI : DFN1C0
      port map(D => \SER_CMD_WORD_R[3]_net_1\, CLK => 
        CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_1, Q => 
        \SER_OUT_RI\);
    
    \SER_CMD_WORD_F[2]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[2]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_9, Q => 
        \SER_CMD_WORD_F[2]_net_1\);
    
    \SER_CMD_WORD_F_RNO[1]\ : MX2
      port map(A => \SER_CMD_WORD_F[0]_net_1\, B => ELK_TX_DAT(2), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_F[1]\);
    
    \SER_CMD_WORD_R[0]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[0]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_6, Q => 
        \SER_CMD_WORD_R[0]_net_1\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    START_RISE : DFN1C0
      port map(D => N_START_RISE, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_9, Q => \START_RISE\);
    
    \SER_CMD_WORD_R[3]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[3]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_6, Q => 
        \SER_CMD_WORD_R[3]_net_1\);
    
    \SER_CMD_WORD_F_RNO[0]\ : NOR2B
      port map(A => \START_RISE\, B => ELK_TX_DAT(0), Y => 
        \N_SER_CMD_WORD_F[0]\);
    
    SER_OUT_RDEL : DFN1C0
      port map(D => \SER_OUT_RI\, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_5, Q => ELK_OUT_R);
    
    \SER_CMD_WORD_F[1]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[1]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_9, Q => 
        \SER_CMD_WORD_F[1]_net_1\);
    
    START_RISE_RNO : NOR2B
      port map(A => \CLK40M_GEN_DEL0\, B => CLK_40M_GL, Y => 
        N_START_RISE);
    
    \SER_CMD_WORD_R_RNO[2]\ : MX2
      port map(A => \SER_CMD_WORD_R[1]_net_1\, B => ELK_TX_DAT(5), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_R[2]\);
    
    SER_OUT_FDEL : DFN1C0
      port map(D => \SER_OUT_FI\, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_8, Q => ELK_OUT_F);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity DDR_BIDIR_LVDS_DUAL_CLK_15 is

    port( DCB_SALT_SEL_c_i : in    std_logic;
          ELK15_DAT_P      : inout std_logic := 'Z';
          ELK15_DAT_N      : inout std_logic := 'Z';
          ELK_OUT_R        : in    std_logic;
          ELK_OUT_F        : in    std_logic;
          CCC_160M_FXD     : in    std_logic;
          CCC_160M_ADJ     : in    std_logic;
          ELK_IN_DDR_R     : out   std_logic;
          ELK_IN_DDR_F     : out   std_logic
        );

end DDR_BIDIR_LVDS_DUAL_CLK_15;

architecture DEF_ARCH of DDR_BIDIR_LVDS_DUAL_CLK_15 is 

  component DDR_REG
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          QR  : out   std_logic;
          QF  : out   std_logic
        );
  end component;

  component DDR_OUT
    port( DR  : in    std_logic := 'U';
          DF  : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component BIBUF_LVDS
    port( PADP : inout   std_logic;
          PADN : inout   std_logic;
          D    : in    std_logic := 'U';
          E    : in    std_logic := 'U';
          Y    : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal DDR_BIDIR_LVDS_DUAL_CLK_15_GND, BIBUF_LVDS_0_Y, 
        DDR_OUT_0_Q, \VCC\ : std_logic;

begin 


    DDR_REG_0 : DDR_REG
      port map(D => BIBUF_LVDS_0_Y, CLK => CCC_160M_ADJ, CLR => 
        DDR_BIDIR_LVDS_DUAL_CLK_15_GND, QR => ELK_IN_DDR_R, QF
         => ELK_IN_DDR_F);
    
    DDR_OUT_0 : DDR_OUT
      port map(DR => ELK_OUT_R, DF => ELK_OUT_F, CLK => 
        CCC_160M_FXD, CLR => DDR_BIDIR_LVDS_DUAL_CLK_15_GND, Q
         => DDR_OUT_0_Q);
    
    BIBUF_LVDS_0 : BIBUF_LVDS
      port map(PADP => ELK15_DAT_P, PADN => ELK15_DAT_N, D => 
        DDR_OUT_0_Q, E => DCB_SALT_SEL_c_i, Y => BIBUF_LVDS_0_Y);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    GND_i : GND
      port map(Y => DDR_BIDIR_LVDS_DUAL_CLK_15_GND);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SYNC_DAT_SEL_15 is

    port( ELK_TX_DAT                : out   std_logic_vector(7 downto 0);
          PATT_ELK_DAT_15           : in    std_logic_vector(7 downto 0);
          OP_MODE_c_6_0             : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_8 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_7 : in    std_logic;
          CLK_40M_GL                : in    std_logic
        );

end SYNC_DAT_SEL_15;

architecture DEF_ARCH of SYNC_DAT_SEL_15 is 

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \N_SERDAT[0]\, \N_SERDAT[1]\, \N_SERDAT[2]\, 
        \N_SERDAT[3]\, \N_SERDAT[4]\, \N_SERDAT[5]\, 
        \N_SERDAT[6]\, \N_SERDAT[7]\, \GND\, \VCC\ : std_logic;

begin 


    \SERDAT_RNO[4]\ : NOR2A
      port map(A => PATT_ELK_DAT_15(4), B => OP_MODE_c_6_0, Y => 
        \N_SERDAT[4]\);
    
    \SERDAT_RNO[0]\ : NOR2A
      port map(A => PATT_ELK_DAT_15(0), B => OP_MODE_c_6_0, Y => 
        \N_SERDAT[0]\);
    
    \SERDAT[6]\ : DFN1C0
      port map(D => \N_SERDAT[6]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_8, Q => ELK_TX_DAT(6));
    
    \SERDAT[4]\ : DFN1C0
      port map(D => \N_SERDAT[4]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_8, Q => ELK_TX_DAT(4));
    
    \SERDAT_RNO[7]\ : OR2
      port map(A => PATT_ELK_DAT_15(7), B => OP_MODE_c_6_0, Y => 
        \N_SERDAT[7]\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \SERDAT_RNO[3]\ : OR2
      port map(A => PATT_ELK_DAT_15(3), B => OP_MODE_c_6_0, Y => 
        \N_SERDAT[3]\);
    
    \SERDAT_RNO[2]\ : OR2
      port map(A => PATT_ELK_DAT_15(2), B => OP_MODE_c_6_0, Y => 
        \N_SERDAT[2]\);
    
    \SERDAT[5]\ : DFN1C0
      port map(D => \N_SERDAT[5]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_8, Q => ELK_TX_DAT(5));
    
    \SERDAT[7]\ : DFN1C0
      port map(D => \N_SERDAT[7]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_8, Q => ELK_TX_DAT(7));
    
    GND_i : GND
      port map(Y => \GND\);
    
    \SERDAT_RNO[5]\ : NOR2A
      port map(A => PATT_ELK_DAT_15(5), B => OP_MODE_c_6_0, Y => 
        \N_SERDAT[5]\);
    
    \SERDAT[0]\ : DFN1C0
      port map(D => \N_SERDAT[0]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_7, Q => ELK_TX_DAT(0));
    
    \SERDAT_RNO[6]\ : NOR2A
      port map(A => PATT_ELK_DAT_15(6), B => OP_MODE_c_6_0, Y => 
        \N_SERDAT[6]\);
    
    \SERDAT[1]\ : DFN1C0
      port map(D => \N_SERDAT[1]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_8, Q => ELK_TX_DAT(1));
    
    \SERDAT_RNO[1]\ : OR2
      port map(A => PATT_ELK_DAT_15(1), B => OP_MODE_c_6_0, Y => 
        \N_SERDAT[1]\);
    
    \SERDAT[3]\ : DFN1C0
      port map(D => \N_SERDAT[3]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_8, Q => ELK_TX_DAT(3));
    
    \SERDAT[2]\ : DFN1C0
      port map(D => \N_SERDAT[2]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_8, Q => ELK_TX_DAT(2));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity ELINK_SLAVE_15_10 is

    port( BIT_OS_SEL_1_0            : in    std_logic;
          BIT_OS_SEL_2              : in    std_logic_vector(2 downto 1);
          BIT_OS_SEL_4_0            : in    std_logic;
          BIT_OS_SEL_3              : in    std_logic_vector(1 downto 0);
          ELK_RX_SER_WORD_15        : out   std_logic_vector(7 downto 0);
          OP_MODE_c_6_0             : in    std_logic;
          PATT_ELK_DAT_15           : in    std_logic_vector(7 downto 0);
          MASTER_DCB_POR_B_i_0_i    : in    std_logic;
          ELK15_DAT_N               : inout std_logic := 'Z';
          ELK15_DAT_P               : inout std_logic := 'Z';
          DCB_SALT_SEL_c_i          : in    std_logic;
          CCC_160M_FXD              : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_5 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_9 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_1 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_6 : in    std_logic;
          CLK_40M_GL                : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_7 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_8 : in    std_logic;
          DEV_RST_B_c_1             : in    std_logic;
          CCC_160M_ADJ              : in    std_logic
        );

end ELINK_SLAVE_15_10;

architecture DEF_ARCH of ELINK_SLAVE_15_10 is 

  component SLAVE_DES320S_1_17_13
    port( ELK_RX_SER_WORD_15     : out   std_logic_vector(7 downto 0);
          BIT_OS_SEL_3           : in    std_logic_vector(1 downto 0) := (others => 'U');
          BIT_OS_SEL_4_0         : in    std_logic := 'U';
          BIT_OS_SEL_2           : in    std_logic_vector(2 downto 1) := (others => 'U');
          BIT_OS_SEL_1_0         : in    std_logic := 'U';
          CLK_40M_GL             : in    std_logic := 'U';
          CCC_160M_FXD           : in    std_logic := 'U';
          ELK_IN_R               : in    std_logic := 'U';
          ELK_IN_F               : in    std_logic := 'U';
          MASTER_DCB_POR_B_i_0_i : in    std_logic := 'U';
          CCC_160M_ADJ           : in    std_logic := 'U'
        );
  end component;

  component SER320M_3_34_15
    port( ELK_TX_DAT                : in    std_logic_vector(7 downto 0) := (others => 'U');
          MASTER_SALT_POR_B_i_0_i_6 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_1 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_9 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_5 : in    std_logic := 'U';
          ELK_OUT_R                 : out   std_logic;
          ELK_OUT_F                 : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_8 : in    std_logic := 'U';
          CCC_160M_FXD              : in    std_logic := 'U';
          CLK_40M_GL                : in    std_logic := 'U'
        );
  end component;

  component DDR_BIDIR_LVDS_DUAL_CLK_15
    port( DCB_SALT_SEL_c_i : in    std_logic := 'U';
          ELK15_DAT_P      : inout   std_logic;
          ELK15_DAT_N      : inout   std_logic;
          ELK_OUT_R        : in    std_logic := 'U';
          ELK_OUT_F        : in    std_logic := 'U';
          CCC_160M_FXD     : in    std_logic := 'U';
          CCC_160M_ADJ     : in    std_logic := 'U';
          ELK_IN_DDR_R     : out   std_logic;
          ELK_IN_DDR_F     : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component SYNC_DAT_SEL_15
    port( ELK_TX_DAT                : out   std_logic_vector(7 downto 0);
          PATT_ELK_DAT_15           : in    std_logic_vector(7 downto 0) := (others => 'U');
          OP_MODE_c_6_0             : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_8 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_7 : in    std_logic := 'U';
          CLK_40M_GL                : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \ELK_IN_F\, ELK_IN_DDR_F, \ELK_IN_R\, ELK_IN_DDR_R, 
        \ELK_TX_DAT[0]\, \ELK_TX_DAT[1]\, \ELK_TX_DAT[2]\, 
        \ELK_TX_DAT[3]\, \ELK_TX_DAT[4]\, \ELK_TX_DAT[5]\, 
        \ELK_TX_DAT[6]\, \ELK_TX_DAT[7]\, ELK_OUT_R, ELK_OUT_F, 
        \GND\, \VCC\ : std_logic;

    for all : SLAVE_DES320S_1_17_13
	Use entity work.SLAVE_DES320S_1_17_13(DEF_ARCH);
    for all : SER320M_3_34_15
	Use entity work.SER320M_3_34_15(DEF_ARCH);
    for all : DDR_BIDIR_LVDS_DUAL_CLK_15
	Use entity work.DDR_BIDIR_LVDS_DUAL_CLK_15(DEF_ARCH);
    for all : SYNC_DAT_SEL_15
	Use entity work.SYNC_DAT_SEL_15(DEF_ARCH);
begin 


    U_SLAVE_1ELK : SLAVE_DES320S_1_17_13
      port map(ELK_RX_SER_WORD_15(7) => ELK_RX_SER_WORD_15(7), 
        ELK_RX_SER_WORD_15(6) => ELK_RX_SER_WORD_15(6), 
        ELK_RX_SER_WORD_15(5) => ELK_RX_SER_WORD_15(5), 
        ELK_RX_SER_WORD_15(4) => ELK_RX_SER_WORD_15(4), 
        ELK_RX_SER_WORD_15(3) => ELK_RX_SER_WORD_15(3), 
        ELK_RX_SER_WORD_15(2) => ELK_RX_SER_WORD_15(2), 
        ELK_RX_SER_WORD_15(1) => ELK_RX_SER_WORD_15(1), 
        ELK_RX_SER_WORD_15(0) => ELK_RX_SER_WORD_15(0), 
        BIT_OS_SEL_3(1) => BIT_OS_SEL_3(1), BIT_OS_SEL_3(0) => 
        BIT_OS_SEL_3(0), BIT_OS_SEL_4_0 => BIT_OS_SEL_4_0, 
        BIT_OS_SEL_2(2) => BIT_OS_SEL_2(2), BIT_OS_SEL_2(1) => 
        BIT_OS_SEL_2(1), BIT_OS_SEL_1_0 => BIT_OS_SEL_1_0, 
        CLK_40M_GL => CLK_40M_GL, CCC_160M_FXD => CCC_160M_FXD, 
        ELK_IN_R => \ELK_IN_R\, ELK_IN_F => \ELK_IN_F\, 
        MASTER_DCB_POR_B_i_0_i => MASTER_DCB_POR_B_i_0_i, 
        CCC_160M_ADJ => CCC_160M_ADJ);
    
    U_ELK1_CMD_TX : SER320M_3_34_15
      port map(ELK_TX_DAT(7) => \ELK_TX_DAT[7]\, ELK_TX_DAT(6)
         => \ELK_TX_DAT[6]\, ELK_TX_DAT(5) => \ELK_TX_DAT[5]\, 
        ELK_TX_DAT(4) => \ELK_TX_DAT[4]\, ELK_TX_DAT(3) => 
        \ELK_TX_DAT[3]\, ELK_TX_DAT(2) => \ELK_TX_DAT[2]\, 
        ELK_TX_DAT(1) => \ELK_TX_DAT[1]\, ELK_TX_DAT(0) => 
        \ELK_TX_DAT[0]\, MASTER_SALT_POR_B_i_0_i_6 => 
        MASTER_SALT_POR_B_i_0_i_6, MASTER_SALT_POR_B_i_0_i_1 => 
        MASTER_SALT_POR_B_i_0_i_1, MASTER_SALT_POR_B_i_0_i_9 => 
        MASTER_SALT_POR_B_i_0_i_9, MASTER_SALT_POR_B_i_0_i_5 => 
        MASTER_SALT_POR_B_i_0_i_5, ELK_OUT_R => ELK_OUT_R, 
        ELK_OUT_F => ELK_OUT_F, MASTER_SALT_POR_B_i_0_i_8 => 
        MASTER_SALT_POR_B_i_0_i_8, CCC_160M_FXD => CCC_160M_FXD, 
        CLK_40M_GL => CLK_40M_GL);
    
    U_DDR_ELK1 : DDR_BIDIR_LVDS_DUAL_CLK_15
      port map(DCB_SALT_SEL_c_i => DCB_SALT_SEL_c_i, ELK15_DAT_P
         => ELK15_DAT_P, ELK15_DAT_N => ELK15_DAT_N, ELK_OUT_R
         => ELK_OUT_R, ELK_OUT_F => ELK_OUT_F, CCC_160M_FXD => 
        CCC_160M_FXD, CCC_160M_ADJ => CCC_160M_ADJ, ELK_IN_DDR_R
         => ELK_IN_DDR_R, ELK_IN_DDR_F => ELK_IN_DDR_F);
    
    ELK_IN_F : DFN1C0
      port map(D => ELK_IN_DDR_F, CLK => CCC_160M_ADJ, CLR => 
        DEV_RST_B_c_1, Q => \ELK_IN_F\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    U_ELK1_SERDAT_SOURCE : SYNC_DAT_SEL_15
      port map(ELK_TX_DAT(7) => \ELK_TX_DAT[7]\, ELK_TX_DAT(6)
         => \ELK_TX_DAT[6]\, ELK_TX_DAT(5) => \ELK_TX_DAT[5]\, 
        ELK_TX_DAT(4) => \ELK_TX_DAT[4]\, ELK_TX_DAT(3) => 
        \ELK_TX_DAT[3]\, ELK_TX_DAT(2) => \ELK_TX_DAT[2]\, 
        ELK_TX_DAT(1) => \ELK_TX_DAT[1]\, ELK_TX_DAT(0) => 
        \ELK_TX_DAT[0]\, PATT_ELK_DAT_15(7) => PATT_ELK_DAT_15(7), 
        PATT_ELK_DAT_15(6) => PATT_ELK_DAT_15(6), 
        PATT_ELK_DAT_15(5) => PATT_ELK_DAT_15(5), 
        PATT_ELK_DAT_15(4) => PATT_ELK_DAT_15(4), 
        PATT_ELK_DAT_15(3) => PATT_ELK_DAT_15(3), 
        PATT_ELK_DAT_15(2) => PATT_ELK_DAT_15(2), 
        PATT_ELK_DAT_15(1) => PATT_ELK_DAT_15(1), 
        PATT_ELK_DAT_15(0) => PATT_ELK_DAT_15(0), OP_MODE_c_6_0
         => OP_MODE_c_6_0, MASTER_SALT_POR_B_i_0_i_8 => 
        MASTER_SALT_POR_B_i_0_i_8, MASTER_SALT_POR_B_i_0_i_7 => 
        MASTER_SALT_POR_B_i_0_i_7, CLK_40M_GL => CLK_40M_GL);
    
    ELK_IN_R : DFN1C0
      port map(D => ELK_IN_DDR_R, CLK => CCC_160M_ADJ, CLR => 
        DEV_RST_B_c_1, Q => \ELK_IN_R\);
    
    GND_i : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity BIDIR_LVDS_IO is

    port( EXT_INT_REF_SEL_c : in    std_logic;
          CLK40M_10NS_REF   : in    std_logic;
          CLK_40M_BUF_RECD  : out   std_logic;
          BIDIR_CLK40M_P    : inout std_logic := 'Z';
          BIDIR_CLK40M_N    : inout std_logic := 'Z'
        );

end BIDIR_LVDS_IO;

architecture DEF_ARCH of BIDIR_LVDS_IO is 

  component INV
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component BIBUF_LVDS
    port( PADP : inout   std_logic;
          PADN : inout   std_logic;
          D    : in    std_logic := 'U';
          E    : in    std_logic := 'U';
          Y    : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal TrienAux, \GND\, \VCC\ : std_logic;

begin 


    Inv_Tri : INV
      port map(A => EXT_INT_REF_SEL_c, Y => TrienAux);
    
    \BIBUF_LVDS[0]\ : BIBUF_LVDS
      port map(PADP => BIDIR_CLK40M_P, PADN => BIDIR_CLK40M_N, D
         => CLK40M_10NS_REF, E => TrienAux, Y => CLK_40M_BUF_RECD);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    GND_i : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity LVDS_BUFOUT is

    port( CLK_40M_BUF_RECD : in    std_logic;
          TX_CLK40M_P      : out   std_logic;
          TX_CLK40M_N      : out   std_logic
        );

end LVDS_BUFOUT;

architecture DEF_ARCH of LVDS_BUFOUT is 

  component OUTBUF_LVDS
    port( D    : in    std_logic := 'U';
          PADP : out   std_logic;
          PADN : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \GND\, \VCC\ : std_logic;

begin 


    \OUTBUF_LVDS[0]\ : OUTBUF_LVDS
      port map(D => CLK_40M_BUF_RECD, PADP => TX_CLK40M_P, PADN
         => TX_CLK40M_N);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    GND_i : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SLAVE_DES320S_1_17_3 is

    port( ELK_RX_SER_WORD_5      : out   std_logic_vector(7 downto 0);
          BIT_OS_SEL_0_0         : in    std_logic;
          BIT_OS_SEL_0_d0        : in    std_logic;
          BIT_OS_SEL_7_0         : in    std_logic;
          BIT_OS_SEL_6           : in    std_logic_vector(2 downto 1);
          BIT_OS_SEL_5           : in    std_logic_vector(2 downto 1);
          CLK_40M_GL             : in    std_logic;
          CCC_160M_FXD           : in    std_logic;
          ELK_IN_R               : in    std_logic;
          ELK_IN_F               : in    std_logic;
          MASTER_DCB_POR_B_i_0_i : in    std_logic;
          CCC_160M_ADJ           : in    std_logic
        );

end SLAVE_DES320S_1_17_3;

architecture DEF_ARCH of SLAVE_DES320S_1_17_3 is 

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal N_17, \ARB_BYTE[0]_net_1\, \ARB_BYTE[4]_net_1\, N_18, 
        \ARB_BYTE[1]_net_1\, \ARB_BYTE[5]_net_1\, N_19, 
        \ARB_BYTE[2]_net_1\, \ARB_BYTE[6]_net_1\, N_20, 
        \ARB_BYTE[3]_net_1\, \ARB_BYTE[7]_net_1\, N_21, 
        \ARB_BYTE[8]_net_1\, N_22, \ARB_BYTE[9]_net_1\, N_23, 
        \ARB_BYTE[10]_net_1\, N_24, \ARB_BYTE[11]_net_1\, N_31, 
        \ARB_BYTE[12]_net_1\, N_32, \ARB_BYTE[13]_net_1\, N_33, 
        N_34, N_35, N_36, N_37, N_38, N_39, N_40, N_56, 
        \ARB_BYTE[14]_net_1\, N_64, \N_RECD_SER_WORD[0]\, 
        \N_RECD_SER_WORD[1]\, \N_RECD_SER_WORD[2]\, 
        \N_RECD_SER_WORD[3]\, \N_RECD_SER_WORD[4]\, 
        \N_RECD_SER_WORD[5]\, \N_RECD_SER_WORD[6]\, 
        \N_RECD_SER_WORD[7]\, \ADJ_SER_IN_F_0DEL\, 
        \ADJ_SER_IN_R_0DEL\, \ADJ_SER_IN_F_1DEL\, 
        \ADJ_SER_IN_R_1DEL\, \Q[0]_net_1\, \ADJ_Q[0]_net_1\, 
        \Q[1]_net_1\, \ADJ_Q[1]_net_1\, \Q[2]_net_1\, 
        \ADJ_Q[2]_net_1\, \Q[3]_net_1\, \ADJ_Q[3]_net_1\, 
        \Q[4]_net_1\, \ADJ_Q[4]_net_1\, \Q[5]_net_1\, 
        \ADJ_Q[5]_net_1\, \Q[6]_net_1\, \ADJ_Q[6]_net_1\, 
        \Q[7]_net_1\, \ADJ_Q[7]_net_1\, \Q[8]_net_1\, 
        \ADJ_Q[8]_net_1\, \Q[9]_net_1\, \ADJ_Q[9]_net_1\, 
        \Q[10]_net_1\, \ADJ_Q[10]_net_1\, \Q[11]_net_1\, 
        \ADJ_Q[11]_net_1\, \Q[12]_net_1\, \ADJ_Q[12]_net_1\, 
        \Q[13]_net_1\, \ADJ_Q[13]_net_1\, \Q[14]_net_1\, 
        \ADJ_Q[14]_net_1\, \ARB_WRD_40M_FIXED[0]_net_1\, 
        \ARB_WRD_40M_FIXED[1]_net_1\, 
        \ARB_WRD_40M_FIXED[2]_net_1\, 
        \ARB_WRD_40M_FIXED[3]_net_1\, 
        \ARB_WRD_40M_FIXED[4]_net_1\, 
        \ARB_WRD_40M_FIXED[5]_net_1\, 
        \ARB_WRD_40M_FIXED[6]_net_1\, 
        \ARB_WRD_40M_FIXED[7]_net_1\, 
        \ARB_WRD_40M_FIXED[8]_net_1\, 
        \ARB_WRD_40M_FIXED[9]_net_1\, 
        \ARB_WRD_40M_FIXED[10]_net_1\, 
        \ARB_WRD_40M_FIXED[11]_net_1\, 
        \ARB_WRD_40M_FIXED[12]_net_1\, 
        \ARB_WRD_40M_FIXED[13]_net_1\, 
        \ARB_WRD_40M_FIXED[14]_net_1\, \GND\, \VCC\ : std_logic;

begin 


    \RECD_SER_WORD_RNO[5]\ : MX2
      port map(A => N_38, B => N_39, S => BIT_OS_SEL_0_0, Y => 
        \N_RECD_SER_WORD[5]\);
    
    \ARB_WRD_40M_FIXED[9]\ : DFN1C0
      port map(D => \Q[9]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[9]_net_1\);
    
    \ADJ_Q[4]\ : DFN1C0
      port map(D => \ADJ_Q[2]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[4]_net_1\);
    
    \ARB_BYTE[6]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[6]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[6]_net_1\);
    
    ADJ_SER_IN_F_1DEL : DFN1C0
      port map(D => \ADJ_SER_IN_F_0DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_F_1DEL\);
    
    \ARB_BYTE[0]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[0]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[0]_net_1\);
    
    \ARB_BYTE_RNIV7F21[6]\ : MX2
      port map(A => N_23, B => N_31, S => BIT_OS_SEL_6(1), Y => 
        N_39);
    
    \Q[11]\ : DFN1C0
      port map(D => \ADJ_Q[11]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[11]_net_1\);
    
    \ADJ_Q[8]\ : DFN1C0
      port map(D => \ADJ_Q[6]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[8]_net_1\);
    
    \ADJ_Q[6]\ : DFN1C0
      port map(D => \ADJ_Q[4]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[6]_net_1\);
    
    \ARB_BYTE_RNI1JGF[2]\ : MX2
      port map(A => N_19, B => N_21, S => BIT_OS_SEL_6(1), Y => 
        N_35);
    
    \ADJ_Q[12]\ : DFN1C0
      port map(D => \ADJ_Q[10]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[12]_net_1\);
    
    \RECD_SER_WORD_RNO_1[0]\ : MX2
      port map(A => \ARB_BYTE[0]_net_1\, B => \ARB_BYTE[4]_net_1\, 
        S => BIT_OS_SEL_5(2), Y => N_17);
    
    \Q[1]\ : DFN1C0
      port map(D => \ADJ_Q[1]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[1]_net_1\);
    
    \ARB_BYTE_RNISBDE[1]\ : MX2
      port map(A => N_18, B => N_20, S => BIT_OS_SEL_5(1), Y => 
        N_34);
    
    \ARB_BYTE[4]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[4]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[4]_net_1\);
    
    \ADJ_Q[2]\ : DFN1C0
      port map(D => \ADJ_Q[0]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[2]_net_1\);
    
    \RECD_SER_WORD_RNO_1[7]\ : MX2
      port map(A => \ARB_BYTE[10]_net_1\, B => 
        \ARB_BYTE[14]_net_1\, S => BIT_OS_SEL_7_0, Y => N_56);
    
    \RECD_SER_WORD[4]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[4]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_5(4));
    
    \Q[5]\ : DFN1C0
      port map(D => \ADJ_Q[5]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[5]_net_1\);
    
    \ARB_BYTE_RNI5NGF[3]\ : MX2
      port map(A => N_20, B => N_22, S => BIT_OS_SEL_6(1), Y => 
        N_36);
    
    \ADJ_Q[11]\ : DFN1C0
      port map(D => \ADJ_Q[9]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[11]_net_1\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \ADJ_Q[3]\ : DFN1C0
      port map(D => \ADJ_Q[1]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[3]_net_1\);
    
    \Q[10]\ : DFN1C0
      port map(D => \ADJ_Q[10]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[10]_net_1\);
    
    \ARB_WRD_40M_FIXED[6]\ : DFN1C0
      port map(D => \Q[6]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[6]_net_1\);
    
    \ARB_WRD_40M_FIXED[1]\ : DFN1C0
      port map(D => \Q[1]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[1]_net_1\);
    
    \RECD_SER_WORD[3]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[3]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_5(3));
    
    \RECD_SER_WORD[0]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[0]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_5(0));
    
    \RECD_SER_WORD_RNO[3]\ : MX2
      port map(A => N_36, B => N_37, S => BIT_OS_SEL_0_0, Y => 
        \N_RECD_SER_WORD[3]\);
    
    \Q[0]\ : DFN1C0
      port map(D => \ADJ_Q[0]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[0]_net_1\);
    
    \RECD_SER_WORD_RNO_0[7]\ : MX2
      port map(A => N_31, B => N_56, S => BIT_OS_SEL_0_d0, Y => 
        N_64);
    
    \Q[7]\ : DFN1C0
      port map(D => \ADJ_Q[7]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[7]_net_1\);
    
    \ARB_BYTE[14]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[14]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[14]_net_1\);
    
    \ARB_WRD_40M_FIXED[2]\ : DFN1C0
      port map(D => \Q[2]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[2]_net_1\);
    
    \ARB_WRD_40M_FIXED[14]\ : DFN1C0
      port map(D => \Q[14]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[14]_net_1\);
    
    \RECD_SER_WORD_RNO[2]\ : MX2
      port map(A => N_35, B => N_36, S => BIT_OS_SEL_0_0, Y => 
        \N_RECD_SER_WORD[2]\);
    
    \ARB_BYTE[2]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[2]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[2]_net_1\);
    
    \ADJ_Q[7]\ : DFN1C0
      port map(D => \ADJ_Q[5]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[7]_net_1\);
    
    \ARB_BYTE[8]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[8]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[8]_net_1\);
    
    \RECD_SER_WORD[5]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[5]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_5(5));
    
    \ARB_BYTE[12]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[12]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[12]_net_1\);
    
    \RECD_SER_WORD[1]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[1]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_5(1));
    
    \Q[3]\ : DFN1C0
      port map(D => \ADJ_Q[3]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[3]_net_1\);
    
    ADJ_SER_IN_F_0DEL : DFN1C0
      port map(D => ELK_IN_F, CLK => CCC_160M_ADJ, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_F_0DEL\);
    
    \RECD_SER_WORD_RNO[7]\ : MX2
      port map(A => N_40, B => N_64, S => BIT_OS_SEL_0_0, Y => 
        \N_RECD_SER_WORD[7]\);
    
    \RECD_SER_WORD_RNO[1]\ : MX2
      port map(A => N_34, B => N_35, S => BIT_OS_SEL_0_0, Y => 
        \N_RECD_SER_WORD[1]\);
    
    \ARB_WRD_40M_FIXED[4]\ : DFN1C0
      port map(D => \Q[4]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[4]_net_1\);
    
    \RECD_SER_WORD_RNO[0]\ : MX2
      port map(A => N_33, B => N_34, S => BIT_OS_SEL_0_0, Y => 
        \N_RECD_SER_WORD[0]\);
    
    \Q[6]\ : DFN1C0
      port map(D => \ADJ_Q[6]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[6]_net_1\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \ARB_WRD_40M_FIXED[8]\ : DFN1C0
      port map(D => \Q[8]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[8]_net_1\);
    
    \ARB_BYTE[11]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[11]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[11]_net_1\);
    
    \Q[9]\ : DFN1C0
      port map(D => \ADJ_Q[9]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[9]_net_1\);
    
    \ARB_BYTE_RNIK10P[5]\ : MX2
      port map(A => N_22, B => N_24, S => BIT_OS_SEL_6(1), Y => 
        N_38);
    
    \Q[14]\ : DFN1C0
      port map(D => \ADJ_Q[14]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[14]_net_1\);
    
    \ARB_BYTE_RNIC3C5[5]\ : MX2
      port map(A => \ARB_BYTE[5]_net_1\, B => \ARB_BYTE[9]_net_1\, 
        S => BIT_OS_SEL_6(2), Y => N_22);
    
    ADJ_SER_IN_R_0DEL : DFN1C0
      port map(D => ELK_IN_R, CLK => CCC_160M_ADJ, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_R_0DEL\);
    
    \Q[13]\ : DFN1C0
      port map(D => \ADJ_Q[13]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[13]_net_1\);
    
    \ARB_BYTE[9]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[9]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[9]_net_1\);
    
    ADJ_SER_IN_R_1DEL : DFN1C0
      port map(D => \ADJ_SER_IN_R_0DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_R_1DEL\);
    
    \ARB_BYTE[10]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[10]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[10]_net_1\);
    
    \ARB_BYTE_RNIN9RE[11]\ : MX2
      port map(A => \ARB_BYTE[7]_net_1\, B => 
        \ARB_BYTE[11]_net_1\, S => BIT_OS_SEL_6(2), Y => N_24);
    
    \ARB_BYTE_RNIGTVO[4]\ : MX2
      port map(A => N_21, B => N_23, S => BIT_OS_SEL_6(1), Y => 
        N_37);
    
    \ADJ_Q[9]\ : DFN1C0
      port map(D => \ADJ_Q[7]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[9]_net_1\);
    
    \RECD_SER_WORD[7]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[7]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_5(7));
    
    \ARB_WRD_40M_FIXED[5]\ : DFN1C0
      port map(D => \Q[5]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[5]_net_1\);
    
    \ARB_WRD_40M_FIXED[12]\ : DFN1C0
      port map(D => \Q[12]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[12]_net_1\);
    
    \ARB_WRD_40M_FIXED[11]\ : DFN1C0
      port map(D => \Q[11]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[11]_net_1\);
    
    \ARB_BYTE_RNI3CF21[13]\ : MX2
      port map(A => N_24, B => N_32, S => BIT_OS_SEL_6(1), Y => 
        N_40);
    
    \ARB_BYTE_RNIL7RE[6]\ : MX2
      port map(A => \ARB_BYTE[6]_net_1\, B => 
        \ARB_BYTE[10]_net_1\, S => BIT_OS_SEL_6(2), Y => N_23);
    
    \ARB_WRD_40M_FIXED[0]\ : DFN1C0
      port map(D => \Q[0]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[0]_net_1\);
    
    \ADJ_Q[10]\ : DFN1C0
      port map(D => \ADJ_Q[8]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[10]_net_1\);
    
    \Q[2]\ : DFN1C0
      port map(D => \ADJ_Q[2]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[2]_net_1\);
    
    \ADJ_Q[1]\ : DFN1C0
      port map(D => \ADJ_SER_IN_F_1DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[1]_net_1\);
    
    \RECD_SER_WORD[6]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[6]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_5(6));
    
    \RECD_SER_WORD[2]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[2]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_5(2));
    
    \ADJ_Q[13]\ : DFN1C0
      port map(D => \ADJ_Q[11]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[13]_net_1\);
    
    \ARB_BYTE_RNIRDRE[13]\ : MX2
      port map(A => \ARB_BYTE[9]_net_1\, B => 
        \ARB_BYTE[13]_net_1\, S => BIT_OS_SEL_6(2), Y => N_32);
    
    \Q[8]\ : DFN1C0
      port map(D => \ADJ_Q[8]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[8]_net_1\);
    
    \ARB_BYTE[5]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[5]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[5]_net_1\);
    
    \ADJ_Q[14]\ : DFN1C0
      port map(D => \ADJ_Q[12]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[14]_net_1\);
    
    \RECD_SER_WORD_RNO[4]\ : MX2
      port map(A => N_37, B => N_38, S => BIT_OS_SEL_0_0, Y => 
        \N_RECD_SER_WORD[4]\);
    
    \Q[12]\ : DFN1C0
      port map(D => \ADJ_Q[12]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[12]_net_1\);
    
    \ARB_BYTE[13]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[13]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[13]_net_1\);
    
    \ARB_BYTE_RNIPBRE[12]\ : MX2
      port map(A => \ARB_BYTE[8]_net_1\, B => 
        \ARB_BYTE[12]_net_1\, S => BIT_OS_SEL_6(2), Y => N_31);
    
    \ARB_WRD_40M_FIXED[3]\ : DFN1C0
      port map(D => \Q[3]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[3]_net_1\);
    
    \ARB_BYTE_RNI6TB5[2]\ : MX2
      port map(A => \ARB_BYTE[2]_net_1\, B => \ARB_BYTE[6]_net_1\, 
        S => BIT_OS_SEL_6(2), Y => N_19);
    
    \ARB_BYTE[7]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[7]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[7]_net_1\);
    
    \RECD_SER_WORD_RNO_0[0]\ : MX2
      port map(A => N_17, B => N_19, S => BIT_OS_SEL_5(1), Y => 
        N_33);
    
    \Q[4]\ : DFN1C0
      port map(D => \ADJ_Q[4]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[4]_net_1\);
    
    \ARB_WRD_40M_FIXED[7]\ : DFN1C0
      port map(D => \Q[7]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[7]_net_1\);
    
    \RECD_SER_WORD_RNO[6]\ : MX2
      port map(A => N_39, B => N_40, S => BIT_OS_SEL_0_0, Y => 
        \N_RECD_SER_WORD[6]\);
    
    \ARB_BYTE_RNIA1C5[4]\ : MX2
      port map(A => \ARB_BYTE[4]_net_1\, B => \ARB_BYTE[8]_net_1\, 
        S => BIT_OS_SEL_6(2), Y => N_21);
    
    \ARB_BYTE[3]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[3]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[3]_net_1\);
    
    \ADJ_Q[5]\ : DFN1C0
      port map(D => \ADJ_Q[3]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[5]_net_1\);
    
    \ARB_BYTE[1]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[1]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[1]_net_1\);
    
    \ARB_WRD_40M_FIXED[13]\ : DFN1C0
      port map(D => \Q[13]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[13]_net_1\);
    
    \ARB_BYTE_RNI8VB5[3]\ : MX2
      port map(A => \ARB_BYTE[3]_net_1\, B => \ARB_BYTE[7]_net_1\, 
        S => BIT_OS_SEL_6(2), Y => N_20);
    
    \ARB_BYTE_RNI4RB5[1]\ : MX2
      port map(A => \ARB_BYTE[1]_net_1\, B => \ARB_BYTE[5]_net_1\, 
        S => BIT_OS_SEL_6(2), Y => N_18);
    
    \ADJ_Q[0]\ : DFN1C0
      port map(D => \ADJ_SER_IN_R_1DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[0]_net_1\);
    
    \ARB_WRD_40M_FIXED[10]\ : DFN1C0
      port map(D => \Q[10]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[10]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SER320M_3_34_5 is

    port( ELK_TX_DAT                 : in    std_logic_vector(7 downto 0);
          MASTER_SALT_POR_B_i_0_i_2  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_6  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_14 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_3  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_5  : in    std_logic;
          ELK_OUT_R                  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_8  : in    std_logic;
          ELK_OUT_F                  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_9  : in    std_logic;
          CCC_160M_FXD               : in    std_logic;
          CLK_40M_GL                 : in    std_logic
        );

end SER320M_3_34_5;

architecture DEF_ARCH of SER320M_3_34_5 is 

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \N_SER_CMD_WORD_R[0]\, \START_RISE\, 
        \N_SER_CMD_WORD_F[0]\, \N_SER_CMD_WORD_R[3]\, 
        \SER_CMD_WORD_R[2]_net_1\, \N_SER_CMD_WORD_R[2]\, 
        \SER_CMD_WORD_R[1]_net_1\, \N_SER_CMD_WORD_R[1]\, 
        \SER_CMD_WORD_R[0]_net_1\, \N_SER_CMD_WORD_F[3]\, 
        \SER_CMD_WORD_F[2]_net_1\, \N_SER_CMD_WORD_F[2]\, 
        \SER_CMD_WORD_F[1]_net_1\, \N_SER_CMD_WORD_F[1]\, 
        \SER_CMD_WORD_F[0]_net_1\, N_START_RISE, 
        \CLK40M_GEN_DEL0\, \SER_OUT_FI\, \SER_OUT_RI\, 
        \SER_CMD_WORD_F[3]_net_1\, \SER_CMD_WORD_R[3]_net_1\, 
        \GND\, \VCC\ : std_logic;

begin 


    SER_OUT_FI : DFN1C0
      port map(D => \SER_CMD_WORD_F[3]_net_1\, CLK => 
        CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_14, Q => 
        \SER_OUT_FI\);
    
    \SER_CMD_WORD_F[3]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[3]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_6, Q => 
        \SER_CMD_WORD_F[3]_net_1\);
    
    \SER_CMD_WORD_R[1]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[1]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_2, Q => 
        \SER_CMD_WORD_R[1]_net_1\);
    
    \SER_CMD_WORD_R[2]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[2]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_2, Q => 
        \SER_CMD_WORD_R[2]_net_1\);
    
    \SER_CMD_WORD_R_RNO[3]\ : MX2
      port map(A => \SER_CMD_WORD_R[2]_net_1\, B => ELK_TX_DAT(7), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_R[3]\);
    
    \SER_CMD_WORD_R_RNO[0]\ : NOR2B
      port map(A => \START_RISE\, B => ELK_TX_DAT(1), Y => 
        \N_SER_CMD_WORD_R[0]\);
    
    \SER_CMD_WORD_F[0]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[0]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_5, Q => 
        \SER_CMD_WORD_F[0]_net_1\);
    
    \SER_CMD_WORD_R_RNO[1]\ : MX2
      port map(A => \SER_CMD_WORD_R[0]_net_1\, B => ELK_TX_DAT(3), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_R[1]\);
    
    \SER_CMD_WORD_F_RNO[2]\ : MX2
      port map(A => \SER_CMD_WORD_F[1]_net_1\, B => ELK_TX_DAT(4), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_F[2]\);
    
    \SER_CMD_WORD_F_RNO[3]\ : MX2
      port map(A => \SER_CMD_WORD_F[2]_net_1\, B => ELK_TX_DAT(6), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_F[3]\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    CLK40M_GEN_DEL0 : DFN1C0
      port map(D => CLK_40M_GL, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_9, Q => \CLK40M_GEN_DEL0\);
    
    SER_OUT_RI : DFN1C0
      port map(D => \SER_CMD_WORD_R[3]_net_1\, CLK => 
        CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_14, Q => 
        \SER_OUT_RI\);
    
    \SER_CMD_WORD_F[2]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[2]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_6, Q => 
        \SER_CMD_WORD_F[2]_net_1\);
    
    \SER_CMD_WORD_F_RNO[1]\ : MX2
      port map(A => \SER_CMD_WORD_F[0]_net_1\, B => ELK_TX_DAT(2), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_F[1]\);
    
    \SER_CMD_WORD_R[0]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[0]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_2, Q => 
        \SER_CMD_WORD_R[0]_net_1\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    START_RISE : DFN1C0
      port map(D => N_START_RISE, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_3, Q => \START_RISE\);
    
    \SER_CMD_WORD_R[3]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[3]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_2, Q => 
        \SER_CMD_WORD_R[3]_net_1\);
    
    \SER_CMD_WORD_F_RNO[0]\ : NOR2B
      port map(A => \START_RISE\, B => ELK_TX_DAT(0), Y => 
        \N_SER_CMD_WORD_F[0]\);
    
    SER_OUT_RDEL : DFN1C0
      port map(D => \SER_OUT_RI\, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_5, Q => ELK_OUT_R);
    
    \SER_CMD_WORD_F[1]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[1]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_5, Q => 
        \SER_CMD_WORD_F[1]_net_1\);
    
    START_RISE_RNO : NOR2B
      port map(A => \CLK40M_GEN_DEL0\, B => CLK_40M_GL, Y => 
        N_START_RISE);
    
    \SER_CMD_WORD_R_RNO[2]\ : MX2
      port map(A => \SER_CMD_WORD_R[1]_net_1\, B => ELK_TX_DAT(5), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_R[2]\);
    
    SER_OUT_FDEL : DFN1C0
      port map(D => \SER_OUT_FI\, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_8, Q => ELK_OUT_F);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity DDR_BIDIR_LVDS_DUAL_CLK_5 is

    port( DCB_SALT_SEL_c_i : in    std_logic;
          ELK5_DAT_P       : inout std_logic := 'Z';
          ELK5_DAT_N       : inout std_logic := 'Z';
          ELK_OUT_R        : in    std_logic;
          ELK_OUT_F        : in    std_logic;
          CCC_160M_FXD     : in    std_logic;
          CCC_160M_ADJ     : in    std_logic;
          ELK_IN_DDR_R     : out   std_logic;
          ELK_IN_DDR_F     : out   std_logic
        );

end DDR_BIDIR_LVDS_DUAL_CLK_5;

architecture DEF_ARCH of DDR_BIDIR_LVDS_DUAL_CLK_5 is 

  component DDR_REG
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          QR  : out   std_logic;
          QF  : out   std_logic
        );
  end component;

  component DDR_OUT
    port( DR  : in    std_logic := 'U';
          DF  : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component BIBUF_LVDS
    port( PADP : inout   std_logic;
          PADN : inout   std_logic;
          D    : in    std_logic := 'U';
          E    : in    std_logic := 'U';
          Y    : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal DDR_BIDIR_LVDS_DUAL_CLK_5_GND, BIBUF_LVDS_0_Y, 
        DDR_OUT_0_Q, \VCC\ : std_logic;

begin 


    DDR_REG_0 : DDR_REG
      port map(D => BIBUF_LVDS_0_Y, CLK => CCC_160M_ADJ, CLR => 
        DDR_BIDIR_LVDS_DUAL_CLK_5_GND, QR => ELK_IN_DDR_R, QF => 
        ELK_IN_DDR_F);
    
    DDR_OUT_0 : DDR_OUT
      port map(DR => ELK_OUT_R, DF => ELK_OUT_F, CLK => 
        CCC_160M_FXD, CLR => DDR_BIDIR_LVDS_DUAL_CLK_5_GND, Q => 
        DDR_OUT_0_Q);
    
    BIBUF_LVDS_0 : BIBUF_LVDS
      port map(PADP => ELK5_DAT_P, PADN => ELK5_DAT_N, D => 
        DDR_OUT_0_Q, E => DCB_SALT_SEL_c_i, Y => BIBUF_LVDS_0_Y);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    GND_i : GND
      port map(Y => DDR_BIDIR_LVDS_DUAL_CLK_5_GND);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SYNC_DAT_SEL_5 is

    port( ELK_TX_DAT                 : out   std_logic_vector(7 downto 0);
          PATT_ELK_DAT_5             : in    std_logic_vector(7 downto 0);
          OP_MODE_c_5_0              : in    std_logic;
          OP_MODE_c_4_0              : in    std_logic;
          MASTER_SALT_POR_B_i_0_i    : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_17 : in    std_logic;
          CLK_40M_GL                 : in    std_logic
        );

end SYNC_DAT_SEL_5;

architecture DEF_ARCH of SYNC_DAT_SEL_5 is 

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \N_SERDAT[0]\, \N_SERDAT[1]\, \N_SERDAT[2]\, 
        \N_SERDAT[3]\, \N_SERDAT[4]\, \N_SERDAT[5]\, 
        \N_SERDAT[6]\, \N_SERDAT[7]\, \GND\, \VCC\ : std_logic;

begin 


    \SERDAT_RNO[4]\ : NOR2A
      port map(A => PATT_ELK_DAT_5(4), B => OP_MODE_c_4_0, Y => 
        \N_SERDAT[4]\);
    
    \SERDAT_RNO[0]\ : NOR2A
      port map(A => PATT_ELK_DAT_5(0), B => OP_MODE_c_4_0, Y => 
        \N_SERDAT[0]\);
    
    \SERDAT[6]\ : DFN1C0
      port map(D => \N_SERDAT[6]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i, Q => ELK_TX_DAT(6));
    
    \SERDAT[4]\ : DFN1C0
      port map(D => \N_SERDAT[4]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i, Q => ELK_TX_DAT(4));
    
    \SERDAT_RNO[7]\ : OR2
      port map(A => PATT_ELK_DAT_5(7), B => OP_MODE_c_5_0, Y => 
        \N_SERDAT[7]\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \SERDAT_RNO[3]\ : OR2
      port map(A => PATT_ELK_DAT_5(3), B => OP_MODE_c_4_0, Y => 
        \N_SERDAT[3]\);
    
    \SERDAT_RNO[2]\ : OR2
      port map(A => PATT_ELK_DAT_5(2), B => OP_MODE_c_4_0, Y => 
        \N_SERDAT[2]\);
    
    \SERDAT[5]\ : DFN1C0
      port map(D => \N_SERDAT[5]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i, Q => ELK_TX_DAT(5));
    
    \SERDAT[7]\ : DFN1C0
      port map(D => \N_SERDAT[7]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i, Q => ELK_TX_DAT(7));
    
    GND_i : GND
      port map(Y => \GND\);
    
    \SERDAT_RNO[5]\ : NOR2A
      port map(A => PATT_ELK_DAT_5(5), B => OP_MODE_c_4_0, Y => 
        \N_SERDAT[5]\);
    
    \SERDAT[0]\ : DFN1C0
      port map(D => \N_SERDAT[0]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_17, Q => ELK_TX_DAT(0));
    
    \SERDAT_RNO[6]\ : NOR2A
      port map(A => PATT_ELK_DAT_5(6), B => OP_MODE_c_5_0, Y => 
        \N_SERDAT[6]\);
    
    \SERDAT[1]\ : DFN1C0
      port map(D => \N_SERDAT[1]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_17, Q => ELK_TX_DAT(1));
    
    \SERDAT_RNO[1]\ : OR2
      port map(A => PATT_ELK_DAT_5(1), B => OP_MODE_c_4_0, Y => 
        \N_SERDAT[1]\);
    
    \SERDAT[3]\ : DFN1C0
      port map(D => \N_SERDAT[3]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_17, Q => ELK_TX_DAT(3));
    
    \SERDAT[2]\ : DFN1C0
      port map(D => \N_SERDAT[2]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_17, Q => ELK_TX_DAT(2));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity ELINK_SLAVE_15_0 is

    port( BIT_OS_SEL_5               : in    std_logic_vector(2 downto 1);
          BIT_OS_SEL_6               : in    std_logic_vector(2 downto 1);
          BIT_OS_SEL_7_0             : in    std_logic;
          BIT_OS_SEL_0_d0            : in    std_logic;
          BIT_OS_SEL_0_0             : in    std_logic;
          ELK_RX_SER_WORD_5          : out   std_logic_vector(7 downto 0);
          OP_MODE_c_4_0              : in    std_logic;
          OP_MODE_c_5_0              : in    std_logic;
          PATT_ELK_DAT_5             : in    std_logic_vector(7 downto 0);
          MASTER_DCB_POR_B_i_0_i     : in    std_logic;
          ELK5_DAT_N                 : inout std_logic := 'Z';
          ELK5_DAT_P                 : inout std_logic := 'Z';
          DCB_SALT_SEL_c_i           : in    std_logic;
          CCC_160M_FXD               : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_9  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_8  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_5  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_3  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_14 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_6  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_2  : in    std_logic;
          CLK_40M_GL                 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_17 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i    : in    std_logic;
          DEV_RST_B_c                : in    std_logic;
          CCC_160M_ADJ               : in    std_logic
        );

end ELINK_SLAVE_15_0;

architecture DEF_ARCH of ELINK_SLAVE_15_0 is 

  component SLAVE_DES320S_1_17_3
    port( ELK_RX_SER_WORD_5      : out   std_logic_vector(7 downto 0);
          BIT_OS_SEL_0_0         : in    std_logic := 'U';
          BIT_OS_SEL_0_d0        : in    std_logic := 'U';
          BIT_OS_SEL_7_0         : in    std_logic := 'U';
          BIT_OS_SEL_6           : in    std_logic_vector(2 downto 1) := (others => 'U');
          BIT_OS_SEL_5           : in    std_logic_vector(2 downto 1) := (others => 'U');
          CLK_40M_GL             : in    std_logic := 'U';
          CCC_160M_FXD           : in    std_logic := 'U';
          ELK_IN_R               : in    std_logic := 'U';
          ELK_IN_F               : in    std_logic := 'U';
          MASTER_DCB_POR_B_i_0_i : in    std_logic := 'U';
          CCC_160M_ADJ           : in    std_logic := 'U'
        );
  end component;

  component SER320M_3_34_5
    port( ELK_TX_DAT                 : in    std_logic_vector(7 downto 0) := (others => 'U');
          MASTER_SALT_POR_B_i_0_i_2  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_6  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_14 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_3  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_5  : in    std_logic := 'U';
          ELK_OUT_R                  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_8  : in    std_logic := 'U';
          ELK_OUT_F                  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_9  : in    std_logic := 'U';
          CCC_160M_FXD               : in    std_logic := 'U';
          CLK_40M_GL                 : in    std_logic := 'U'
        );
  end component;

  component DDR_BIDIR_LVDS_DUAL_CLK_5
    port( DCB_SALT_SEL_c_i : in    std_logic := 'U';
          ELK5_DAT_P       : inout   std_logic;
          ELK5_DAT_N       : inout   std_logic;
          ELK_OUT_R        : in    std_logic := 'U';
          ELK_OUT_F        : in    std_logic := 'U';
          CCC_160M_FXD     : in    std_logic := 'U';
          CCC_160M_ADJ     : in    std_logic := 'U';
          ELK_IN_DDR_R     : out   std_logic;
          ELK_IN_DDR_F     : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component SYNC_DAT_SEL_5
    port( ELK_TX_DAT                 : out   std_logic_vector(7 downto 0);
          PATT_ELK_DAT_5             : in    std_logic_vector(7 downto 0) := (others => 'U');
          OP_MODE_c_5_0              : in    std_logic := 'U';
          OP_MODE_c_4_0              : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i    : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_17 : in    std_logic := 'U';
          CLK_40M_GL                 : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \ELK_IN_F\, ELK_IN_DDR_F, \ELK_IN_R\, ELK_IN_DDR_R, 
        \ELK_TX_DAT[0]\, \ELK_TX_DAT[1]\, \ELK_TX_DAT[2]\, 
        \ELK_TX_DAT[3]\, \ELK_TX_DAT[4]\, \ELK_TX_DAT[5]\, 
        \ELK_TX_DAT[6]\, \ELK_TX_DAT[7]\, ELK_OUT_R, ELK_OUT_F, 
        \GND\, \VCC\ : std_logic;

    for all : SLAVE_DES320S_1_17_3
	Use entity work.SLAVE_DES320S_1_17_3(DEF_ARCH);
    for all : SER320M_3_34_5
	Use entity work.SER320M_3_34_5(DEF_ARCH);
    for all : DDR_BIDIR_LVDS_DUAL_CLK_5
	Use entity work.DDR_BIDIR_LVDS_DUAL_CLK_5(DEF_ARCH);
    for all : SYNC_DAT_SEL_5
	Use entity work.SYNC_DAT_SEL_5(DEF_ARCH);
begin 


    U_SLAVE_1ELK : SLAVE_DES320S_1_17_3
      port map(ELK_RX_SER_WORD_5(7) => ELK_RX_SER_WORD_5(7), 
        ELK_RX_SER_WORD_5(6) => ELK_RX_SER_WORD_5(6), 
        ELK_RX_SER_WORD_5(5) => ELK_RX_SER_WORD_5(5), 
        ELK_RX_SER_WORD_5(4) => ELK_RX_SER_WORD_5(4), 
        ELK_RX_SER_WORD_5(3) => ELK_RX_SER_WORD_5(3), 
        ELK_RX_SER_WORD_5(2) => ELK_RX_SER_WORD_5(2), 
        ELK_RX_SER_WORD_5(1) => ELK_RX_SER_WORD_5(1), 
        ELK_RX_SER_WORD_5(0) => ELK_RX_SER_WORD_5(0), 
        BIT_OS_SEL_0_0 => BIT_OS_SEL_0_0, BIT_OS_SEL_0_d0 => 
        BIT_OS_SEL_0_d0, BIT_OS_SEL_7_0 => BIT_OS_SEL_7_0, 
        BIT_OS_SEL_6(2) => BIT_OS_SEL_6(2), BIT_OS_SEL_6(1) => 
        BIT_OS_SEL_6(1), BIT_OS_SEL_5(2) => BIT_OS_SEL_5(2), 
        BIT_OS_SEL_5(1) => BIT_OS_SEL_5(1), CLK_40M_GL => 
        CLK_40M_GL, CCC_160M_FXD => CCC_160M_FXD, ELK_IN_R => 
        \ELK_IN_R\, ELK_IN_F => \ELK_IN_F\, 
        MASTER_DCB_POR_B_i_0_i => MASTER_DCB_POR_B_i_0_i, 
        CCC_160M_ADJ => CCC_160M_ADJ);
    
    U_ELK1_CMD_TX : SER320M_3_34_5
      port map(ELK_TX_DAT(7) => \ELK_TX_DAT[7]\, ELK_TX_DAT(6)
         => \ELK_TX_DAT[6]\, ELK_TX_DAT(5) => \ELK_TX_DAT[5]\, 
        ELK_TX_DAT(4) => \ELK_TX_DAT[4]\, ELK_TX_DAT(3) => 
        \ELK_TX_DAT[3]\, ELK_TX_DAT(2) => \ELK_TX_DAT[2]\, 
        ELK_TX_DAT(1) => \ELK_TX_DAT[1]\, ELK_TX_DAT(0) => 
        \ELK_TX_DAT[0]\, MASTER_SALT_POR_B_i_0_i_2 => 
        MASTER_SALT_POR_B_i_0_i_2, MASTER_SALT_POR_B_i_0_i_6 => 
        MASTER_SALT_POR_B_i_0_i_6, MASTER_SALT_POR_B_i_0_i_14 => 
        MASTER_SALT_POR_B_i_0_i_14, MASTER_SALT_POR_B_i_0_i_3 => 
        MASTER_SALT_POR_B_i_0_i_3, MASTER_SALT_POR_B_i_0_i_5 => 
        MASTER_SALT_POR_B_i_0_i_5, ELK_OUT_R => ELK_OUT_R, 
        MASTER_SALT_POR_B_i_0_i_8 => MASTER_SALT_POR_B_i_0_i_8, 
        ELK_OUT_F => ELK_OUT_F, MASTER_SALT_POR_B_i_0_i_9 => 
        MASTER_SALT_POR_B_i_0_i_9, CCC_160M_FXD => CCC_160M_FXD, 
        CLK_40M_GL => CLK_40M_GL);
    
    U_DDR_ELK1 : DDR_BIDIR_LVDS_DUAL_CLK_5
      port map(DCB_SALT_SEL_c_i => DCB_SALT_SEL_c_i, ELK5_DAT_P
         => ELK5_DAT_P, ELK5_DAT_N => ELK5_DAT_N, ELK_OUT_R => 
        ELK_OUT_R, ELK_OUT_F => ELK_OUT_F, CCC_160M_FXD => 
        CCC_160M_FXD, CCC_160M_ADJ => CCC_160M_ADJ, ELK_IN_DDR_R
         => ELK_IN_DDR_R, ELK_IN_DDR_F => ELK_IN_DDR_F);
    
    ELK_IN_F : DFN1C0
      port map(D => ELK_IN_DDR_F, CLK => CCC_160M_ADJ, CLR => 
        DEV_RST_B_c, Q => \ELK_IN_F\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    U_ELK1_SERDAT_SOURCE : SYNC_DAT_SEL_5
      port map(ELK_TX_DAT(7) => \ELK_TX_DAT[7]\, ELK_TX_DAT(6)
         => \ELK_TX_DAT[6]\, ELK_TX_DAT(5) => \ELK_TX_DAT[5]\, 
        ELK_TX_DAT(4) => \ELK_TX_DAT[4]\, ELK_TX_DAT(3) => 
        \ELK_TX_DAT[3]\, ELK_TX_DAT(2) => \ELK_TX_DAT[2]\, 
        ELK_TX_DAT(1) => \ELK_TX_DAT[1]\, ELK_TX_DAT(0) => 
        \ELK_TX_DAT[0]\, PATT_ELK_DAT_5(7) => PATT_ELK_DAT_5(7), 
        PATT_ELK_DAT_5(6) => PATT_ELK_DAT_5(6), PATT_ELK_DAT_5(5)
         => PATT_ELK_DAT_5(5), PATT_ELK_DAT_5(4) => 
        PATT_ELK_DAT_5(4), PATT_ELK_DAT_5(3) => PATT_ELK_DAT_5(3), 
        PATT_ELK_DAT_5(2) => PATT_ELK_DAT_5(2), PATT_ELK_DAT_5(1)
         => PATT_ELK_DAT_5(1), PATT_ELK_DAT_5(0) => 
        PATT_ELK_DAT_5(0), OP_MODE_c_5_0 => OP_MODE_c_5_0, 
        OP_MODE_c_4_0 => OP_MODE_c_4_0, MASTER_SALT_POR_B_i_0_i
         => MASTER_SALT_POR_B_i_0_i, MASTER_SALT_POR_B_i_0_i_17
         => MASTER_SALT_POR_B_i_0_i_17, CLK_40M_GL => CLK_40M_GL);
    
    ELK_IN_R : DFN1C0
      port map(D => ELK_IN_DDR_R, CLK => CCC_160M_ADJ, CLR => 
        DEV_RST_B_c, Q => \ELK_IN_R\);
    
    GND_i : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SLAVE_DES320S_1_17_8 is

    port( ELK_RX_SER_WORD_10     : out   std_logic_vector(7 downto 0);
          BIT_OS_SEL_0_0         : in    std_logic;
          BIT_OS_SEL_0_d0        : in    std_logic;
          BIT_OS_SEL_7_0         : in    std_logic;
          BIT_OS_SEL_5           : in    std_logic_vector(2 downto 1);
          BIT_OS_SEL_6_0         : in    std_logic;
          CLK_40M_GL             : in    std_logic;
          CCC_160M_FXD           : in    std_logic;
          ELK_IN_R               : in    std_logic;
          ELK_IN_F               : in    std_logic;
          MASTER_DCB_POR_B_i_0_i : in    std_logic;
          CCC_160M_ADJ           : in    std_logic
        );

end SLAVE_DES320S_1_17_8;

architecture DEF_ARCH of SLAVE_DES320S_1_17_8 is 

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal N_17, \ARB_BYTE[0]_net_1\, \ARB_BYTE[4]_net_1\, N_18, 
        \ARB_BYTE[1]_net_1\, \ARB_BYTE[5]_net_1\, N_19, 
        \ARB_BYTE[2]_net_1\, \ARB_BYTE[6]_net_1\, N_20, 
        \ARB_BYTE[3]_net_1\, \ARB_BYTE[7]_net_1\, N_21, 
        \ARB_BYTE[8]_net_1\, N_22, \ARB_BYTE[9]_net_1\, N_23, 
        \ARB_BYTE[10]_net_1\, N_24, \ARB_BYTE[11]_net_1\, N_31, 
        \ARB_BYTE[12]_net_1\, N_32, \ARB_BYTE[13]_net_1\, N_33, 
        N_34, N_35, N_36, N_37, N_38, N_39, N_40, N_56, 
        \ARB_BYTE[14]_net_1\, N_64, \N_RECD_SER_WORD[0]\, 
        \N_RECD_SER_WORD[1]\, \N_RECD_SER_WORD[2]\, 
        \N_RECD_SER_WORD[3]\, \N_RECD_SER_WORD[4]\, 
        \N_RECD_SER_WORD[5]\, \N_RECD_SER_WORD[6]\, 
        \N_RECD_SER_WORD[7]\, \ADJ_SER_IN_F_0DEL\, 
        \ADJ_SER_IN_R_0DEL\, \ADJ_SER_IN_F_1DEL\, 
        \ADJ_SER_IN_R_1DEL\, \Q[0]_net_1\, \ADJ_Q[0]_net_1\, 
        \Q[1]_net_1\, \ADJ_Q[1]_net_1\, \Q[2]_net_1\, 
        \ADJ_Q[2]_net_1\, \Q[3]_net_1\, \ADJ_Q[3]_net_1\, 
        \Q[4]_net_1\, \ADJ_Q[4]_net_1\, \Q[5]_net_1\, 
        \ADJ_Q[5]_net_1\, \Q[6]_net_1\, \ADJ_Q[6]_net_1\, 
        \Q[7]_net_1\, \ADJ_Q[7]_net_1\, \Q[8]_net_1\, 
        \ADJ_Q[8]_net_1\, \Q[9]_net_1\, \ADJ_Q[9]_net_1\, 
        \Q[10]_net_1\, \ADJ_Q[10]_net_1\, \Q[11]_net_1\, 
        \ADJ_Q[11]_net_1\, \Q[12]_net_1\, \ADJ_Q[12]_net_1\, 
        \Q[13]_net_1\, \ADJ_Q[13]_net_1\, \Q[14]_net_1\, 
        \ADJ_Q[14]_net_1\, \ARB_WRD_40M_FIXED[0]_net_1\, 
        \ARB_WRD_40M_FIXED[1]_net_1\, 
        \ARB_WRD_40M_FIXED[2]_net_1\, 
        \ARB_WRD_40M_FIXED[3]_net_1\, 
        \ARB_WRD_40M_FIXED[4]_net_1\, 
        \ARB_WRD_40M_FIXED[5]_net_1\, 
        \ARB_WRD_40M_FIXED[6]_net_1\, 
        \ARB_WRD_40M_FIXED[7]_net_1\, 
        \ARB_WRD_40M_FIXED[8]_net_1\, 
        \ARB_WRD_40M_FIXED[9]_net_1\, 
        \ARB_WRD_40M_FIXED[10]_net_1\, 
        \ARB_WRD_40M_FIXED[11]_net_1\, 
        \ARB_WRD_40M_FIXED[12]_net_1\, 
        \ARB_WRD_40M_FIXED[13]_net_1\, 
        \ARB_WRD_40M_FIXED[14]_net_1\, \GND\, \VCC\ : std_logic;

begin 


    \RECD_SER_WORD_RNO[5]\ : MX2
      port map(A => N_38, B => N_39, S => BIT_OS_SEL_0_0, Y => 
        \N_RECD_SER_WORD[5]\);
    
    \ARB_WRD_40M_FIXED[9]\ : DFN1C0
      port map(D => \Q[9]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[9]_net_1\);
    
    \ADJ_Q[4]\ : DFN1C0
      port map(D => \ADJ_Q[2]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[4]_net_1\);
    
    \ARB_BYTE[6]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[6]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[6]_net_1\);
    
    ADJ_SER_IN_F_1DEL : DFN1C0
      port map(D => \ADJ_SER_IN_F_0DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_F_1DEL\);
    
    \ARB_BYTE[0]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[0]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[0]_net_1\);
    
    \Q[11]\ : DFN1C0
      port map(D => \ADJ_Q[11]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[11]_net_1\);
    
    \ADJ_Q[8]\ : DFN1C0
      port map(D => \ADJ_Q[6]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[8]_net_1\);
    
    \ARB_BYTE_RNICL9P[10]\ : MX2
      port map(A => \ARB_BYTE[6]_net_1\, B => 
        \ARB_BYTE[10]_net_1\, S => BIT_OS_SEL_5(2), Y => N_23);
    
    \ARB_BYTE_RNIJUCQ[13]\ : MX2
      port map(A => \ARB_BYTE[9]_net_1\, B => 
        \ARB_BYTE[13]_net_1\, S => BIT_OS_SEL_6_0, Y => N_32);
    
    \ADJ_Q[6]\ : DFN1C0
      port map(D => \ADJ_Q[4]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[6]_net_1\);
    
    \ADJ_Q[12]\ : DFN1C0
      port map(D => \ADJ_Q[10]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[12]_net_1\);
    
    \RECD_SER_WORD_RNO_1[0]\ : MX2
      port map(A => \ARB_BYTE[0]_net_1\, B => \ARB_BYTE[4]_net_1\, 
        S => BIT_OS_SEL_5(2), Y => N_17);
    
    \Q[1]\ : DFN1C0
      port map(D => \ADJ_Q[1]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[1]_net_1\);
    
    \ARB_BYTE_RNIEN9P[11]\ : MX2
      port map(A => \ARB_BYTE[7]_net_1\, B => 
        \ARB_BYTE[11]_net_1\, S => BIT_OS_SEL_5(2), Y => N_24);
    
    \ARB_BYTE_RNI1E7T1[11]\ : MX2
      port map(A => N_22, B => N_24, S => BIT_OS_SEL_5(1), Y => 
        N_38);
    
    \ARB_BYTE_RNIV0801[3]\ : MX2
      port map(A => \ARB_BYTE[3]_net_1\, B => \ARB_BYTE[7]_net_1\, 
        S => BIT_OS_SEL_5(2), Y => N_20);
    
    \ARB_BYTE[4]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[4]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[4]_net_1\);
    
    \ARB_BYTE_RNI35801[5]\ : MX2
      port map(A => \ARB_BYTE[5]_net_1\, B => \ARB_BYTE[9]_net_1\, 
        S => BIT_OS_SEL_5(2), Y => N_22);
    
    \ADJ_Q[2]\ : DFN1C0
      port map(D => \ADJ_Q[0]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[2]_net_1\);
    
    \RECD_SER_WORD_RNO_1[7]\ : MX2
      port map(A => \ARB_BYTE[10]_net_1\, B => 
        \ARB_BYTE[14]_net_1\, S => BIT_OS_SEL_7_0, Y => N_56);
    
    \RECD_SER_WORD[4]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[4]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_10(4));
    
    \Q[5]\ : DFN1C0
      port map(D => \ADJ_Q[5]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[5]_net_1\);
    
    \ADJ_Q[11]\ : DFN1C0
      port map(D => \ADJ_Q[9]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[11]_net_1\);
    
    \ARB_BYTE_RNIIN542[3]\ : MX2
      port map(A => N_20, B => N_22, S => BIT_OS_SEL_5(1), Y => 
        N_36);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \ADJ_Q[3]\ : DFN1C0
      port map(D => \ADJ_Q[1]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[3]_net_1\);
    
    \Q[10]\ : DFN1C0
      port map(D => \ADJ_Q[10]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[10]_net_1\);
    
    \ARB_WRD_40M_FIXED[6]\ : DFN1C0
      port map(D => \Q[6]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[6]_net_1\);
    
    \ARB_BYTE_RNI13801[4]\ : MX2
      port map(A => \ARB_BYTE[4]_net_1\, B => \ARB_BYTE[8]_net_1\, 
        S => BIT_OS_SEL_5(2), Y => N_21);
    
    \ARB_WRD_40M_FIXED[1]\ : DFN1C0
      port map(D => \Q[1]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[1]_net_1\);
    
    \RECD_SER_WORD[3]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[3]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_10(3));
    
    \RECD_SER_WORD[0]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[0]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_10(0));
    
    \RECD_SER_WORD_RNO[3]\ : MX2
      port map(A => N_36, B => N_37, S => BIT_OS_SEL_0_0, Y => 
        \N_RECD_SER_WORD[3]\);
    
    \Q[0]\ : DFN1C0
      port map(D => \ADJ_Q[0]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[0]_net_1\);
    
    \RECD_SER_WORD_RNO_0[7]\ : MX2
      port map(A => N_31, B => N_56, S => BIT_OS_SEL_0_d0, Y => 
        N_64);
    
    \Q[7]\ : DFN1C0
      port map(D => \ADJ_Q[7]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[7]_net_1\);
    
    \ARB_BYTE[14]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[14]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[14]_net_1\);
    
    \ARB_WRD_40M_FIXED[2]\ : DFN1C0
      port map(D => \Q[2]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[2]_net_1\);
    
    \ARB_WRD_40M_FIXED[14]\ : DFN1C0
      port map(D => \Q[14]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[14]_net_1\);
    
    \RECD_SER_WORD_RNO[2]\ : MX2
      port map(A => N_35, B => N_36, S => BIT_OS_SEL_0_0, Y => 
        \N_RECD_SER_WORD[2]\);
    
    \ARB_BYTE[2]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[2]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[2]_net_1\);
    
    \ADJ_Q[7]\ : DFN1C0
      port map(D => \ADJ_Q[5]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[7]_net_1\);
    
    \ARB_BYTE[8]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[8]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[8]_net_1\);
    
    \ARB_BYTE_RNIEJ542[2]\ : MX2
      port map(A => N_19, B => N_21, S => BIT_OS_SEL_5(1), Y => 
        N_35);
    
    \RECD_SER_WORD[5]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[5]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_10(5));
    
    \ARB_BYTE[12]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[12]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[12]_net_1\);
    
    \ARB_BYTE_RNITU701[2]\ : MX2
      port map(A => \ARB_BYTE[2]_net_1\, B => \ARB_BYTE[6]_net_1\, 
        S => BIT_OS_SEL_5(2), Y => N_19);
    
    \RECD_SER_WORD[1]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[1]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_10(1));
    
    \Q[3]\ : DFN1C0
      port map(D => \ADJ_Q[3]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[3]_net_1\);
    
    \ARB_BYTE_RNIRS701[1]\ : MX2
      port map(A => \ARB_BYTE[1]_net_1\, B => \ARB_BYTE[5]_net_1\, 
        S => BIT_OS_SEL_5(2), Y => N_18);
    
    ADJ_SER_IN_F_0DEL : DFN1C0
      port map(D => ELK_IN_F, CLK => CCC_160M_ADJ, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_F_0DEL\);
    
    \RECD_SER_WORD_RNO[7]\ : MX2
      port map(A => N_40, B => N_64, S => BIT_OS_SEL_0_0, Y => 
        \N_RECD_SER_WORD[7]\);
    
    \RECD_SER_WORD_RNO[1]\ : MX2
      port map(A => N_34, B => N_35, S => BIT_OS_SEL_0_0, Y => 
        \N_RECD_SER_WORD[1]\);
    
    \ARB_WRD_40M_FIXED[4]\ : DFN1C0
      port map(D => \Q[4]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[4]_net_1\);
    
    \RECD_SER_WORD_RNO[0]\ : MX2
      port map(A => N_33, B => N_34, S => BIT_OS_SEL_0_0, Y => 
        \N_RECD_SER_WORD[0]\);
    
    \Q[6]\ : DFN1C0
      port map(D => \ADJ_Q[6]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[6]_net_1\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \ARB_WRD_40M_FIXED[8]\ : DFN1C0
      port map(D => \Q[8]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[8]_net_1\);
    
    \ARB_BYTE[11]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[11]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[11]_net_1\);
    
    \Q[9]\ : DFN1C0
      port map(D => \ADJ_Q[9]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[9]_net_1\);
    
    \Q[14]\ : DFN1C0
      port map(D => \ADJ_Q[14]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[14]_net_1\);
    
    ADJ_SER_IN_R_0DEL : DFN1C0
      port map(D => ELK_IN_R, CLK => CCC_160M_ADJ, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_R_0DEL\);
    
    \Q[13]\ : DFN1C0
      port map(D => \ADJ_Q[13]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[13]_net_1\);
    
    \ARB_BYTE[9]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[9]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[9]_net_1\);
    
    ADJ_SER_IN_R_1DEL : DFN1C0
      port map(D => \ADJ_SER_IN_R_0DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_SER_IN_R_1DEL\);
    
    \ARB_BYTE[10]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[10]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[10]_net_1\);
    
    \ARB_BYTE_RNIT97T1[10]\ : MX2
      port map(A => N_21, B => N_23, S => BIT_OS_SEL_5(1), Y => 
        N_37);
    
    \ADJ_Q[9]\ : DFN1C0
      port map(D => \ADJ_Q[7]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[9]_net_1\);
    
    \RECD_SER_WORD[7]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[7]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_10(7));
    
    \ARB_WRD_40M_FIXED[5]\ : DFN1C0
      port map(D => \Q[5]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[5]_net_1\);
    
    \ARB_WRD_40M_FIXED[12]\ : DFN1C0
      port map(D => \Q[12]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[12]_net_1\);
    
    \ARB_WRD_40M_FIXED[11]\ : DFN1C0
      port map(D => \Q[11]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[11]_net_1\);
    
    \ARB_WRD_40M_FIXED[0]\ : DFN1C0
      port map(D => \Q[0]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[0]_net_1\);
    
    \ADJ_Q[10]\ : DFN1C0
      port map(D => \ADJ_Q[8]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[10]_net_1\);
    
    \Q[2]\ : DFN1C0
      port map(D => \ADJ_Q[2]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[2]_net_1\);
    
    \ADJ_Q[1]\ : DFN1C0
      port map(D => \ADJ_SER_IN_F_1DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[1]_net_1\);
    
    \RECD_SER_WORD[6]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[6]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_10(6));
    
    \ARB_BYTE_RNIH7CN1[13]\ : MX2
      port map(A => N_24, B => N_32, S => BIT_OS_SEL_5(1), Y => 
        N_40);
    
    \RECD_SER_WORD[2]\ : DFN1C0
      port map(D => \N_RECD_SER_WORD[2]\, CLK => CLK_40M_GL, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => ELK_RX_SER_WORD_10(2));
    
    \ADJ_Q[13]\ : DFN1C0
      port map(D => \ADJ_Q[11]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[13]_net_1\);
    
    \Q[8]\ : DFN1C0
      port map(D => \ADJ_Q[8]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[8]_net_1\);
    
    \ARB_BYTE[5]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[5]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[5]_net_1\);
    
    \ADJ_Q[14]\ : DFN1C0
      port map(D => \ADJ_Q[12]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[14]_net_1\);
    
    \RECD_SER_WORD_RNO[4]\ : MX2
      port map(A => N_37, B => N_38, S => BIT_OS_SEL_0_0, Y => 
        \N_RECD_SER_WORD[4]\);
    
    \Q[12]\ : DFN1C0
      port map(D => \ADJ_Q[12]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[12]_net_1\);
    
    \ARB_BYTE_RNID3CN1[10]\ : MX2
      port map(A => N_23, B => N_31, S => BIT_OS_SEL_5(1), Y => 
        N_39);
    
    \ARB_BYTE[13]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[13]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[13]_net_1\);
    
    \ARB_WRD_40M_FIXED[3]\ : DFN1C0
      port map(D => \Q[3]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[3]_net_1\);
    
    \ARB_BYTE[7]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[7]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[7]_net_1\);
    
    \RECD_SER_WORD_RNO_0[0]\ : MX2
      port map(A => N_17, B => N_19, S => BIT_OS_SEL_5(1), Y => 
        N_33);
    
    \ARB_BYTE_RNIAF542[1]\ : MX2
      port map(A => N_18, B => N_20, S => BIT_OS_SEL_5(1), Y => 
        N_34);
    
    \Q[4]\ : DFN1C0
      port map(D => \ADJ_Q[4]_net_1\, CLK => CCC_160M_FXD, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \Q[4]_net_1\);
    
    \ARB_WRD_40M_FIXED[7]\ : DFN1C0
      port map(D => \Q[7]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => \ARB_WRD_40M_FIXED[7]_net_1\);
    
    \RECD_SER_WORD_RNO[6]\ : MX2
      port map(A => N_39, B => N_40, S => BIT_OS_SEL_0_0, Y => 
        \N_RECD_SER_WORD[6]\);
    
    \ARB_BYTE[3]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[3]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[3]_net_1\);
    
    \ADJ_Q[5]\ : DFN1C0
      port map(D => \ADJ_Q[3]_net_1\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[5]_net_1\);
    
    \ARB_BYTE_RNIHSCQ[12]\ : MX2
      port map(A => \ARB_BYTE[8]_net_1\, B => 
        \ARB_BYTE[12]_net_1\, S => BIT_OS_SEL_6_0, Y => N_31);
    
    \ARB_BYTE[1]\ : DFN1C0
      port map(D => \ARB_WRD_40M_FIXED[1]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_BYTE[1]_net_1\);
    
    \ARB_WRD_40M_FIXED[13]\ : DFN1C0
      port map(D => \Q[13]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[13]_net_1\);
    
    \ADJ_Q[0]\ : DFN1C0
      port map(D => \ADJ_SER_IN_R_1DEL\, CLK => CCC_160M_ADJ, CLR
         => MASTER_DCB_POR_B_i_0_i, Q => \ADJ_Q[0]_net_1\);
    
    \ARB_WRD_40M_FIXED[10]\ : DFN1C0
      port map(D => \Q[10]_net_1\, CLK => CLK_40M_GL, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \ARB_WRD_40M_FIXED[10]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SER320M_3_34_10 is

    port( ELK_TX_DAT                 : in    std_logic_vector(7 downto 0);
          MASTER_SALT_POR_B_i_0_i_3  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_6  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_11 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_1  : in    std_logic;
          ELK_OUT_R                  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_8  : in    std_logic;
          ELK_OUT_F                  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_5  : in    std_logic;
          CCC_160M_FXD               : in    std_logic;
          CLK_40M_GL                 : in    std_logic
        );

end SER320M_3_34_10;

architecture DEF_ARCH of SER320M_3_34_10 is 

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \N_SER_CMD_WORD_R[0]\, \START_RISE\, 
        \N_SER_CMD_WORD_F[0]\, \N_SER_CMD_WORD_R[3]\, 
        \SER_CMD_WORD_R[2]_net_1\, \N_SER_CMD_WORD_R[2]\, 
        \SER_CMD_WORD_R[1]_net_1\, \N_SER_CMD_WORD_R[1]\, 
        \SER_CMD_WORD_R[0]_net_1\, \N_SER_CMD_WORD_F[3]\, 
        \SER_CMD_WORD_F[2]_net_1\, \N_SER_CMD_WORD_F[2]\, 
        \SER_CMD_WORD_F[1]_net_1\, \N_SER_CMD_WORD_F[1]\, 
        \SER_CMD_WORD_F[0]_net_1\, N_START_RISE, 
        \CLK40M_GEN_DEL0\, \SER_OUT_FI\, \SER_OUT_RI\, 
        \SER_CMD_WORD_F[3]_net_1\, \SER_CMD_WORD_R[3]_net_1\, 
        \GND\, \VCC\ : std_logic;

begin 


    SER_OUT_FI : DFN1C0
      port map(D => \SER_CMD_WORD_F[3]_net_1\, CLK => 
        CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_11, Q => 
        \SER_OUT_FI\);
    
    \SER_CMD_WORD_F[3]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[3]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_6, Q => 
        \SER_CMD_WORD_F[3]_net_1\);
    
    \SER_CMD_WORD_R[1]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[1]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_3, Q => 
        \SER_CMD_WORD_R[1]_net_1\);
    
    \SER_CMD_WORD_R[2]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[2]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_3, Q => 
        \SER_CMD_WORD_R[2]_net_1\);
    
    \SER_CMD_WORD_R_RNO[3]\ : MX2
      port map(A => \SER_CMD_WORD_R[2]_net_1\, B => ELK_TX_DAT(7), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_R[3]\);
    
    \SER_CMD_WORD_R_RNO[0]\ : NOR2B
      port map(A => \START_RISE\, B => ELK_TX_DAT(1), Y => 
        \N_SER_CMD_WORD_R[0]\);
    
    \SER_CMD_WORD_F[0]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[0]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_6, Q => 
        \SER_CMD_WORD_F[0]_net_1\);
    
    \SER_CMD_WORD_R_RNO[1]\ : MX2
      port map(A => \SER_CMD_WORD_R[0]_net_1\, B => ELK_TX_DAT(3), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_R[1]\);
    
    \SER_CMD_WORD_F_RNO[2]\ : MX2
      port map(A => \SER_CMD_WORD_F[1]_net_1\, B => ELK_TX_DAT(4), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_F[2]\);
    
    \SER_CMD_WORD_F_RNO[3]\ : MX2
      port map(A => \SER_CMD_WORD_F[2]_net_1\, B => ELK_TX_DAT(6), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_F[3]\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    CLK40M_GEN_DEL0 : DFN1C0
      port map(D => CLK_40M_GL, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_5, Q => \CLK40M_GEN_DEL0\);
    
    SER_OUT_RI : DFN1C0
      port map(D => \SER_CMD_WORD_R[3]_net_1\, CLK => 
        CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_11, Q => 
        \SER_OUT_RI\);
    
    \SER_CMD_WORD_F[2]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[2]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_6, Q => 
        \SER_CMD_WORD_F[2]_net_1\);
    
    \SER_CMD_WORD_F_RNO[1]\ : MX2
      port map(A => \SER_CMD_WORD_F[0]_net_1\, B => ELK_TX_DAT(2), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_F[1]\);
    
    \SER_CMD_WORD_R[0]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[0]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_3, Q => 
        \SER_CMD_WORD_R[0]_net_1\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    START_RISE : DFN1C0
      port map(D => N_START_RISE, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_1, Q => \START_RISE\);
    
    \SER_CMD_WORD_R[3]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_R[3]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_3, Q => 
        \SER_CMD_WORD_R[3]_net_1\);
    
    \SER_CMD_WORD_F_RNO[0]\ : NOR2B
      port map(A => \START_RISE\, B => ELK_TX_DAT(0), Y => 
        \N_SER_CMD_WORD_F[0]\);
    
    SER_OUT_RDEL : DFN1C0
      port map(D => \SER_OUT_RI\, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_5, Q => ELK_OUT_R);
    
    \SER_CMD_WORD_F[1]\ : DFN1C0
      port map(D => \N_SER_CMD_WORD_F[1]\, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_6, Q => 
        \SER_CMD_WORD_F[1]_net_1\);
    
    START_RISE_RNO : NOR2B
      port map(A => \CLK40M_GEN_DEL0\, B => CLK_40M_GL, Y => 
        N_START_RISE);
    
    \SER_CMD_WORD_R_RNO[2]\ : MX2
      port map(A => \SER_CMD_WORD_R[1]_net_1\, B => ELK_TX_DAT(5), 
        S => \START_RISE\, Y => \N_SER_CMD_WORD_R[2]\);
    
    SER_OUT_FDEL : DFN1C0
      port map(D => \SER_OUT_FI\, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_8, Q => ELK_OUT_F);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity DDR_BIDIR_LVDS_DUAL_CLK_10 is

    port( DCB_SALT_SEL_c_i : in    std_logic;
          ELK10_DAT_P      : inout std_logic := 'Z';
          ELK10_DAT_N      : inout std_logic := 'Z';
          ELK_OUT_R        : in    std_logic;
          ELK_OUT_F        : in    std_logic;
          CCC_160M_FXD     : in    std_logic;
          CCC_160M_ADJ     : in    std_logic;
          ELK_IN_DDR_R     : out   std_logic;
          ELK_IN_DDR_F     : out   std_logic
        );

end DDR_BIDIR_LVDS_DUAL_CLK_10;

architecture DEF_ARCH of DDR_BIDIR_LVDS_DUAL_CLK_10 is 

  component DDR_REG
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          QR  : out   std_logic;
          QF  : out   std_logic
        );
  end component;

  component DDR_OUT
    port( DR  : in    std_logic := 'U';
          DF  : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component BIBUF_LVDS
    port( PADP : inout   std_logic;
          PADN : inout   std_logic;
          D    : in    std_logic := 'U';
          E    : in    std_logic := 'U';
          Y    : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal DDR_BIDIR_LVDS_DUAL_CLK_10_GND, BIBUF_LVDS_0_Y, 
        DDR_OUT_0_Q, \VCC\ : std_logic;

begin 


    DDR_REG_0 : DDR_REG
      port map(D => BIBUF_LVDS_0_Y, CLK => CCC_160M_ADJ, CLR => 
        DDR_BIDIR_LVDS_DUAL_CLK_10_GND, QR => ELK_IN_DDR_R, QF
         => ELK_IN_DDR_F);
    
    DDR_OUT_0 : DDR_OUT
      port map(DR => ELK_OUT_R, DF => ELK_OUT_F, CLK => 
        CCC_160M_FXD, CLR => DDR_BIDIR_LVDS_DUAL_CLK_10_GND, Q
         => DDR_OUT_0_Q);
    
    BIBUF_LVDS_0 : BIBUF_LVDS
      port map(PADP => ELK10_DAT_P, PADN => ELK10_DAT_N, D => 
        DDR_OUT_0_Q, E => DCB_SALT_SEL_c_i, Y => BIBUF_LVDS_0_Y);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    GND_i : GND
      port map(Y => DDR_BIDIR_LVDS_DUAL_CLK_10_GND);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity SYNC_DAT_SEL_10 is

    port( ELK_TX_DAT                 : out   std_logic_vector(7 downto 0);
          PATT_ELK_DAT_10            : in    std_logic_vector(7 downto 0);
          OP_MODE_c_3_0              : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_17 : in    std_logic;
          CLK_40M_GL                 : in    std_logic
        );

end SYNC_DAT_SEL_10;

architecture DEF_ARCH of SYNC_DAT_SEL_10 is 

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \N_SERDAT[0]\, \N_SERDAT[1]\, \N_SERDAT[2]\, 
        \N_SERDAT[3]\, \N_SERDAT[4]\, \N_SERDAT[5]\, 
        \N_SERDAT[6]\, \N_SERDAT[7]\, \GND\, \VCC\ : std_logic;

begin 


    \SERDAT_RNO[4]\ : NOR2A
      port map(A => PATT_ELK_DAT_10(4), B => OP_MODE_c_3_0, Y => 
        \N_SERDAT[4]\);
    
    \SERDAT_RNO[0]\ : NOR2A
      port map(A => PATT_ELK_DAT_10(0), B => OP_MODE_c_3_0, Y => 
        \N_SERDAT[0]\);
    
    \SERDAT[6]\ : DFN1C0
      port map(D => \N_SERDAT[6]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_17, Q => ELK_TX_DAT(6));
    
    \SERDAT[4]\ : DFN1C0
      port map(D => \N_SERDAT[4]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_17, Q => ELK_TX_DAT(4));
    
    \SERDAT_RNO[7]\ : OR2
      port map(A => PATT_ELK_DAT_10(7), B => OP_MODE_c_3_0, Y => 
        \N_SERDAT[7]\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \SERDAT_RNO[3]\ : OR2
      port map(A => PATT_ELK_DAT_10(3), B => OP_MODE_c_3_0, Y => 
        \N_SERDAT[3]\);
    
    \SERDAT_RNO[2]\ : OR2
      port map(A => PATT_ELK_DAT_10(2), B => OP_MODE_c_3_0, Y => 
        \N_SERDAT[2]\);
    
    \SERDAT[5]\ : DFN1C0
      port map(D => \N_SERDAT[5]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_17, Q => ELK_TX_DAT(5));
    
    \SERDAT[7]\ : DFN1C0
      port map(D => \N_SERDAT[7]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_17, Q => ELK_TX_DAT(7));
    
    GND_i : GND
      port map(Y => \GND\);
    
    \SERDAT_RNO[5]\ : NOR2A
      port map(A => PATT_ELK_DAT_10(5), B => OP_MODE_c_3_0, Y => 
        \N_SERDAT[5]\);
    
    \SERDAT[0]\ : DFN1C0
      port map(D => \N_SERDAT[0]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_17, Q => ELK_TX_DAT(0));
    
    \SERDAT_RNO[6]\ : NOR2A
      port map(A => PATT_ELK_DAT_10(6), B => OP_MODE_c_3_0, Y => 
        \N_SERDAT[6]\);
    
    \SERDAT[1]\ : DFN1C0
      port map(D => \N_SERDAT[1]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_17, Q => ELK_TX_DAT(1));
    
    \SERDAT_RNO[1]\ : OR2
      port map(A => PATT_ELK_DAT_10(1), B => OP_MODE_c_3_0, Y => 
        \N_SERDAT[1]\);
    
    \SERDAT[3]\ : DFN1C0
      port map(D => \N_SERDAT[3]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_17, Q => ELK_TX_DAT(3));
    
    \SERDAT[2]\ : DFN1C0
      port map(D => \N_SERDAT[2]\, CLK => CLK_40M_GL, CLR => 
        MASTER_SALT_POR_B_i_0_i_17, Q => ELK_TX_DAT(2));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity ELINK_SLAVE_15_5 is

    port( BIT_OS_SEL_6_0             : in    std_logic;
          BIT_OS_SEL_5               : in    std_logic_vector(2 downto 1);
          BIT_OS_SEL_7_0             : in    std_logic;
          BIT_OS_SEL_0_d0            : in    std_logic;
          BIT_OS_SEL_0_0             : in    std_logic;
          ELK_RX_SER_WORD_10         : out   std_logic_vector(7 downto 0);
          OP_MODE_c_3_0              : in    std_logic;
          PATT_ELK_DAT_10            : in    std_logic_vector(7 downto 0);
          MASTER_DCB_POR_B_i_0_i     : in    std_logic;
          ELK10_DAT_N                : inout std_logic := 'Z';
          ELK10_DAT_P                : inout std_logic := 'Z';
          DCB_SALT_SEL_c_i           : in    std_logic;
          CCC_160M_FXD               : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_5  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_8  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_1  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_11 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_6  : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_3  : in    std_logic;
          CLK_40M_GL                 : in    std_logic;
          MASTER_SALT_POR_B_i_0_i_17 : in    std_logic;
          DEV_RST_B_c_0              : in    std_logic;
          CCC_160M_ADJ               : in    std_logic
        );

end ELINK_SLAVE_15_5;

architecture DEF_ARCH of ELINK_SLAVE_15_5 is 

  component SLAVE_DES320S_1_17_8
    port( ELK_RX_SER_WORD_10     : out   std_logic_vector(7 downto 0);
          BIT_OS_SEL_0_0         : in    std_logic := 'U';
          BIT_OS_SEL_0_d0        : in    std_logic := 'U';
          BIT_OS_SEL_7_0         : in    std_logic := 'U';
          BIT_OS_SEL_5           : in    std_logic_vector(2 downto 1) := (others => 'U');
          BIT_OS_SEL_6_0         : in    std_logic := 'U';
          CLK_40M_GL             : in    std_logic := 'U';
          CCC_160M_FXD           : in    std_logic := 'U';
          ELK_IN_R               : in    std_logic := 'U';
          ELK_IN_F               : in    std_logic := 'U';
          MASTER_DCB_POR_B_i_0_i : in    std_logic := 'U';
          CCC_160M_ADJ           : in    std_logic := 'U'
        );
  end component;

  component SER320M_3_34_10
    port( ELK_TX_DAT                 : in    std_logic_vector(7 downto 0) := (others => 'U');
          MASTER_SALT_POR_B_i_0_i_3  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_6  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_11 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_1  : in    std_logic := 'U';
          ELK_OUT_R                  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_8  : in    std_logic := 'U';
          ELK_OUT_F                  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_5  : in    std_logic := 'U';
          CCC_160M_FXD               : in    std_logic := 'U';
          CLK_40M_GL                 : in    std_logic := 'U'
        );
  end component;

  component DDR_BIDIR_LVDS_DUAL_CLK_10
    port( DCB_SALT_SEL_c_i : in    std_logic := 'U';
          ELK10_DAT_P      : inout   std_logic;
          ELK10_DAT_N      : inout   std_logic;
          ELK_OUT_R        : in    std_logic := 'U';
          ELK_OUT_F        : in    std_logic := 'U';
          CCC_160M_FXD     : in    std_logic := 'U';
          CCC_160M_ADJ     : in    std_logic := 'U';
          ELK_IN_DDR_R     : out   std_logic;
          ELK_IN_DDR_F     : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component SYNC_DAT_SEL_10
    port( ELK_TX_DAT                 : out   std_logic_vector(7 downto 0);
          PATT_ELK_DAT_10            : in    std_logic_vector(7 downto 0) := (others => 'U');
          OP_MODE_c_3_0              : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_17 : in    std_logic := 'U';
          CLK_40M_GL                 : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \ELK_IN_F\, ELK_IN_DDR_F, \ELK_IN_R\, ELK_IN_DDR_R, 
        \ELK_TX_DAT[0]\, \ELK_TX_DAT[1]\, \ELK_TX_DAT[2]\, 
        \ELK_TX_DAT[3]\, \ELK_TX_DAT[4]\, \ELK_TX_DAT[5]\, 
        \ELK_TX_DAT[6]\, \ELK_TX_DAT[7]\, ELK_OUT_R, ELK_OUT_F, 
        \GND\, \VCC\ : std_logic;

    for all : SLAVE_DES320S_1_17_8
	Use entity work.SLAVE_DES320S_1_17_8(DEF_ARCH);
    for all : SER320M_3_34_10
	Use entity work.SER320M_3_34_10(DEF_ARCH);
    for all : DDR_BIDIR_LVDS_DUAL_CLK_10
	Use entity work.DDR_BIDIR_LVDS_DUAL_CLK_10(DEF_ARCH);
    for all : SYNC_DAT_SEL_10
	Use entity work.SYNC_DAT_SEL_10(DEF_ARCH);
begin 


    U_SLAVE_1ELK : SLAVE_DES320S_1_17_8
      port map(ELK_RX_SER_WORD_10(7) => ELK_RX_SER_WORD_10(7), 
        ELK_RX_SER_WORD_10(6) => ELK_RX_SER_WORD_10(6), 
        ELK_RX_SER_WORD_10(5) => ELK_RX_SER_WORD_10(5), 
        ELK_RX_SER_WORD_10(4) => ELK_RX_SER_WORD_10(4), 
        ELK_RX_SER_WORD_10(3) => ELK_RX_SER_WORD_10(3), 
        ELK_RX_SER_WORD_10(2) => ELK_RX_SER_WORD_10(2), 
        ELK_RX_SER_WORD_10(1) => ELK_RX_SER_WORD_10(1), 
        ELK_RX_SER_WORD_10(0) => ELK_RX_SER_WORD_10(0), 
        BIT_OS_SEL_0_0 => BIT_OS_SEL_0_0, BIT_OS_SEL_0_d0 => 
        BIT_OS_SEL_0_d0, BIT_OS_SEL_7_0 => BIT_OS_SEL_7_0, 
        BIT_OS_SEL_5(2) => BIT_OS_SEL_5(2), BIT_OS_SEL_5(1) => 
        BIT_OS_SEL_5(1), BIT_OS_SEL_6_0 => BIT_OS_SEL_6_0, 
        CLK_40M_GL => CLK_40M_GL, CCC_160M_FXD => CCC_160M_FXD, 
        ELK_IN_R => \ELK_IN_R\, ELK_IN_F => \ELK_IN_F\, 
        MASTER_DCB_POR_B_i_0_i => MASTER_DCB_POR_B_i_0_i, 
        CCC_160M_ADJ => CCC_160M_ADJ);
    
    U_ELK1_CMD_TX : SER320M_3_34_10
      port map(ELK_TX_DAT(7) => \ELK_TX_DAT[7]\, ELK_TX_DAT(6)
         => \ELK_TX_DAT[6]\, ELK_TX_DAT(5) => \ELK_TX_DAT[5]\, 
        ELK_TX_DAT(4) => \ELK_TX_DAT[4]\, ELK_TX_DAT(3) => 
        \ELK_TX_DAT[3]\, ELK_TX_DAT(2) => \ELK_TX_DAT[2]\, 
        ELK_TX_DAT(1) => \ELK_TX_DAT[1]\, ELK_TX_DAT(0) => 
        \ELK_TX_DAT[0]\, MASTER_SALT_POR_B_i_0_i_3 => 
        MASTER_SALT_POR_B_i_0_i_3, MASTER_SALT_POR_B_i_0_i_6 => 
        MASTER_SALT_POR_B_i_0_i_6, MASTER_SALT_POR_B_i_0_i_11 => 
        MASTER_SALT_POR_B_i_0_i_11, MASTER_SALT_POR_B_i_0_i_1 => 
        MASTER_SALT_POR_B_i_0_i_1, ELK_OUT_R => ELK_OUT_R, 
        MASTER_SALT_POR_B_i_0_i_8 => MASTER_SALT_POR_B_i_0_i_8, 
        ELK_OUT_F => ELK_OUT_F, MASTER_SALT_POR_B_i_0_i_5 => 
        MASTER_SALT_POR_B_i_0_i_5, CCC_160M_FXD => CCC_160M_FXD, 
        CLK_40M_GL => CLK_40M_GL);
    
    U_DDR_ELK1 : DDR_BIDIR_LVDS_DUAL_CLK_10
      port map(DCB_SALT_SEL_c_i => DCB_SALT_SEL_c_i, ELK10_DAT_P
         => ELK10_DAT_P, ELK10_DAT_N => ELK10_DAT_N, ELK_OUT_R
         => ELK_OUT_R, ELK_OUT_F => ELK_OUT_F, CCC_160M_FXD => 
        CCC_160M_FXD, CCC_160M_ADJ => CCC_160M_ADJ, ELK_IN_DDR_R
         => ELK_IN_DDR_R, ELK_IN_DDR_F => ELK_IN_DDR_F);
    
    ELK_IN_F : DFN1C0
      port map(D => ELK_IN_DDR_F, CLK => CCC_160M_ADJ, CLR => 
        DEV_RST_B_c_0, Q => \ELK_IN_F\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    U_ELK1_SERDAT_SOURCE : SYNC_DAT_SEL_10
      port map(ELK_TX_DAT(7) => \ELK_TX_DAT[7]\, ELK_TX_DAT(6)
         => \ELK_TX_DAT[6]\, ELK_TX_DAT(5) => \ELK_TX_DAT[5]\, 
        ELK_TX_DAT(4) => \ELK_TX_DAT[4]\, ELK_TX_DAT(3) => 
        \ELK_TX_DAT[3]\, ELK_TX_DAT(2) => \ELK_TX_DAT[2]\, 
        ELK_TX_DAT(1) => \ELK_TX_DAT[1]\, ELK_TX_DAT(0) => 
        \ELK_TX_DAT[0]\, PATT_ELK_DAT_10(7) => PATT_ELK_DAT_10(7), 
        PATT_ELK_DAT_10(6) => PATT_ELK_DAT_10(6), 
        PATT_ELK_DAT_10(5) => PATT_ELK_DAT_10(5), 
        PATT_ELK_DAT_10(4) => PATT_ELK_DAT_10(4), 
        PATT_ELK_DAT_10(3) => PATT_ELK_DAT_10(3), 
        PATT_ELK_DAT_10(2) => PATT_ELK_DAT_10(2), 
        PATT_ELK_DAT_10(1) => PATT_ELK_DAT_10(1), 
        PATT_ELK_DAT_10(0) => PATT_ELK_DAT_10(0), OP_MODE_c_3_0
         => OP_MODE_c_3_0, MASTER_SALT_POR_B_i_0_i_17 => 
        MASTER_SALT_POR_B_i_0_i_17, CLK_40M_GL => CLK_40M_GL);
    
    ELK_IN_R : DFN1C0
      port map(D => ELK_IN_DDR_R, CLK => CCC_160M_ADJ, CLR => 
        DEV_RST_B_c_0, Q => \ELK_IN_R\);
    
    GND_i : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity TOP_COMET is

    port( CLK200_P        : in    std_logic;
          CLK200_N        : in    std_logic;
          DEV_RST_B       : in    std_logic;
          DCB_SALT_SEL    : in    std_logic;
          EXTCLK_40MHZ    : out   std_logic;
          EXT_INT_REF_SEL : in    std_logic;
          ALL_PLL_LOCK    : out   std_logic;
          P_MASTER_POR_B  : out   std_logic;
          P_USB_MASTER_EN : out   std_logic;
          P_CLK_40M_GL    : out   std_logic;
          P_CCC_160M_FXD  : out   std_logic;
          P_CCC_160M_ADJ  : out   std_logic;
          P_ELK0_SYNC_DET : out   std_logic;
          P_TFC_SYNC_DET  : out   std_logic;
          P_OP_MODE1_SPE  : out   std_logic;
          P_OP_MODE2_TE   : out   std_logic;
          P_OP_MODE5_AAE  : out   std_logic;
          P_OP_MODE6_EE   : out   std_logic;
          BIDIR_CLK40M_P  : inout std_logic := 'Z';
          BIDIR_CLK40M_N  : inout std_logic := 'Z';
          TX_CLK40M_P     : out   std_logic;
          TX_CLK40M_N     : out   std_logic;
          USBCLK60MHZ     : in    std_logic;
          BIDIR_USB_ADBUS : inout std_logic_vector(7 downto 0) := (others => 'Z');
          USB_OE_B        : out   std_logic;
          P_USB_RXF_B     : in    std_logic;
          USB_RD_B        : out   std_logic;
          P_USB_TXE_B     : in    std_logic;
          USB_WR_B        : out   std_logic;
          USB_SIWU_B      : out   std_logic;
          TFC_DAT_0P      : inout std_logic := 'Z';
          TFC_DAT_0N      : inout std_logic := 'Z';
          REF_CLK_0P      : inout std_logic := 'Z';
          REF_CLK_0N      : inout std_logic := 'Z';
          ELK0_DAT_P      : inout std_logic := 'Z';
          ELK0_DAT_N      : inout std_logic := 'Z';
          ELK1_DAT_P      : inout std_logic := 'Z';
          ELK1_DAT_N      : inout std_logic := 'Z';
          ELK2_DAT_P      : inout std_logic := 'Z';
          ELK2_DAT_N      : inout std_logic := 'Z';
          ELK3_DAT_P      : inout std_logic := 'Z';
          ELK3_DAT_N      : inout std_logic := 'Z';
          ELK4_DAT_P      : inout std_logic := 'Z';
          ELK4_DAT_N      : inout std_logic := 'Z';
          ELK5_DAT_P      : inout std_logic := 'Z';
          ELK5_DAT_N      : inout std_logic := 'Z';
          ELK6_DAT_P      : inout std_logic := 'Z';
          ELK6_DAT_N      : inout std_logic := 'Z';
          ELK7_DAT_P      : inout std_logic := 'Z';
          ELK7_DAT_N      : inout std_logic := 'Z';
          ELK8_DAT_P      : inout std_logic := 'Z';
          ELK8_DAT_N      : inout std_logic := 'Z';
          ELK9_DAT_P      : inout std_logic := 'Z';
          ELK9_DAT_N      : inout std_logic := 'Z';
          ELK10_DAT_P     : inout std_logic := 'Z';
          ELK10_DAT_N     : inout std_logic := 'Z';
          ELK11_DAT_P     : inout std_logic := 'Z';
          ELK11_DAT_N     : inout std_logic := 'Z';
          ELK12_DAT_P     : inout std_logic := 'Z';
          ELK12_DAT_N     : inout std_logic := 'Z';
          ELK13_DAT_P     : inout std_logic := 'Z';
          ELK13_DAT_N     : inout std_logic := 'Z';
          ELK14_DAT_P     : inout std_logic := 'Z';
          ELK14_DAT_N     : inout std_logic := 'Z';
          ELK15_DAT_P     : inout std_logic := 'Z';
          ELK15_DAT_N     : inout std_logic := 'Z';
          ELK16_DAT_P     : inout std_logic := 'Z';
          ELK16_DAT_N     : inout std_logic := 'Z';
          ELK17_DAT_P     : inout std_logic := 'Z';
          ELK17_DAT_N     : inout std_logic := 'Z';
          ELK18_DAT_P     : inout std_logic := 'Z';
          ELK18_DAT_N     : inout std_logic := 'Z';
          ELK19_DAT_P     : inout std_logic := 'Z';
          ELK19_DAT_N     : inout std_logic := 'Z'
        );

end TOP_COMET;

architecture DEF_ARCH of TOP_COMET is 

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component INBUF
    port( PAD : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component ELINK_SLAVE_INV_2
    port( BIT_OS_SEL_0_d0            : in    std_logic := 'U';
          BIT_OS_SEL_0_0             : in    std_logic := 'U';
          BIT_OS_SEL_1               : in    std_logic_vector(2 downto 0) := (others => 'U');
          BIT_OS_SEL_2_0             : in    std_logic := 'U';
          ELK_RX_SER_WORD_1          : out   std_logic_vector(7 downto 0);
          OP_MODE_c_5_0              : in    std_logic := 'U';
          PATT_ELK_DAT_1             : in    std_logic_vector(7 downto 0) := (others => 'U');
          MASTER_DCB_POR_B_i_0_i     : in    std_logic := 'U';
          ELK1_DAT_N                 : inout   std_logic;
          ELK1_DAT_P                 : inout   std_logic;
          DCB_SALT_SEL_c_i           : in    std_logic := 'U';
          CCC_160M_FXD               : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_14 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_7  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_1  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_16 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_4  : in    std_logic := 'U';
          CLK_40M_GL                 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_11 : in    std_logic := 'U';
          DEV_RST_B_c_0              : in    std_logic := 'U';
          CCC_160M_ADJ               : in    std_logic := 'U'
        );
  end component;

  component OUTBUF
    port( D   : in    std_logic := 'U';
          PAD : out   std_logic
        );
  end component;

  component ELINK_SLAVE_INV_2_0
    port( BIT_OS_SEL_7_0             : in    std_logic := 'U';
          BIT_OS_SEL_6_0             : in    std_logic := 'U';
          BIT_OS_SEL_0_d0            : in    std_logic := 'U';
          BIT_OS_SEL_0               : in    std_logic_vector(2 downto 1) := (others => 'U');
          BIT_OS_SEL_1_0             : in    std_logic := 'U';
          ELK_RX_SER_WORD_3          : out   std_logic_vector(7 downto 0);
          OP_MODE_c_5_0              : in    std_logic := 'U';
          PATT_ELK_DAT_3             : in    std_logic_vector(7 downto 0) := (others => 'U');
          MASTER_DCB_POR_B_i_0_i     : in    std_logic := 'U';
          ELK3_DAT_N                 : inout   std_logic;
          ELK3_DAT_P                 : inout   std_logic;
          DCB_SALT_SEL_c_i           : in    std_logic := 'U';
          CCC_160M_FXD               : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_8  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_5  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_2  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_3  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_16 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_12 : in    std_logic := 'U';
          CLK_40M_GL                 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_14 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_15 : in    std_logic := 'U';
          DEV_RST_B_c                : in    std_logic := 'U';
          CCC_160M_ADJ               : in    std_logic := 'U'
        );
  end component;

  component USB_INTERFACE
    port( OP_MODE_c_6_0          : out   std_logic;
          OP_MODE_c_5_0          : out   std_logic;
          OP_MODE_c_4_0          : out   std_logic;
          OP_MODE_c_3_0          : out   std_logic;
          OP_MODE_c_2_0          : out   std_logic;
          OP_MODE_c_1_0          : out   std_logic;
          OP_MODE_c_0_0          : out   std_logic;
          OP_MODE_c_1_d0         : out   std_logic;
          OP_MODE_c_5_d0         : out   std_logic;
          OP_MODE_c_4_d0         : out   std_logic;
          OP_MODE_c_0_d0         : out   std_logic;
          OP_MODE_0_0            : out   std_logic;
          OP_MODE_0_4            : out   std_logic;
          ELKS_STOP_ADDR         : out   std_logic_vector(7 downto 0);
          ELKS_STRT_ADDR         : out   std_logic_vector(7 downto 0);
          TFC_STOP_ADDR_0        : out   std_logic_vector(7 downto 0);
          TFC_STRT_ADDR_0        : out   std_logic_vector(7 downto 0);
          BIDIR_USB_ADBUS        : inout   std_logic_vector(7 downto 0);
          PATT_ELK_DAT_19        : out   std_logic_vector(7 downto 0);
          ELK_RX_SER_WORD_19     : in    std_logic_vector(7 downto 0) := (others => 'U');
          PATT_ELK_DAT_18        : out   std_logic_vector(7 downto 0);
          ELK_RX_SER_WORD_18     : in    std_logic_vector(7 downto 0) := (others => 'U');
          PATT_ELK_DAT_17        : out   std_logic_vector(7 downto 0);
          ELK_RX_SER_WORD_17     : in    std_logic_vector(7 downto 0) := (others => 'U');
          PATT_ELK_DAT_16        : out   std_logic_vector(7 downto 0);
          ELK_RX_SER_WORD_16     : in    std_logic_vector(7 downto 0) := (others => 'U');
          PATT_ELK_DAT_15        : out   std_logic_vector(7 downto 0);
          ELK_RX_SER_WORD_15     : in    std_logic_vector(7 downto 0) := (others => 'U');
          PATT_ELK_DAT_14        : out   std_logic_vector(7 downto 0);
          ELK_RX_SER_WORD_14     : in    std_logic_vector(7 downto 0) := (others => 'U');
          PATT_ELK_DAT_13        : out   std_logic_vector(7 downto 0);
          ELK_RX_SER_WORD_13     : in    std_logic_vector(7 downto 0) := (others => 'U');
          PATT_ELK_DAT_12        : out   std_logic_vector(7 downto 0);
          ELK_RX_SER_WORD_12     : in    std_logic_vector(7 downto 0) := (others => 'U');
          PATT_ELK_DAT_11        : out   std_logic_vector(7 downto 0);
          ELK_RX_SER_WORD_11     : in    std_logic_vector(7 downto 0) := (others => 'U');
          PATT_ELK_DAT_10        : out   std_logic_vector(7 downto 0);
          ELK_RX_SER_WORD_10     : in    std_logic_vector(7 downto 0) := (others => 'U');
          PATT_ELK_DAT_9         : out   std_logic_vector(7 downto 0);
          ELK_RX_SER_WORD_9      : in    std_logic_vector(7 downto 0) := (others => 'U');
          PATT_ELK_DAT_8         : out   std_logic_vector(7 downto 0);
          ELK_RX_SER_WORD_8      : in    std_logic_vector(7 downto 0) := (others => 'U');
          PATT_ELK_DAT_7         : out   std_logic_vector(7 downto 0);
          ELK_RX_SER_WORD_7      : in    std_logic_vector(7 downto 0) := (others => 'U');
          PATT_ELK_DAT_6         : out   std_logic_vector(7 downto 0);
          ELK_RX_SER_WORD_6      : in    std_logic_vector(7 downto 0) := (others => 'U');
          PATT_ELK_DAT_5         : out   std_logic_vector(7 downto 0);
          ELK_RX_SER_WORD_5      : in    std_logic_vector(7 downto 0) := (others => 'U');
          PATT_ELK_DAT_4         : out   std_logic_vector(7 downto 0);
          ELK_RX_SER_WORD_4      : in    std_logic_vector(7 downto 0) := (others => 'U');
          PATT_ELK_DAT_3         : out   std_logic_vector(7 downto 0);
          ELK_RX_SER_WORD_3      : in    std_logic_vector(7 downto 0) := (others => 'U');
          PATT_ELK_DAT_2         : out   std_logic_vector(7 downto 0);
          ELK_RX_SER_WORD_2      : in    std_logic_vector(7 downto 0) := (others => 'U');
          PATT_ELK_DAT_1         : out   std_logic_vector(7 downto 0);
          ELKS_ADDRB_0_0         : in    std_logic := 'U';
          ELKS_ADDRB_0_2         : in    std_logic := 'U';
          ELKS_ADDRB_0_4         : in    std_logic := 'U';
          ELK_RX_SER_WORD_1      : in    std_logic_vector(7 downto 0) := (others => 'U');
          PATT_ELK_DAT_0         : out   std_logic_vector(7 downto 0);
          ELKS_ADDRB             : in    std_logic_vector(7 downto 0) := (others => 'U');
          ELK_RX_SER_WORD_0      : in    std_logic_vector(7 downto 0) := (others => 'U');
          PATT_TFC_DAT           : out   std_logic_vector(7 downto 0);
          TFC_ADDRB              : in    std_logic_vector(7 downto 0) := (others => 'U');
          TFC_RX_SER_WORD        : in    std_logic_vector(7 downto 0) := (others => 'U');
          P_MASTER_POR_B_c_0_0   : in    std_logic := 'U';
          P_MASTER_POR_B_c_1     : in    std_logic := 'U';
          P_MASTER_POR_B_c       : in    std_logic := 'U';
          P_MASTER_POR_B_c_6     : in    std_logic := 'U';
          P_MASTER_POR_B_c_24    : in    std_logic := 'U';
          P_MASTER_POR_B_c_3     : in    std_logic := 'U';
          P_MASTER_POR_B_c_26    : in    std_logic := 'U';
          P_MASTER_POR_B_c_33    : in    std_logic := 'U';
          P_MASTER_POR_B_c_22_0  : in    std_logic := 'U';
          P_MASTER_POR_B_c_28    : in    std_logic := 'U';
          P_MASTER_POR_B_c_23    : in    std_logic := 'U';
          P_MASTER_POR_B_c_19    : in    std_logic := 'U';
          P_MASTER_POR_B_c_24_0  : in    std_logic := 'U';
          P_MASTER_POR_B_c_25    : in    std_logic := 'U';
          P_MASTER_POR_B_c_29    : in    std_logic := 'U';
          P_MASTER_POR_B_c_30    : in    std_logic := 'U';
          P_MASTER_POR_B_c_27    : in    std_logic := 'U';
          P_MASTER_POR_B_c_17    : in    std_logic := 'U';
          P_MASTER_POR_B_c_32    : in    std_logic := 'U';
          P_MASTER_POR_B_c_32_0  : in    std_logic := 'U';
          P_MASTER_POR_B_c_21    : in    std_logic := 'U';
          P_MASTER_POR_B_c_22    : in    std_logic := 'U';
          ELKS_RAM_BLKB_EN       : in    std_logic := 'U';
          ELKS_RWB               : in    std_logic := 'U';
          TFC_RAM_BLKB_EN        : in    std_logic := 'U';
          CLK_40M_GL             : in    std_logic := 'U';
          TFC_RWB                : in    std_logic := 'U';
          P_USB_MASTER_EN_c_1    : in    std_logic := 'U';
          P_USB_MASTER_EN_c_0    : in    std_logic := 'U';
          P_USB_MASTER_EN_c_2    : in    std_logic := 'U';
          P_USB_MASTER_EN_c_20   : in    std_logic := 'U';
          P_USB_MASTER_EN_c_6    : in    std_logic := 'U';
          P_USB_MASTER_EN_c_9    : in    std_logic := 'U';
          P_USB_MASTER_EN_c_11   : in    std_logic := 'U';
          P_USB_MASTER_EN_c_12   : in    std_logic := 'U';
          P_USB_MASTER_EN_c_14   : in    std_logic := 'U';
          P_USB_MASTER_EN_c_18   : in    std_logic := 'U';
          P_USB_MASTER_EN_c_7    : in    std_logic := 'U';
          P_USB_MASTER_EN_c_21   : in    std_logic := 'U';
          P_USB_MASTER_EN_c_17   : in    std_logic := 'U';
          P_USB_MASTER_EN_c_15   : in    std_logic := 'U';
          P_USB_MASTER_EN_c_4    : in    std_logic := 'U';
          USB_WR_BI              : out   std_logic;
          P_USB_MASTER_EN_c_3    : in    std_logic := 'U';
          P_USB_MASTER_EN_c_8    : in    std_logic := 'U';
          USB_SIWU_BI            : out   std_logic;
          P_USB_MASTER_EN_c_19   : in    std_logic := 'U';
          USB_OE_BI              : out   std_logic;
          USB_RD_BI              : out   std_logic;
          P_USB_MASTER_EN_c_13   : in    std_logic := 'U';
          P_USB_MASTER_EN_c_5    : in    std_logic := 'U';
          P_USB_MASTER_EN_c_10   : in    std_logic := 'U';
          P_USB_MASTER_EN_c_22   : in    std_logic := 'U';
          P_USB_TXE_B_c          : in    std_logic := 'U';
          P_USB_MASTER_EN_c_16   : in    std_logic := 'U';
          P_USB_MASTER_EN_c_22_0 : in    std_logic := 'U';
          P_USB_MASTER_EN_c_2_0  : in    std_logic := 'U';
          P_USB_MASTER_EN_c_1_0  : in    std_logic := 'U';
          P_USB_MASTER_EN_c      : in    std_logic := 'U';
          P_USB_RXF_B_c          : in    std_logic := 'U';
          CLK60MHZ               : in    std_logic := 'U'
        );
  end component;

  component SYNC_DAT_SEL
    port( TFC_TX_DAT             : out   std_logic_vector(7 downto 0);
          PATT_TFC_DAT           : in    std_logic_vector(7 downto 0) := (others => 'U');
          OP_MODE_c_0_0          : in    std_logic := 'U';
          MASTER_DCB_POR_B_i_0_i : in    std_logic := 'U';
          CLK_40M_GL             : in    std_logic := 'U'
        );
  end component;

  component CLK_FXD_40_160_A60M
    port( USBCLK60MHZ_c    : in    std_logic := 'U';
          CCC_MAIN_LOCK    : out   std_logic;
          CLK60MHZ_1       : out   std_logic;
          CCC_160M_FXD_1   : out   std_logic;
          CLK_40M_GL_1     : out   std_logic;
          CLK_40M_BUF_RECD : in    std_logic := 'U'
        );
  end component;

  component ELINK_SLAVE_15_13
    port( BIT_OS_SEL_0               : in    std_logic_vector(2 downto 1) := (others => 'U');
          BIT_OS_SEL_1               : in    std_logic_vector(2 downto 1) := (others => 'U');
          BIT_OS_SEL_2               : in    std_logic_vector(1 downto 0) := (others => 'U');
          ELK_RX_SER_WORD_18         : out   std_logic_vector(7 downto 0);
          OP_MODE_c_1_0              : in    std_logic := 'U';
          OP_MODE_c_2_0              : in    std_logic := 'U';
          PATT_ELK_DAT_18            : in    std_logic_vector(7 downto 0) := (others => 'U');
          MASTER_DCB_POR_B_i_0_i     : in    std_logic := 'U';
          ELK18_DAT_N                : inout   std_logic;
          ELK18_DAT_P                : inout   std_logic;
          DCB_SALT_SEL_c_i           : in    std_logic := 'U';
          CCC_160M_FXD               : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_9  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_4  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_1  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_17 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_3  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_0  : in    std_logic := 'U';
          CLK_40M_GL                 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_13 : in    std_logic := 'U';
          DEV_RST_B_c_0              : in    std_logic := 'U';
          CCC_160M_ADJ               : in    std_logic := 'U'
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component tristate_buf_1
    port( P_USB_MASTER_EN_c : in    std_logic := 'U';
          USB_OE_BI         : in    std_logic := 'U';
          USB_OE_B          : out   std_logic
        );
  end component;

  component BIDIR_LVDS_IO_0
    port( DCB_SALT_SEL_c : in    std_logic := 'U';
          CLK_40M_GL     : in    std_logic := 'U';
          EXTCLK_40MHZ_c : out   std_logic;
          REF_CLK_0P     : inout   std_logic;
          REF_CLK_0N     : inout   std_logic
        );
  end component;

  component ELINK_SLAVE_15_6
    port( BIT_OS_SEL_4               : in    std_logic_vector(2 downto 1) := (others => 'U');
          BIT_OS_SEL_5               : in    std_logic_vector(2 downto 1) := (others => 'U');
          BIT_OS_SEL_7_0             : in    std_logic := 'U';
          BIT_OS_SEL_6_0             : in    std_logic := 'U';
          BIT_OS_SEL_0               : in    std_logic := 'U';
          ELK_RX_SER_WORD_11         : out   std_logic_vector(7 downto 0);
          OP_MODE_c_0                : in    std_logic := 'U';
          PATT_ELK_DAT_11            : in    std_logic_vector(7 downto 0) := (others => 'U');
          MASTER_DCB_POR_B_i_0_i     : in    std_logic := 'U';
          ELK11_DAT_N                : inout   std_logic;
          ELK11_DAT_P                : inout   std_logic;
          DCB_SALT_SEL_c_i           : in    std_logic := 'U';
          CCC_160M_FXD               : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_5  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_16 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_10 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_2  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_11 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_7  : in    std_logic := 'U';
          CLK_40M_GL                 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_0  : in    std_logic := 'U';
          DEV_RST_B_c_0              : in    std_logic := 'U';
          CCC_160M_ADJ               : in    std_logic := 'U'
        );
  end component;

  component GP_PATT_GEN_1_0
    port( ELKS_ADDRB            : out   std_logic_vector(7 downto 0);
          ELK_RX_SER_WORD_0     : in    std_logic_vector(7 downto 0) := (others => 'U');
          ELKS_STOP_ADDR        : in    std_logic_vector(7 downto 0) := (others => 'U');
          ELKS_STRT_ADDR        : in    std_logic_vector(7 downto 0) := (others => 'U');
          OP_MODE_0             : in    std_logic := 'U';
          OP_MODE_c_0           : in    std_logic := 'U';
          ELKS_ADDRB_0_0        : out   std_logic;
          ELKS_ADDRB_0_2        : out   std_logic;
          ELKS_ADDRB_0_4        : out   std_logic;
          P_MASTER_POR_B_c_32   : in    std_logic := 'U';
          P_MASTER_POR_B_c_26   : in    std_logic := 'U';
          P_MASTER_POR_B_c_25   : in    std_logic := 'U';
          P_MASTER_POR_B_c_23   : in    std_logic := 'U';
          P_MASTER_POR_B_c_7    : in    std_logic := 'U';
          P_MASTER_POR_B_c_11   : in    std_logic := 'U';
          P_MASTER_POR_B_c_29   : in    std_logic := 'U';
          DCB_SALT_SEL_c_i      : in    std_logic := 'U';
          P_MASTER_POR_B_c_2    : in    std_logic := 'U';
          P_MASTER_POR_B_c_12   : in    std_logic := 'U';
          ELKS_RWB              : out   std_logic;
          P_MASTER_POR_B_c_13   : in    std_logic := 'U';
          ELKS_RAM_BLKB_EN      : out   std_logic;
          P_USB_MASTER_EN_c     : in    std_logic := 'U';
          ALIGN_ACTIVE          : in    std_logic := 'U';
          P_MASTER_POR_B_c_34_0 : in    std_logic := 'U';
          P_MASTER_POR_B_c_32_0 : in    std_logic := 'U';
          P_MASTER_POR_B_c_31_0 : in    std_logic := 'U';
          CLK_40M_GL            : in    std_logic := 'U'
        );
  end component;

  component BUFF
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SER320M_3_34
    port( TFC_TX_DAT             : in    std_logic_vector(7 downto 0) := (others => 'U');
          TFC_OUT_R              : out   std_logic;
          TFC_OUT_F              : out   std_logic;
          MASTER_DCB_POR_B_i_0_i : in    std_logic := 'U';
          CCC_160M_FXD           : in    std_logic := 'U';
          CLK_40M_GL             : in    std_logic := 'U'
        );
  end component;

  component SER320M_3_34_0
    port( ELK0_TX_DAT                : in    std_logic_vector(7 downto 0) := (others => 'U');
          MASTER_SALT_POR_B_i_0_i_17 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_3  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_7  : in    std_logic := 'U';
          ELK0_OUT_R_i_0             : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_10 : in    std_logic := 'U';
          ELK0_OUT_F_i_0             : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_5  : in    std_logic := 'U';
          CLK_40M_GL                 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_13 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_14 : in    std_logic := 'U';
          CCC_160M_FXD               : in    std_logic := 'U'
        );
  end component;

  component ELINK_SLAVE_15_7
    port( BIT_OS_SEL_3_0             : in    std_logic := 'U';
          BIT_OS_SEL_4               : in    std_logic_vector(2 downto 1) := (others => 'U');
          BIT_OS_SEL_6               : in    std_logic_vector(2 downto 1) := (others => 'U');
          BIT_OS_SEL_5_0             : in    std_logic := 'U';
          ELK_RX_SER_WORD_12         : out   std_logic_vector(7 downto 0);
          OP_MODE_c_2_0              : in    std_logic := 'U';
          OP_MODE_c_3_0              : in    std_logic := 'U';
          PATT_ELK_DAT_12            : in    std_logic_vector(7 downto 0) := (others => 'U');
          MASTER_DCB_POR_B_i_0_i     : in    std_logic := 'U';
          ELK12_DAT_N                : inout   std_logic;
          ELK12_DAT_P                : inout   std_logic;
          DCB_SALT_SEL_c_i           : in    std_logic := 'U';
          CCC_160M_FXD               : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_6  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_12 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_8  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_0  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_10 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_15 : in    std_logic := 'U';
          CLK_40M_GL                 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_2  : in    std_logic := 'U';
          DEV_RST_B_c                : in    std_logic := 'U';
          CCC_160M_ADJ               : in    std_logic := 'U'
        );
  end component;

  component ELINK_SLAVE_15_8
    port( BIT_OS_SEL_2_0             : in    std_logic := 'U';
          BIT_OS_SEL_3               : in    std_logic_vector(2 downto 1) := (others => 'U');
          BIT_OS_SEL_6_0             : in    std_logic := 'U';
          BIT_OS_SEL_5_0             : in    std_logic := 'U';
          BIT_OS_SEL_4_0             : in    std_logic := 'U';
          ELK_RX_SER_WORD_13         : out   std_logic_vector(7 downto 0);
          OP_MODE_c_6_0              : in    std_logic := 'U';
          OP_MODE_c_0                : in    std_logic := 'U';
          PATT_ELK_DAT_13            : in    std_logic_vector(7 downto 0) := (others => 'U');
          MASTER_DCB_POR_B_i_0_i     : in    std_logic := 'U';
          ELK13_DAT_N                : inout   std_logic;
          ELK13_DAT_P                : inout   std_logic;
          DCB_SALT_SEL_c_i           : in    std_logic := 'U';
          CCC_160M_FXD               : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_6  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_1  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_9  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_16 : in    std_logic := 'U';
          CLK_40M_GL                 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_4  : in    std_logic := 'U';
          DEV_RST_B_c                : in    std_logic := 'U';
          CCC_160M_ADJ               : in    std_logic := 'U'
        );
  end component;

  component SYNC_DAT_SEL_0
    port( ELK0_TX_DAT                : out   std_logic_vector(7 downto 0);
          PATT_ELK_DAT_0             : in    std_logic_vector(7 downto 0) := (others => 'U');
          OP_MODE_c_4_0              : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_10 : in    std_logic := 'U';
          CLK_40M_GL                 : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component EXEC_MODE_CNTL
    port( CLK60MHZ                   : in    std_logic := 'U';
          P_USB_MASTER_EN_c_1_0      : out   std_logic;
          P_USB_MASTER_EN_c_2_0      : out   std_logic;
          P_USB_MASTER_EN_c_22_0     : out   std_logic;
          P_USB_MASTER_EN_c_22       : out   std_logic;
          P_USB_MASTER_EN_c_21       : out   std_logic;
          P_USB_MASTER_EN_c_20       : out   std_logic;
          P_USB_MASTER_EN_c_19       : out   std_logic;
          P_USB_MASTER_EN_c_18       : out   std_logic;
          P_USB_MASTER_EN_c_17       : out   std_logic;
          P_USB_MASTER_EN_c_16       : out   std_logic;
          P_USB_MASTER_EN_c_15       : out   std_logic;
          P_USB_MASTER_EN_c_14       : out   std_logic;
          P_USB_MASTER_EN_c_13       : out   std_logic;
          P_USB_MASTER_EN_c_12       : out   std_logic;
          P_USB_MASTER_EN_c_11       : out   std_logic;
          P_USB_MASTER_EN_c_10       : out   std_logic;
          P_USB_MASTER_EN_c_9        : out   std_logic;
          P_USB_MASTER_EN_c_8        : out   std_logic;
          P_USB_MASTER_EN_c_7        : out   std_logic;
          P_USB_MASTER_EN_c_6        : out   std_logic;
          P_USB_MASTER_EN_c_5        : out   std_logic;
          P_USB_MASTER_EN_c_4        : out   std_logic;
          P_USB_MASTER_EN_c_3        : out   std_logic;
          P_USB_MASTER_EN_c_2        : out   std_logic;
          P_USB_MASTER_EN_c_1        : out   std_logic;
          P_USB_MASTER_EN_c_0        : out   std_logic;
          P_USB_MASTER_EN_c          : out   std_logic;
          P_MASTER_POR_B_c           : out   std_logic;
          CCC_MAIN_LOCK              : in    std_logic := 'U';
          DCB_SALT_SEL_c             : in    std_logic := 'U';
          DEV_RST_B_c_1              : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i    : out   std_logic;
          MASTER_DCB_POR_B_i_0_i     : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_0  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_1  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_2  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_3  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_4  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_5  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_6  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_7  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_8  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_9  : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_10 : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_11 : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_12 : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_13 : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_14 : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_15 : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_16 : out   std_logic;
          MASTER_SALT_POR_B_i_0_i_17 : out   std_logic;
          P_MASTER_POR_B_c_1         : out   std_logic;
          P_MASTER_POR_B_c_2         : out   std_logic;
          P_MASTER_POR_B_c_3         : out   std_logic;
          P_MASTER_POR_B_c_4         : out   std_logic;
          P_MASTER_POR_B_c_5         : out   std_logic;
          P_MASTER_POR_B_c_6         : out   std_logic;
          P_MASTER_POR_B_c_7         : out   std_logic;
          P_MASTER_POR_B_c_8         : out   std_logic;
          P_MASTER_POR_B_c_9         : out   std_logic;
          P_MASTER_POR_B_c_10        : out   std_logic;
          P_MASTER_POR_B_c_11        : out   std_logic;
          P_MASTER_POR_B_c_12        : out   std_logic;
          P_MASTER_POR_B_c_13        : out   std_logic;
          P_MASTER_POR_B_c_14        : out   std_logic;
          P_MASTER_POR_B_c_15        : out   std_logic;
          P_MASTER_POR_B_c_16        : out   std_logic;
          P_MASTER_POR_B_c_17        : out   std_logic;
          P_MASTER_POR_B_c_18        : out   std_logic;
          P_MASTER_POR_B_c_19        : out   std_logic;
          P_MASTER_POR_B_c_20        : out   std_logic;
          P_MASTER_POR_B_c_21        : out   std_logic;
          P_MASTER_POR_B_c_22        : out   std_logic;
          P_MASTER_POR_B_c_23        : out   std_logic;
          P_MASTER_POR_B_c_24        : out   std_logic;
          P_MASTER_POR_B_c_25        : out   std_logic;
          P_MASTER_POR_B_c_26        : out   std_logic;
          P_MASTER_POR_B_c_27        : out   std_logic;
          P_MASTER_POR_B_c_28        : out   std_logic;
          P_MASTER_POR_B_c_29        : out   std_logic;
          P_MASTER_POR_B_c_30        : out   std_logic;
          P_MASTER_POR_B_c_31        : out   std_logic;
          P_MASTER_POR_B_c_32        : out   std_logic;
          P_MASTER_POR_B_c_33        : out   std_logic;
          P_MASTER_POR_B_c_34        : out   std_logic;
          P_MASTER_POR_B_c_34_0      : out   std_logic;
          P_MASTER_POR_B_c_32_0      : out   std_logic;
          P_MASTER_POR_B_c_31_0      : out   std_logic;
          P_MASTER_POR_B_c_27_0      : out   std_logic;
          P_MASTER_POR_B_c_27_1      : out   std_logic;
          P_MASTER_POR_B_c_24_0      : out   std_logic;
          P_MASTER_POR_B_c_22_0      : out   std_logic;
          P_MASTER_POR_B_c_17_0      : out   std_logic;
          P_MASTER_POR_B_c_16_0      : out   std_logic;
          DEV_RST_B_c                : in    std_logic := 'U';
          CCC_160M_FXD               : in    std_logic := 'U';
          CLK_40M_GL                 : in    std_logic := 'U';
          P_MASTER_POR_B_c_0_0       : out   std_logic
        );
  end component;

  component ELINK_SLAVE_15_2
    port( BIT_OS_SEL_4               : in    std_logic_vector(2 downto 1) := (others => 'U');
          BIT_OS_SEL_6               : in    std_logic_vector(2 downto 1) := (others => 'U');
          BIT_OS_SEL_5_2             : in    std_logic := 'U';
          BIT_OS_SEL_5_0             : in    std_logic := 'U';
          BIT_OS_SEL_0               : in    std_logic := 'U';
          ELK_RX_SER_WORD_7          : out   std_logic_vector(7 downto 0);
          OP_MODE_c_4_0              : in    std_logic := 'U';
          PATT_ELK_DAT_7             : in    std_logic_vector(7 downto 0) := (others => 'U');
          MASTER_DCB_POR_B_i_0_i     : in    std_logic := 'U';
          ELK7_DAT_N                 : inout   std_logic;
          ELK7_DAT_P                 : inout   std_logic;
          DCB_SALT_SEL_c_i           : in    std_logic := 'U';
          CCC_160M_FXD               : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_11 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_12 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_8  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_2  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_13 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_14 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_10 : in    std_logic := 'U';
          CLK_40M_GL                 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_3  : in    std_logic := 'U';
          DEV_RST_B_c_1              : in    std_logic := 'U';
          CCC_160M_ADJ               : in    std_logic := 'U'
        );
  end component;

  component ELINK_SLAVE_15_9
    port( BIT_OS_SEL_2               : in    std_logic_vector(2 downto 1) := (others => 'U');
          BIT_OS_SEL_5_0             : in    std_logic := 'U';
          BIT_OS_SEL_3_0             : in    std_logic := 'U';
          BIT_OS_SEL_4               : in    std_logic_vector(1 downto 0) := (others => 'U');
          ELK_RX_SER_WORD_14         : out   std_logic_vector(7 downto 0);
          OP_MODE_c_2_0              : in    std_logic := 'U';
          PATT_ELK_DAT_14            : in    std_logic_vector(7 downto 0) := (others => 'U');
          MASTER_DCB_POR_B_i_0_i     : in    std_logic := 'U';
          ELK14_DAT_N                : inout   std_logic;
          ELK14_DAT_P                : inout   std_logic;
          DCB_SALT_SEL_c_i           : in    std_logic := 'U';
          CCC_160M_FXD               : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_7  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_15 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_12 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_0  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_10 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_5  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_2  : in    std_logic := 'U';
          CLK_40M_GL                 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_6  : in    std_logic := 'U';
          DEV_RST_B_c                : in    std_logic := 'U';
          CCC_160M_ADJ               : in    std_logic := 'U'
        );
  end component;

  component tristate_buf_0
    port( P_USB_MASTER_EN_c : in    std_logic := 'U';
          USB_WR_BI         : in    std_logic := 'U';
          USB_WR_B          : out   std_logic
        );
  end component;

  component ELINK_SLAVE_15
    port( BIT_OS_SEL_7_0             : in    std_logic := 'U';
          BIT_OS_SEL                 : in    std_logic_vector(2 downto 1) := (others => 'U');
          BIT_OS_SEL_0_0             : in    std_logic := 'U';
          BIT_OS_SEL_1               : in    std_logic_vector(1 downto 0) := (others => 'U');
          ELK_RX_SER_WORD_2          : out   std_logic_vector(7 downto 0);
          OP_MODE_c_1_0              : in    std_logic := 'U';
          PATT_ELK_DAT_2             : in    std_logic_vector(7 downto 0) := (others => 'U');
          MASTER_DCB_POR_B_i_0_i     : in    std_logic := 'U';
          ELK2_DAT_N                 : inout   std_logic;
          ELK2_DAT_P                 : inout   std_logic;
          DCB_SALT_SEL_c_i           : in    std_logic := 'U';
          CCC_160M_FXD               : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_8  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_12 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_5  : in    std_logic := 'U';
          CLK_40M_GL                 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_13 : in    std_logic := 'U';
          DEV_RST_B_c_0              : in    std_logic := 'U';
          CCC_160M_ADJ               : in    std_logic := 'U'
        );
  end component;

  component ELINK_SLAVE_INV_2_1
    port( BIT_OS_SEL_7_0             : in    std_logic := 'U';
          BIT_OS_SEL_6               : in    std_logic_vector(2 downto 1) := (others => 'U');
          BIT_OS_SEL_0_d0            : in    std_logic := 'U';
          BIT_OS_SEL_0               : in    std_logic_vector(1 downto 0) := (others => 'U');
          BIT_OS_SEL_1_0             : in    std_logic := 'U';
          ELK_RX_SER_WORD_4          : out   std_logic_vector(7 downto 0);
          OP_MODE_c_1_0              : in    std_logic := 'U';
          PATT_ELK_DAT_4             : in    std_logic_vector(7 downto 0) := (others => 'U');
          MASTER_DCB_POR_B_i_0_i     : in    std_logic := 'U';
          ELK4_DAT_N                 : inout   std_logic;
          ELK4_DAT_P                 : inout   std_logic;
          DCB_SALT_SEL_c_i           : in    std_logic := 'U';
          CCC_160M_FXD               : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_4  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_9  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_13 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_1  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_17 : in    std_logic := 'U';
          CLK_40M_GL                 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_16 : in    std_logic := 'U';
          DEV_RST_B_c                : in    std_logic := 'U';
          CCC_160M_ADJ               : in    std_logic := 'U'
        );
  end component;

  component DDR_BIDIR_LVDS_DUAL_CLK
    port( DCB_SALT_SEL_c : in    std_logic := 'U';
          TFC_DAT_0P     : inout   std_logic;
          TFC_DAT_0N     : inout   std_logic;
          TFC_OUT_R      : in    std_logic := 'U';
          TFC_OUT_F      : in    std_logic := 'U';
          CCC_160M_FXD   : in    std_logic := 'U';
          CCC_160M_ADJ   : in    std_logic := 'U';
          TFC_IN_DDR_R   : out   std_logic;
          TFC_IN_DDR_F   : out   std_logic
        );
  end component;

  component tristate_buf
    port( P_USB_MASTER_EN_c : in    std_logic := 'U';
          USB_RD_BI         : in    std_logic := 'U';
          USB_RD_B          : out   std_logic
        );
  end component;

  component REF_CLK_DIV_GEN
    port( DEV_RST_B_c_1   : in    std_logic := 'U';
          Y               : in    std_logic := 'U';
          CLK40M_10NS_REF : out   std_logic
        );
  end component;

  component ELINK_SLAVE_15_1
    port( BIT_OS_SEL_5               : in    std_logic_vector(2 downto 1) := (others => 'U');
          BIT_OS_SEL_7_0             : in    std_logic := 'U';
          BIT_OS_SEL_6_0             : in    std_logic := 'U';
          BIT_OS_SEL_0               : in    std_logic := 'U';
          ELK_RX_SER_WORD_6          : out   std_logic_vector(7 downto 0);
          OP_MODE_c_0_0              : in    std_logic := 'U';
          OP_MODE_c_1_0              : in    std_logic := 'U';
          PATT_ELK_DAT_6             : in    std_logic_vector(7 downto 0) := (others => 'U');
          MASTER_DCB_POR_B_i_0_i     : in    std_logic := 'U';
          ELK6_DAT_N                 : inout   std_logic;
          ELK6_DAT_P                 : inout   std_logic;
          DCB_SALT_SEL_c_i           : in    std_logic := 'U';
          CCC_160M_FXD               : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_10 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_16 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_12 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_3  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_9  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_6  : in    std_logic := 'U';
          CLK_40M_GL                 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_1  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_2  : in    std_logic := 'U';
          DEV_RST_B_c_1              : in    std_logic := 'U';
          CCC_160M_ADJ               : in    std_logic := 'U'
        );
  end component;

  component TOP_MASTER_DES320M
    port( BIT_OS_SEL_7_0        : out   std_logic;
          BIT_OS_SEL_6          : out   std_logic_vector(2 downto 1);
          BIT_OS_SEL_5          : out   std_logic_vector(2 downto 0);
          BIT_OS_SEL_4          : out   std_logic_vector(2 downto 0);
          BIT_OS_SEL_3          : out   std_logic_vector(2 downto 0);
          BIT_OS_SEL_2          : out   std_logic_vector(2 downto 0);
          BIT_OS_SEL_1          : out   std_logic_vector(2 downto 0);
          BIT_OS_SEL_0          : out   std_logic_vector(2 downto 0);
          OP_MODE_c_0           : in    std_logic := 'U';
          BIT_OS_SEL            : out   std_logic_vector(2 downto 0);
          TFC_RX_SER_WORD       : out   std_logic_vector(7 downto 0);
          ELK_RX_SER_WORD_0     : out   std_logic_vector(7 downto 0);
          P_MASTER_POR_B_c_27_0 : in    std_logic := 'U';
          P_MASTER_POR_B_c_27_1 : in    std_logic := 'U';
          P_MASTER_POR_B_c_16_0 : in    std_logic := 'U';
          P_MASTER_POR_B_c_17_0 : in    std_logic := 'U';
          P_MASTER_POR_B_c_24_0 : in    std_logic := 'U';
          TFC_SYNC_DET_1        : out   std_logic;
          ELK0_SYNC_DET_1       : out   std_logic;
          DCB_SALT_SEL_c        : in    std_logic := 'U';
          TFC_IN_R              : in    std_logic := 'U';
          ELK0_IN_R             : in    std_logic := 'U';
          TFC_IN_F              : in    std_logic := 'U';
          ELK0_IN_F             : in    std_logic := 'U';
          ALL_PLL_LOCK_c        : out   std_logic;
          CCC_MAIN_LOCK         : in    std_logic := 'U';
          P_MASTER_POR_B_c_31_0 : in    std_logic := 'U';
          P_MASTER_POR_B_c_26   : in    std_logic := 'U';
          P_MASTER_POR_B_c_32   : in    std_logic := 'U';
          P_MASTER_POR_B_c_24   : in    std_logic := 'U';
          P_MASTER_POR_B_c_5    : in    std_logic := 'U';
          P_MASTER_POR_B_c_4    : in    std_logic := 'U';
          P_MASTER_POR_B_c_2    : in    std_logic := 'U';
          P_MASTER_POR_B_c_3    : in    std_logic := 'U';
          P_MASTER_POR_B_c_9    : in    std_logic := 'U';
          P_MASTER_POR_B_c_21   : in    std_logic := 'U';
          P_MASTER_POR_B_c_15   : in    std_logic := 'U';
          P_MASTER_POR_B_c_16   : in    std_logic := 'U';
          P_MASTER_POR_B_c_12   : in    std_logic := 'U';
          P_MASTER_POR_B_c_11   : in    std_logic := 'U';
          P_MASTER_POR_B_c_7    : in    std_logic := 'U';
          ALIGN_ACTIVE          : out   std_logic;
          P_MASTER_POR_B_c_27   : in    std_logic := 'U';
          P_MASTER_POR_B_c_10   : in    std_logic := 'U';
          P_MASTER_POR_B_c_17   : in    std_logic := 'U';
          P_MASTER_POR_B_c_1    : in    std_logic := 'U';
          P_MASTER_POR_B_c_20   : in    std_logic := 'U';
          P_MASTER_POR_B_c_8    : in    std_logic := 'U';
          P_MASTER_POR_B_c_29   : in    std_logic := 'U';
          P_MASTER_POR_B_c_30   : in    std_logic := 'U';
          P_MASTER_POR_B_c_28   : in    std_logic := 'U';
          P_MASTER_POR_B_c_34_0 : in    std_logic := 'U';
          P_MASTER_POR_B_c_32_0 : in    std_logic := 'U';
          CCC_160M_FXD          : in    std_logic := 'U';
          P_MASTER_POR_B_c_23   : in    std_logic := 'U';
          P_MASTER_POR_B_c      : in    std_logic := 'U';
          CLK_40M_BUF_RECD      : in    std_logic := 'U';
          CLK_40M_GL            : in    std_logic := 'U';
          P_MASTER_POR_B_c_22_0 : in    std_logic := 'U';
          P_MASTER_POR_B_c_14   : in    std_logic := 'U';
          P_MASTER_POR_B_c_6    : in    std_logic := 'U';
          P_MASTER_POR_B_c_25   : in    std_logic := 'U';
          P_MASTER_POR_B_c_13   : in    std_logic := 'U';
          P_MASTER_POR_B_c_22   : in    std_logic := 'U';
          P_MASTER_POR_B_c_31   : in    std_logic := 'U';
          P_MASTER_POR_B_c_33   : in    std_logic := 'U';
          P_MASTER_POR_B_c_18   : in    std_logic := 'U';
          P_MASTER_POR_B_c_19   : in    std_logic := 'U';
          P_MASTER_POR_B_c_34   : in    std_logic := 'U';
          CCC_160M_ADJ          : out   std_logic
        );
  end component;

  component ELINK_SLAVE_15_11
    port( BIT_OS_SEL_1               : in    std_logic_vector(2 downto 1) := (others => 'U');
          BIT_OS_SEL_2_0             : in    std_logic := 'U';
          BIT_OS_SEL_3               : in    std_logic_vector(2 downto 0) := (others => 'U');
          ELK_RX_SER_WORD_16         : out   std_logic_vector(7 downto 0);
          OP_MODE_c_2_0              : in    std_logic := 'U';
          PATT_ELK_DAT_16            : in    std_logic_vector(7 downto 0) := (others => 'U');
          MASTER_DCB_POR_B_i_0_i     : in    std_logic := 'U';
          ELK16_DAT_N                : inout   std_logic;
          ELK16_DAT_P                : inout   std_logic;
          DCB_SALT_SEL_c_i           : in    std_logic := 'U';
          CCC_160M_FXD               : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_8  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_1  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_16 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_0  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_10 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_14 : in    std_logic := 'U';
          CLK_40M_GL                 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_9  : in    std_logic := 'U';
          DEV_RST_B_c_1              : in    std_logic := 'U';
          CCC_160M_ADJ               : in    std_logic := 'U'
        );
  end component;

  component tristate_buf_2
    port( P_USB_MASTER_EN_c : in    std_logic := 'U';
          USB_SIWU_BI       : in    std_logic := 'U';
          USB_SIWU_B        : out   std_logic
        );
  end component;

  component INV
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DDR_BIDIR_LVDS_DUAL_CLK_0
    port( DCB_SALT_SEL_c_i : in    std_logic := 'U';
          ELK0_DAT_P       : inout   std_logic;
          ELK0_DAT_N       : inout   std_logic;
          ELK0_OUT_R_i_0   : in    std_logic := 'U';
          ELK0_OUT_F_i_0   : in    std_logic := 'U';
          CCC_160M_FXD     : in    std_logic := 'U';
          CCC_160M_ADJ     : in    std_logic := 'U';
          ELK0_IN_DDR_F_i  : out   std_logic;
          ELK0_IN_DDR_R_i  : out   std_logic
        );
  end component;

  component LVDS_CLK_IN
    port( CLK200_N : in    std_logic := 'U';
          CLK200_P : in    std_logic := 'U';
          Y        : out   std_logic
        );
  end component;

  component ELINK_SLAVE_15_14
    port( BIT_OS_SEL_0_d0            : in    std_logic := 'U';
          BIT_OS_SEL_0               : in    std_logic_vector(2 downto 1) := (others => 'U');
          BIT_OS_SEL_1               : in    std_logic_vector(2 downto 1) := (others => 'U');
          BIT_OS_SEL_2_0             : in    std_logic := 'U';
          ELK_RX_SER_WORD_19         : out   std_logic_vector(7 downto 0);
          OP_MODE_c_5_0              : in    std_logic := 'U';
          OP_MODE_c_6_0              : in    std_logic := 'U';
          PATT_ELK_DAT_19            : in    std_logic_vector(7 downto 0) := (others => 'U');
          MASTER_DCB_POR_B_i_0_i     : in    std_logic := 'U';
          ELK19_DAT_N                : inout   std_logic;
          ELK19_DAT_P                : inout   std_logic;
          DCB_SALT_SEL_c_i           : in    std_logic := 'U';
          CCC_160M_FXD               : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_10 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_16 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_12 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_8  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_0  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_7  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_4  : in    std_logic := 'U';
          CLK_40M_GL                 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_15 : in    std_logic := 'U';
          DEV_RST_B_c_0              : in    std_logic := 'U';
          CCC_160M_ADJ               : in    std_logic := 'U'
        );
  end component;

  component ELINK_SLAVE_15_4
    port( BIT_OS_SEL_2               : in    std_logic_vector(2 downto 1) := (others => 'U');
          BIT_OS_SEL_3               : in    std_logic_vector(2 downto 1) := (others => 'U');
          BIT_OS_SEL_5               : in    std_logic_vector(2 downto 1) := (others => 'U');
          BIT_OS_SEL_4_0             : in    std_logic := 'U';
          ELK_RX_SER_WORD_9          : out   std_logic_vector(7 downto 0);
          OP_MODE_c_3_0              : in    std_logic := 'U';
          PATT_ELK_DAT_9             : in    std_logic_vector(7 downto 0) := (others => 'U');
          MASTER_DCB_POR_B_i_0_i     : in    std_logic := 'U';
          ELK9_DAT_N                 : inout   std_logic;
          ELK9_DAT_P                 : inout   std_logic;
          DCB_SALT_SEL_c_i           : in    std_logic := 'U';
          CCC_160M_FXD               : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_12 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_16 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_13 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_2  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_3  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_4  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_0  : in    std_logic := 'U';
          CLK_40M_GL                 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_7  : in    std_logic := 'U';
          DEV_RST_B_c_0              : in    std_logic := 'U';
          CCC_160M_ADJ               : in    std_logic := 'U'
        );
  end component;

  component GP_PATT_GEN_1
    port( TFC_ADDRB              : out   std_logic_vector(7 downto 0);
          TFC_RX_SER_WORD        : in    std_logic_vector(7 downto 0) := (others => 'U');
          TFC_STOP_ADDR          : in    std_logic_vector(7 downto 0) := (others => 'U');
          TFC_STRT_ADDR          : in    std_logic_vector(7 downto 0) := (others => 'U');
          OP_MODE_0              : in    std_logic := 'U';
          OP_MODE_c_0            : in    std_logic := 'U';
          P_MASTER_POR_B_c_24    : in    std_logic := 'U';
          P_MASTER_POR_B_c       : in    std_logic := 'U';
          P_MASTER_POR_B_c_31    : in    std_logic := 'U';
          P_MASTER_POR_B_c_30    : in    std_logic := 'U';
          P_MASTER_POR_B_c_1     : in    std_logic := 'U';
          P_MASTER_POR_B_c_5     : in    std_logic := 'U';
          P_MASTER_POR_B_c_4     : in    std_logic := 'U';
          P_MASTER_POR_B_c_28    : in    std_logic := 'U';
          DCB_SALT_SEL_c         : in    std_logic := 'U';
          P_MASTER_POR_B_c_15    : in    std_logic := 'U';
          P_MASTER_POR_B_c_16_0  : in    std_logic := 'U';
          TFC_RWB                : out   std_logic;
          P_MASTER_POR_B_c_9     : in    std_logic := 'U';
          TFC_RAM_BLKB_EN        : out   std_logic;
          P_USB_MASTER_EN_c_22_0 : in    std_logic := 'U';
          ALIGN_ACTIVE           : in    std_logic := 'U';
          P_MASTER_POR_B_c_27_1  : in    std_logic := 'U';
          CLK_40M_GL             : in    std_logic := 'U'
        );
  end component;

  component ELINK_SLAVE_15_3
    port( BIT_OS_SEL_4_0             : in    std_logic := 'U';
          BIT_OS_SEL_3               : in    std_logic_vector(2 downto 1) := (others => 'U');
          BIT_OS_SEL_6_0             : in    std_logic := 'U';
          BIT_OS_SEL_5               : in    std_logic_vector(1 downto 0) := (others => 'U');
          ELK_RX_SER_WORD_8          : out   std_logic_vector(7 downto 0);
          OP_MODE_c_0_0              : in    std_logic := 'U';
          PATT_ELK_DAT_8             : in    std_logic_vector(7 downto 0) := (others => 'U');
          MASTER_DCB_POR_B_i_0_i     : in    std_logic := 'U';
          ELK8_DAT_N                 : inout   std_logic;
          ELK8_DAT_P                 : inout   std_logic;
          DCB_SALT_SEL_c_i           : in    std_logic := 'U';
          CCC_160M_FXD               : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_12 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_2  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_3  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i    : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_15 : in    std_logic := 'U';
          CLK_40M_GL                 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_5  : in    std_logic := 'U';
          DEV_RST_B_c_1              : in    std_logic := 'U';
          DEV_RST_B_c_0              : in    std_logic := 'U';
          CCC_160M_ADJ               : in    std_logic := 'U'
        );
  end component;

  component ELINK_SLAVE_15_12
    port( BIT_OS_SEL_0_0             : in    std_logic := 'U';
          BIT_OS_SEL_1_0             : in    std_logic := 'U';
          BIT_OS_SEL_2               : in    std_logic_vector(2 downto 0) := (others => 'U');
          BIT_OS_SEL_3_0             : in    std_logic := 'U';
          ELK_RX_SER_WORD_17         : out   std_logic_vector(7 downto 0);
          OP_MODE_c_6_0              : in    std_logic := 'U';
          PATT_ELK_DAT_17            : in    std_logic_vector(7 downto 0) := (others => 'U');
          MASTER_DCB_POR_B_i_0_i     : in    std_logic := 'U';
          ELK17_DAT_N                : inout   std_logic;
          ELK17_DAT_P                : inout   std_logic;
          DCB_SALT_SEL_c_i           : in    std_logic := 'U';
          CCC_160M_FXD               : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_9  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_8  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_0  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_17 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_14 : in    std_logic := 'U';
          CLK_40M_GL                 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_11 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_12 : in    std_logic := 'U';
          DEV_RST_B_c_1              : in    std_logic := 'U';
          CCC_160M_ADJ               : in    std_logic := 'U'
        );
  end component;

  component ELINK_SLAVE_15_10
    port( BIT_OS_SEL_1_0            : in    std_logic := 'U';
          BIT_OS_SEL_2              : in    std_logic_vector(2 downto 1) := (others => 'U');
          BIT_OS_SEL_4_0            : in    std_logic := 'U';
          BIT_OS_SEL_3              : in    std_logic_vector(1 downto 0) := (others => 'U');
          ELK_RX_SER_WORD_15        : out   std_logic_vector(7 downto 0);
          OP_MODE_c_6_0             : in    std_logic := 'U';
          PATT_ELK_DAT_15           : in    std_logic_vector(7 downto 0) := (others => 'U');
          MASTER_DCB_POR_B_i_0_i    : in    std_logic := 'U';
          ELK15_DAT_N               : inout   std_logic;
          ELK15_DAT_P               : inout   std_logic;
          DCB_SALT_SEL_c_i          : in    std_logic := 'U';
          CCC_160M_FXD              : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_5 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_9 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_1 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_6 : in    std_logic := 'U';
          CLK_40M_GL                : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_7 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_8 : in    std_logic := 'U';
          DEV_RST_B_c_1             : in    std_logic := 'U';
          CCC_160M_ADJ              : in    std_logic := 'U'
        );
  end component;

  component BIDIR_LVDS_IO
    port( EXT_INT_REF_SEL_c : in    std_logic := 'U';
          CLK40M_10NS_REF   : in    std_logic := 'U';
          CLK_40M_BUF_RECD  : out   std_logic;
          BIDIR_CLK40M_P    : inout   std_logic;
          BIDIR_CLK40M_N    : inout   std_logic
        );
  end component;

  component LVDS_BUFOUT
    port( CLK_40M_BUF_RECD : in    std_logic := 'U';
          TX_CLK40M_P      : out   std_logic;
          TX_CLK40M_N      : out   std_logic
        );
  end component;

  component ELINK_SLAVE_15_0
    port( BIT_OS_SEL_5               : in    std_logic_vector(2 downto 1) := (others => 'U');
          BIT_OS_SEL_6               : in    std_logic_vector(2 downto 1) := (others => 'U');
          BIT_OS_SEL_7_0             : in    std_logic := 'U';
          BIT_OS_SEL_0_d0            : in    std_logic := 'U';
          BIT_OS_SEL_0_0             : in    std_logic := 'U';
          ELK_RX_SER_WORD_5          : out   std_logic_vector(7 downto 0);
          OP_MODE_c_4_0              : in    std_logic := 'U';
          OP_MODE_c_5_0              : in    std_logic := 'U';
          PATT_ELK_DAT_5             : in    std_logic_vector(7 downto 0) := (others => 'U');
          MASTER_DCB_POR_B_i_0_i     : in    std_logic := 'U';
          ELK5_DAT_N                 : inout   std_logic;
          ELK5_DAT_P                 : inout   std_logic;
          DCB_SALT_SEL_c_i           : in    std_logic := 'U';
          CCC_160M_FXD               : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_9  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_8  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_5  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_3  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_14 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_6  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_2  : in    std_logic := 'U';
          CLK_40M_GL                 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_17 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i    : in    std_logic := 'U';
          DEV_RST_B_c                : in    std_logic := 'U';
          CCC_160M_ADJ               : in    std_logic := 'U'
        );
  end component;

  component ELINK_SLAVE_15_5
    port( BIT_OS_SEL_6_0             : in    std_logic := 'U';
          BIT_OS_SEL_5               : in    std_logic_vector(2 downto 1) := (others => 'U');
          BIT_OS_SEL_7_0             : in    std_logic := 'U';
          BIT_OS_SEL_0_d0            : in    std_logic := 'U';
          BIT_OS_SEL_0_0             : in    std_logic := 'U';
          ELK_RX_SER_WORD_10         : out   std_logic_vector(7 downto 0);
          OP_MODE_c_3_0              : in    std_logic := 'U';
          PATT_ELK_DAT_10            : in    std_logic_vector(7 downto 0) := (others => 'U');
          MASTER_DCB_POR_B_i_0_i     : in    std_logic := 'U';
          ELK10_DAT_N                : inout   std_logic;
          ELK10_DAT_P                : inout   std_logic;
          DCB_SALT_SEL_c_i           : in    std_logic := 'U';
          CCC_160M_FXD               : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_5  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_8  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_1  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_11 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_6  : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_3  : in    std_logic := 'U';
          CLK_40M_GL                 : in    std_logic := 'U';
          MASTER_SALT_POR_B_i_0_i_17 : in    std_logic := 'U';
          DEV_RST_B_c_0              : in    std_logic := 'U';
          CCC_160M_ADJ               : in    std_logic := 'U'
        );
  end component;

    signal Y, CLK40M_10NS_REF, CLK_40M_BUF_RECD, CCC_MAIN_LOCK, 
        CLK60MHZ, \VCC\, \GND\, \PATT_TFC_DAT[0]\, 
        \PATT_TFC_DAT[1]\, \PATT_TFC_DAT[2]\, \PATT_TFC_DAT[3]\, 
        \PATT_TFC_DAT[4]\, \PATT_TFC_DAT[5]\, \PATT_TFC_DAT[6]\, 
        \PATT_TFC_DAT[7]\, \TFC_TX_DAT[0]\, \TFC_TX_DAT[1]\, 
        \TFC_TX_DAT[2]\, \TFC_TX_DAT[3]\, \TFC_TX_DAT[4]\, 
        \TFC_TX_DAT[5]\, \TFC_TX_DAT[6]\, \TFC_TX_DAT[7]\, 
        TFC_OUT_R, TFC_OUT_F, TFC_IN_DDR_R, TFC_IN_DDR_F, 
        \PATT_ELK_DAT_0[0]\, \PATT_ELK_DAT_0[1]\, 
        \PATT_ELK_DAT_0[2]\, \PATT_ELK_DAT_0[3]\, 
        \PATT_ELK_DAT_0[4]\, \PATT_ELK_DAT_0[5]\, 
        \PATT_ELK_DAT_0[6]\, \PATT_ELK_DAT_0[7]\, 
        \ELK0_TX_DAT[0]\, \ELK0_TX_DAT[1]\, \ELK0_TX_DAT[2]\, 
        \ELK0_TX_DAT[3]\, \ELK0_TX_DAT[4]\, \ELK0_TX_DAT[5]\, 
        \ELK0_TX_DAT[6]\, \ELK0_TX_DAT[7]\, \ELK0_IN_R\, 
        \ELK0_IN_F\, \TFC_IN_R\, \TFC_IN_F\, \TFC_RX_SER_WORD[0]\, 
        \TFC_RX_SER_WORD[1]\, \TFC_RX_SER_WORD[2]\, 
        \TFC_RX_SER_WORD[3]\, \TFC_RX_SER_WORD[4]\, 
        \TFC_RX_SER_WORD[5]\, \TFC_RX_SER_WORD[6]\, 
        \TFC_RX_SER_WORD[7]\, \ELK_RX_SER_WORD_0[0]\, 
        \ELK_RX_SER_WORD_0[1]\, \ELK_RX_SER_WORD_0[2]\, 
        \ELK_RX_SER_WORD_0[3]\, \ELK_RX_SER_WORD_0[4]\, 
        \ELK_RX_SER_WORD_0[5]\, \ELK_RX_SER_WORD_0[6]\, 
        \ELK_RX_SER_WORD_0[7]\, \BIT_OS_SEL[0]\, \BIT_OS_SEL[1]\, 
        \BIT_OS_SEL[2]\, ALIGN_ACTIVE, \PATT_ELK_DAT_1[0]\, 
        \PATT_ELK_DAT_1[1]\, \PATT_ELK_DAT_1[2]\, 
        \PATT_ELK_DAT_1[3]\, \PATT_ELK_DAT_1[4]\, 
        \PATT_ELK_DAT_1[5]\, \PATT_ELK_DAT_1[6]\, 
        \PATT_ELK_DAT_1[7]\, \ELK_RX_SER_WORD_1[0]\, 
        \ELK_RX_SER_WORD_1[1]\, \ELK_RX_SER_WORD_1[2]\, 
        \ELK_RX_SER_WORD_1[3]\, \ELK_RX_SER_WORD_1[4]\, 
        \ELK_RX_SER_WORD_1[5]\, \ELK_RX_SER_WORD_1[6]\, 
        \ELK_RX_SER_WORD_1[7]\, \PATT_ELK_DAT_2[0]\, 
        \PATT_ELK_DAT_2[1]\, \PATT_ELK_DAT_2[2]\, 
        \PATT_ELK_DAT_2[3]\, \PATT_ELK_DAT_2[4]\, 
        \PATT_ELK_DAT_2[5]\, \PATT_ELK_DAT_2[6]\, 
        \PATT_ELK_DAT_2[7]\, \ELK_RX_SER_WORD_2[0]\, 
        \ELK_RX_SER_WORD_2[1]\, \ELK_RX_SER_WORD_2[2]\, 
        \ELK_RX_SER_WORD_2[3]\, \ELK_RX_SER_WORD_2[4]\, 
        \ELK_RX_SER_WORD_2[5]\, \ELK_RX_SER_WORD_2[6]\, 
        \ELK_RX_SER_WORD_2[7]\, \PATT_ELK_DAT_3[0]\, 
        \PATT_ELK_DAT_3[1]\, \PATT_ELK_DAT_3[2]\, 
        \PATT_ELK_DAT_3[3]\, \PATT_ELK_DAT_3[4]\, 
        \PATT_ELK_DAT_3[5]\, \PATT_ELK_DAT_3[6]\, 
        \PATT_ELK_DAT_3[7]\, \ELK_RX_SER_WORD_3[0]\, 
        \ELK_RX_SER_WORD_3[1]\, \ELK_RX_SER_WORD_3[2]\, 
        \ELK_RX_SER_WORD_3[3]\, \ELK_RX_SER_WORD_3[4]\, 
        \ELK_RX_SER_WORD_3[5]\, \ELK_RX_SER_WORD_3[6]\, 
        \ELK_RX_SER_WORD_3[7]\, \PATT_ELK_DAT_4[0]\, 
        \PATT_ELK_DAT_4[1]\, \PATT_ELK_DAT_4[2]\, 
        \PATT_ELK_DAT_4[3]\, \PATT_ELK_DAT_4[4]\, 
        \PATT_ELK_DAT_4[5]\, \PATT_ELK_DAT_4[6]\, 
        \PATT_ELK_DAT_4[7]\, \ELK_RX_SER_WORD_4[0]\, 
        \ELK_RX_SER_WORD_4[1]\, \ELK_RX_SER_WORD_4[2]\, 
        \ELK_RX_SER_WORD_4[3]\, \ELK_RX_SER_WORD_4[4]\, 
        \ELK_RX_SER_WORD_4[5]\, \ELK_RX_SER_WORD_4[6]\, 
        \ELK_RX_SER_WORD_4[7]\, \PATT_ELK_DAT_5[0]\, 
        \PATT_ELK_DAT_5[1]\, \PATT_ELK_DAT_5[2]\, 
        \PATT_ELK_DAT_5[3]\, \PATT_ELK_DAT_5[4]\, 
        \PATT_ELK_DAT_5[5]\, \PATT_ELK_DAT_5[6]\, 
        \PATT_ELK_DAT_5[7]\, \ELK_RX_SER_WORD_5[0]\, 
        \ELK_RX_SER_WORD_5[1]\, \ELK_RX_SER_WORD_5[2]\, 
        \ELK_RX_SER_WORD_5[3]\, \ELK_RX_SER_WORD_5[4]\, 
        \ELK_RX_SER_WORD_5[5]\, \ELK_RX_SER_WORD_5[6]\, 
        \ELK_RX_SER_WORD_5[7]\, \PATT_ELK_DAT_6[0]\, 
        \PATT_ELK_DAT_6[1]\, \PATT_ELK_DAT_6[2]\, 
        \PATT_ELK_DAT_6[3]\, \PATT_ELK_DAT_6[4]\, 
        \PATT_ELK_DAT_6[5]\, \PATT_ELK_DAT_6[6]\, 
        \PATT_ELK_DAT_6[7]\, \ELK_RX_SER_WORD_6[0]\, 
        \ELK_RX_SER_WORD_6[1]\, \ELK_RX_SER_WORD_6[2]\, 
        \ELK_RX_SER_WORD_6[3]\, \ELK_RX_SER_WORD_6[4]\, 
        \ELK_RX_SER_WORD_6[5]\, \ELK_RX_SER_WORD_6[6]\, 
        \ELK_RX_SER_WORD_6[7]\, \PATT_ELK_DAT_7[0]\, 
        \PATT_ELK_DAT_7[1]\, \PATT_ELK_DAT_7[2]\, 
        \PATT_ELK_DAT_7[3]\, \PATT_ELK_DAT_7[4]\, 
        \PATT_ELK_DAT_7[5]\, \PATT_ELK_DAT_7[6]\, 
        \PATT_ELK_DAT_7[7]\, \ELK_RX_SER_WORD_7[0]\, 
        \ELK_RX_SER_WORD_7[1]\, \ELK_RX_SER_WORD_7[2]\, 
        \ELK_RX_SER_WORD_7[3]\, \ELK_RX_SER_WORD_7[4]\, 
        \ELK_RX_SER_WORD_7[5]\, \ELK_RX_SER_WORD_7[6]\, 
        \ELK_RX_SER_WORD_7[7]\, \PATT_ELK_DAT_8[0]\, 
        \PATT_ELK_DAT_8[1]\, \PATT_ELK_DAT_8[2]\, 
        \PATT_ELK_DAT_8[3]\, \PATT_ELK_DAT_8[4]\, 
        \PATT_ELK_DAT_8[5]\, \PATT_ELK_DAT_8[6]\, 
        \PATT_ELK_DAT_8[7]\, \ELK_RX_SER_WORD_8[0]\, 
        \ELK_RX_SER_WORD_8[1]\, \ELK_RX_SER_WORD_8[2]\, 
        \ELK_RX_SER_WORD_8[3]\, \ELK_RX_SER_WORD_8[4]\, 
        \ELK_RX_SER_WORD_8[5]\, \ELK_RX_SER_WORD_8[6]\, 
        \ELK_RX_SER_WORD_8[7]\, \PATT_ELK_DAT_9[0]\, 
        \PATT_ELK_DAT_9[1]\, \PATT_ELK_DAT_9[2]\, 
        \PATT_ELK_DAT_9[3]\, \PATT_ELK_DAT_9[4]\, 
        \PATT_ELK_DAT_9[5]\, \PATT_ELK_DAT_9[6]\, 
        \PATT_ELK_DAT_9[7]\, \ELK_RX_SER_WORD_9[0]\, 
        \ELK_RX_SER_WORD_9[1]\, \ELK_RX_SER_WORD_9[2]\, 
        \ELK_RX_SER_WORD_9[3]\, \ELK_RX_SER_WORD_9[4]\, 
        \ELK_RX_SER_WORD_9[5]\, \ELK_RX_SER_WORD_9[6]\, 
        \ELK_RX_SER_WORD_9[7]\, \PATT_ELK_DAT_10[0]\, 
        \PATT_ELK_DAT_10[1]\, \PATT_ELK_DAT_10[2]\, 
        \PATT_ELK_DAT_10[3]\, \PATT_ELK_DAT_10[4]\, 
        \PATT_ELK_DAT_10[5]\, \PATT_ELK_DAT_10[6]\, 
        \PATT_ELK_DAT_10[7]\, \ELK_RX_SER_WORD_10[0]\, 
        \ELK_RX_SER_WORD_10[1]\, \ELK_RX_SER_WORD_10[2]\, 
        \ELK_RX_SER_WORD_10[3]\, \ELK_RX_SER_WORD_10[4]\, 
        \ELK_RX_SER_WORD_10[5]\, \ELK_RX_SER_WORD_10[6]\, 
        \ELK_RX_SER_WORD_10[7]\, \PATT_ELK_DAT_11[0]\, 
        \PATT_ELK_DAT_11[1]\, \PATT_ELK_DAT_11[2]\, 
        \PATT_ELK_DAT_11[3]\, \PATT_ELK_DAT_11[4]\, 
        \PATT_ELK_DAT_11[5]\, \PATT_ELK_DAT_11[6]\, 
        \PATT_ELK_DAT_11[7]\, \ELK_RX_SER_WORD_11[0]\, 
        \ELK_RX_SER_WORD_11[1]\, \ELK_RX_SER_WORD_11[2]\, 
        \ELK_RX_SER_WORD_11[3]\, \ELK_RX_SER_WORD_11[4]\, 
        \ELK_RX_SER_WORD_11[5]\, \ELK_RX_SER_WORD_11[6]\, 
        \ELK_RX_SER_WORD_11[7]\, \PATT_ELK_DAT_12[0]\, 
        \PATT_ELK_DAT_12[1]\, \PATT_ELK_DAT_12[2]\, 
        \PATT_ELK_DAT_12[3]\, \PATT_ELK_DAT_12[4]\, 
        \PATT_ELK_DAT_12[5]\, \PATT_ELK_DAT_12[6]\, 
        \PATT_ELK_DAT_12[7]\, \ELK_RX_SER_WORD_12[0]\, 
        \ELK_RX_SER_WORD_12[1]\, \ELK_RX_SER_WORD_12[2]\, 
        \ELK_RX_SER_WORD_12[3]\, \ELK_RX_SER_WORD_12[4]\, 
        \ELK_RX_SER_WORD_12[5]\, \ELK_RX_SER_WORD_12[6]\, 
        \ELK_RX_SER_WORD_12[7]\, \PATT_ELK_DAT_13[0]\, 
        \PATT_ELK_DAT_13[1]\, \PATT_ELK_DAT_13[2]\, 
        \PATT_ELK_DAT_13[3]\, \PATT_ELK_DAT_13[4]\, 
        \PATT_ELK_DAT_13[5]\, \PATT_ELK_DAT_13[6]\, 
        \PATT_ELK_DAT_13[7]\, \ELK_RX_SER_WORD_13[0]\, 
        \ELK_RX_SER_WORD_13[1]\, \ELK_RX_SER_WORD_13[2]\, 
        \ELK_RX_SER_WORD_13[3]\, \ELK_RX_SER_WORD_13[4]\, 
        \ELK_RX_SER_WORD_13[5]\, \ELK_RX_SER_WORD_13[6]\, 
        \ELK_RX_SER_WORD_13[7]\, \PATT_ELK_DAT_14[0]\, 
        \PATT_ELK_DAT_14[1]\, \PATT_ELK_DAT_14[2]\, 
        \PATT_ELK_DAT_14[3]\, \PATT_ELK_DAT_14[4]\, 
        \PATT_ELK_DAT_14[5]\, \PATT_ELK_DAT_14[6]\, 
        \PATT_ELK_DAT_14[7]\, \ELK_RX_SER_WORD_14[0]\, 
        \ELK_RX_SER_WORD_14[1]\, \ELK_RX_SER_WORD_14[2]\, 
        \ELK_RX_SER_WORD_14[3]\, \ELK_RX_SER_WORD_14[4]\, 
        \ELK_RX_SER_WORD_14[5]\, \ELK_RX_SER_WORD_14[6]\, 
        \ELK_RX_SER_WORD_14[7]\, \PATT_ELK_DAT_15[0]\, 
        \PATT_ELK_DAT_15[1]\, \PATT_ELK_DAT_15[2]\, 
        \PATT_ELK_DAT_15[3]\, \PATT_ELK_DAT_15[4]\, 
        \PATT_ELK_DAT_15[5]\, \PATT_ELK_DAT_15[6]\, 
        \PATT_ELK_DAT_15[7]\, \ELK_RX_SER_WORD_15[0]\, 
        \ELK_RX_SER_WORD_15[1]\, \ELK_RX_SER_WORD_15[2]\, 
        \ELK_RX_SER_WORD_15[3]\, \ELK_RX_SER_WORD_15[4]\, 
        \ELK_RX_SER_WORD_15[5]\, \ELK_RX_SER_WORD_15[6]\, 
        \ELK_RX_SER_WORD_15[7]\, \PATT_ELK_DAT_16[0]\, 
        \PATT_ELK_DAT_16[1]\, \PATT_ELK_DAT_16[2]\, 
        \PATT_ELK_DAT_16[3]\, \PATT_ELK_DAT_16[4]\, 
        \PATT_ELK_DAT_16[5]\, \PATT_ELK_DAT_16[6]\, 
        \PATT_ELK_DAT_16[7]\, \ELK_RX_SER_WORD_16[0]\, 
        \ELK_RX_SER_WORD_16[1]\, \ELK_RX_SER_WORD_16[2]\, 
        \ELK_RX_SER_WORD_16[3]\, \ELK_RX_SER_WORD_16[4]\, 
        \ELK_RX_SER_WORD_16[5]\, \ELK_RX_SER_WORD_16[6]\, 
        \ELK_RX_SER_WORD_16[7]\, \PATT_ELK_DAT_17[0]\, 
        \PATT_ELK_DAT_17[1]\, \PATT_ELK_DAT_17[2]\, 
        \PATT_ELK_DAT_17[3]\, \PATT_ELK_DAT_17[4]\, 
        \PATT_ELK_DAT_17[5]\, \PATT_ELK_DAT_17[6]\, 
        \PATT_ELK_DAT_17[7]\, \ELK_RX_SER_WORD_17[0]\, 
        \ELK_RX_SER_WORD_17[1]\, \ELK_RX_SER_WORD_17[2]\, 
        \ELK_RX_SER_WORD_17[3]\, \ELK_RX_SER_WORD_17[4]\, 
        \ELK_RX_SER_WORD_17[5]\, \ELK_RX_SER_WORD_17[6]\, 
        \ELK_RX_SER_WORD_17[7]\, \PATT_ELK_DAT_18[0]\, 
        \PATT_ELK_DAT_18[1]\, \PATT_ELK_DAT_18[2]\, 
        \PATT_ELK_DAT_18[3]\, \PATT_ELK_DAT_18[4]\, 
        \PATT_ELK_DAT_18[5]\, \PATT_ELK_DAT_18[6]\, 
        \PATT_ELK_DAT_18[7]\, \ELK_RX_SER_WORD_18[0]\, 
        \ELK_RX_SER_WORD_18[1]\, \ELK_RX_SER_WORD_18[2]\, 
        \ELK_RX_SER_WORD_18[3]\, \ELK_RX_SER_WORD_18[4]\, 
        \ELK_RX_SER_WORD_18[5]\, \ELK_RX_SER_WORD_18[6]\, 
        \ELK_RX_SER_WORD_18[7]\, \PATT_ELK_DAT_19[0]\, 
        \PATT_ELK_DAT_19[1]\, \PATT_ELK_DAT_19[2]\, 
        \PATT_ELK_DAT_19[3]\, \PATT_ELK_DAT_19[4]\, 
        \PATT_ELK_DAT_19[5]\, \PATT_ELK_DAT_19[6]\, 
        \PATT_ELK_DAT_19[7]\, \ELK_RX_SER_WORD_19[0]\, 
        \ELK_RX_SER_WORD_19[1]\, \ELK_RX_SER_WORD_19[2]\, 
        \ELK_RX_SER_WORD_19[3]\, \ELK_RX_SER_WORD_19[4]\, 
        \ELK_RX_SER_WORD_19[5]\, \ELK_RX_SER_WORD_19[6]\, 
        \ELK_RX_SER_WORD_19[7]\, USB_OE_BI, USB_RD_BI, USB_WR_BI, 
        USB_SIWU_BI, \TFC_STRT_ADDR[0]\, \TFC_STRT_ADDR[1]\, 
        \TFC_STRT_ADDR[2]\, \TFC_STRT_ADDR[3]\, 
        \TFC_STRT_ADDR[4]\, \TFC_STRT_ADDR[5]\, 
        \TFC_STRT_ADDR[6]\, \TFC_STRT_ADDR[7]\, 
        \TFC_STOP_ADDR[0]\, \TFC_STOP_ADDR[1]\, 
        \TFC_STOP_ADDR[2]\, \TFC_STOP_ADDR[3]\, 
        \TFC_STOP_ADDR[4]\, \TFC_STOP_ADDR[5]\, 
        \TFC_STOP_ADDR[6]\, \TFC_STOP_ADDR[7]\, \TFC_ADDRB[0]\, 
        \TFC_ADDRB[1]\, \TFC_ADDRB[2]\, \TFC_ADDRB[3]\, 
        \TFC_ADDRB[4]\, \TFC_ADDRB[5]\, \TFC_ADDRB[6]\, 
        \TFC_ADDRB[7]\, TFC_RAM_BLKB_EN, TFC_RWB, 
        \ELKS_STRT_ADDR[0]\, \ELKS_STRT_ADDR[1]\, 
        \ELKS_STRT_ADDR[2]\, \ELKS_STRT_ADDR[3]\, 
        \ELKS_STRT_ADDR[4]\, \ELKS_STRT_ADDR[5]\, 
        \ELKS_STRT_ADDR[6]\, \ELKS_STRT_ADDR[7]\, 
        \ELKS_STOP_ADDR[0]\, \ELKS_STOP_ADDR[1]\, 
        \ELKS_STOP_ADDR[2]\, \ELKS_STOP_ADDR[3]\, 
        \ELKS_STOP_ADDR[4]\, \ELKS_STOP_ADDR[5]\, 
        \ELKS_STOP_ADDR[6]\, \ELKS_STOP_ADDR[7]\, \ELKS_ADDRB[0]\, 
        \ELKS_ADDRB[1]\, \ELKS_ADDRB[2]\, \ELKS_ADDRB[3]\, 
        \ELKS_ADDRB[4]\, \ELKS_ADDRB[5]\, \ELKS_ADDRB[6]\, 
        \ELKS_ADDRB[7]\, ELKS_RAM_BLKB_EN, ELKS_RWB, \OP_MODE[0]\, 
        \OP_MODE[4]\, \SYNC_STAT_DET.ELK0_SYNC_DET_1\, 
        \SYNC_STAT_DET.TFC_SYNC_DET_1\, DEV_RST_B_c, 
        DCB_SALT_SEL_c, EXTCLK_40MHZ_c, EXT_INT_REF_SEL_c, 
        ALL_PLL_LOCK_c, P_MASTER_POR_B_c, P_USB_MASTER_EN_c, 
        CLK_40M_GL, CCC_160M_FXD, CCC_160M_ADJ, P_ELK0_SYNC_DET_c, 
        P_TFC_SYNC_DET_c, \OP_MODE_c[1]\, \OP_MODE_c[2]\, 
        \OP_MODE_c[5]\, \OP_MODE_c[6]\, USBCLK60MHZ_c, 
        P_USB_RXF_B_c, P_USB_TXE_B_c, ELK0_OUT_R_i_0, 
        ELK0_OUT_F_i_0, MASTER_DCB_POR_B_i_0_i, 
        MASTER_SALT_POR_B_i_0_i, DCB_SALT_SEL_c_i, 
        ELK0_IN_DDR_F_i, ELK0_IN_DDR_R_i, 
        MASTER_SALT_POR_B_i_0_i_0, MASTER_SALT_POR_B_i_0_i_1, 
        MASTER_SALT_POR_B_i_0_i_2, MASTER_SALT_POR_B_i_0_i_3, 
        MASTER_SALT_POR_B_i_0_i_4, MASTER_SALT_POR_B_i_0_i_5, 
        MASTER_SALT_POR_B_i_0_i_6, MASTER_SALT_POR_B_i_0_i_7, 
        MASTER_SALT_POR_B_i_0_i_8, MASTER_SALT_POR_B_i_0_i_9, 
        MASTER_SALT_POR_B_i_0_i_10, MASTER_SALT_POR_B_i_0_i_11, 
        MASTER_SALT_POR_B_i_0_i_12, MASTER_SALT_POR_B_i_0_i_13, 
        MASTER_SALT_POR_B_i_0_i_14, MASTER_SALT_POR_B_i_0_i_15, 
        MASTER_SALT_POR_B_i_0_i_16, MASTER_SALT_POR_B_i_0_i_17, 
        \OP_MODE_c_0[1]\, \OP_MODE_c_1[1]\, \OP_MODE_c_2[1]\, 
        \OP_MODE_c_3[1]\, \OP_MODE_c_4[1]\, \OP_MODE_c_5[1]\, 
        \OP_MODE_c_6[1]\, P_USB_MASTER_EN_c_0, 
        P_USB_MASTER_EN_c_1, P_USB_MASTER_EN_c_2, 
        P_USB_MASTER_EN_c_3, P_USB_MASTER_EN_c_4, 
        P_USB_MASTER_EN_c_5, P_USB_MASTER_EN_c_6, 
        P_USB_MASTER_EN_c_7, P_USB_MASTER_EN_c_8, 
        P_USB_MASTER_EN_c_9, P_USB_MASTER_EN_c_10, 
        P_USB_MASTER_EN_c_11, P_USB_MASTER_EN_c_12, 
        P_USB_MASTER_EN_c_13, P_USB_MASTER_EN_c_14, 
        P_USB_MASTER_EN_c_15, P_USB_MASTER_EN_c_16, 
        P_USB_MASTER_EN_c_17, P_USB_MASTER_EN_c_18, 
        P_USB_MASTER_EN_c_19, P_USB_MASTER_EN_c_20, 
        P_USB_MASTER_EN_c_21, P_USB_MASTER_EN_c_22, 
        P_MASTER_POR_B_c_1, P_MASTER_POR_B_c_2, 
        P_MASTER_POR_B_c_3, P_MASTER_POR_B_c_4, 
        P_MASTER_POR_B_c_5, P_MASTER_POR_B_c_6, 
        P_MASTER_POR_B_c_7, P_MASTER_POR_B_c_8, 
        P_MASTER_POR_B_c_9, P_MASTER_POR_B_c_10, 
        P_MASTER_POR_B_c_11, P_MASTER_POR_B_c_12, 
        P_MASTER_POR_B_c_13, P_MASTER_POR_B_c_14, 
        P_MASTER_POR_B_c_15, P_MASTER_POR_B_c_16, 
        P_MASTER_POR_B_c_17, P_MASTER_POR_B_c_18, 
        P_MASTER_POR_B_c_19, P_MASTER_POR_B_c_20, 
        P_MASTER_POR_B_c_21, P_MASTER_POR_B_c_22, 
        P_MASTER_POR_B_c_23, P_MASTER_POR_B_c_24, 
        P_MASTER_POR_B_c_25, P_MASTER_POR_B_c_26, 
        P_MASTER_POR_B_c_27, P_MASTER_POR_B_c_28, 
        P_MASTER_POR_B_c_29, P_MASTER_POR_B_c_30, 
        P_MASTER_POR_B_c_31, P_MASTER_POR_B_c_32, 
        P_MASTER_POR_B_c_33, P_MASTER_POR_B_c_34, DEV_RST_B_c_0, 
        DEV_RST_B_c_1, \ELKS_ADDRB_0[6]\, \ELKS_ADDRB_0[4]\, 
        \ELKS_ADDRB_0[2]\, \BIT_OS_SEL_0[2]\, \BIT_OS_SEL_1[2]\, 
        \BIT_OS_SEL_2[2]\, \BIT_OS_SEL_3[2]\, \BIT_OS_SEL_4[2]\, 
        \BIT_OS_SEL_5[2]\, \BIT_OS_SEL_6[2]\, \BIT_OS_SEL_7[2]\, 
        \BIT_OS_SEL_0[1]\, \BIT_OS_SEL_1[1]\, \BIT_OS_SEL_2[1]\, 
        \BIT_OS_SEL_3[1]\, \BIT_OS_SEL_4[1]\, \BIT_OS_SEL_5[1]\, 
        \BIT_OS_SEL_6[1]\, \BIT_OS_SEL_0[0]\, \BIT_OS_SEL_1[0]\, 
        \BIT_OS_SEL_2[0]\, \BIT_OS_SEL_3[0]\, \BIT_OS_SEL_4[0]\, 
        \BIT_OS_SEL_5[0]\, P_MASTER_POR_B_c_34_0, 
        P_MASTER_POR_B_c_32_0, P_MASTER_POR_B_c_31_0, 
        P_MASTER_POR_B_c_27_0, P_MASTER_POR_B_c_27_1, 
        P_MASTER_POR_B_c_24_0, P_MASTER_POR_B_c_22_0, 
        P_MASTER_POR_B_c_17_0, P_MASTER_POR_B_c_16_0, 
        P_USB_MASTER_EN_c_22_0, P_USB_MASTER_EN_c_2_0, 
        P_USB_MASTER_EN_c_1_0, P_MASTER_POR_B_c_0_0 : std_logic;

    for all : ELINK_SLAVE_INV_2
	Use entity work.ELINK_SLAVE_INV_2(DEF_ARCH);
    for all : ELINK_SLAVE_INV_2_0
	Use entity work.ELINK_SLAVE_INV_2_0(DEF_ARCH);
    for all : USB_INTERFACE
	Use entity work.USB_INTERFACE(DEF_ARCH);
    for all : SYNC_DAT_SEL
	Use entity work.SYNC_DAT_SEL(DEF_ARCH);
    for all : CLK_FXD_40_160_A60M
	Use entity work.CLK_FXD_40_160_A60M(DEF_ARCH);
    for all : ELINK_SLAVE_15_13
	Use entity work.ELINK_SLAVE_15_13(DEF_ARCH);
    for all : tristate_buf_1
	Use entity work.tristate_buf_1(DEF_ARCH);
    for all : BIDIR_LVDS_IO_0
	Use entity work.BIDIR_LVDS_IO_0(DEF_ARCH);
    for all : ELINK_SLAVE_15_6
	Use entity work.ELINK_SLAVE_15_6(DEF_ARCH);
    for all : GP_PATT_GEN_1_0
	Use entity work.GP_PATT_GEN_1_0(DEF_ARCH);
    for all : SER320M_3_34
	Use entity work.SER320M_3_34(DEF_ARCH);
    for all : SER320M_3_34_0
	Use entity work.SER320M_3_34_0(DEF_ARCH);
    for all : ELINK_SLAVE_15_7
	Use entity work.ELINK_SLAVE_15_7(DEF_ARCH);
    for all : ELINK_SLAVE_15_8
	Use entity work.ELINK_SLAVE_15_8(DEF_ARCH);
    for all : SYNC_DAT_SEL_0
	Use entity work.SYNC_DAT_SEL_0(DEF_ARCH);
    for all : EXEC_MODE_CNTL
	Use entity work.EXEC_MODE_CNTL(DEF_ARCH);
    for all : ELINK_SLAVE_15_2
	Use entity work.ELINK_SLAVE_15_2(DEF_ARCH);
    for all : ELINK_SLAVE_15_9
	Use entity work.ELINK_SLAVE_15_9(DEF_ARCH);
    for all : tristate_buf_0
	Use entity work.tristate_buf_0(DEF_ARCH);
    for all : ELINK_SLAVE_15
	Use entity work.ELINK_SLAVE_15(DEF_ARCH);
    for all : ELINK_SLAVE_INV_2_1
	Use entity work.ELINK_SLAVE_INV_2_1(DEF_ARCH);
    for all : DDR_BIDIR_LVDS_DUAL_CLK
	Use entity work.DDR_BIDIR_LVDS_DUAL_CLK(DEF_ARCH);
    for all : tristate_buf
	Use entity work.tristate_buf(DEF_ARCH);
    for all : REF_CLK_DIV_GEN
	Use entity work.REF_CLK_DIV_GEN(DEF_ARCH);
    for all : ELINK_SLAVE_15_1
	Use entity work.ELINK_SLAVE_15_1(DEF_ARCH);
    for all : TOP_MASTER_DES320M
	Use entity work.TOP_MASTER_DES320M(DEF_ARCH);
    for all : ELINK_SLAVE_15_11
	Use entity work.ELINK_SLAVE_15_11(DEF_ARCH);
    for all : tristate_buf_2
	Use entity work.tristate_buf_2(DEF_ARCH);
    for all : DDR_BIDIR_LVDS_DUAL_CLK_0
	Use entity work.DDR_BIDIR_LVDS_DUAL_CLK_0(DEF_ARCH);
    for all : LVDS_CLK_IN
	Use entity work.LVDS_CLK_IN(DEF_ARCH);
    for all : ELINK_SLAVE_15_14
	Use entity work.ELINK_SLAVE_15_14(DEF_ARCH);
    for all : ELINK_SLAVE_15_4
	Use entity work.ELINK_SLAVE_15_4(DEF_ARCH);
    for all : GP_PATT_GEN_1
	Use entity work.GP_PATT_GEN_1(DEF_ARCH);
    for all : ELINK_SLAVE_15_3
	Use entity work.ELINK_SLAVE_15_3(DEF_ARCH);
    for all : ELINK_SLAVE_15_12
	Use entity work.ELINK_SLAVE_15_12(DEF_ARCH);
    for all : ELINK_SLAVE_15_10
	Use entity work.ELINK_SLAVE_15_10(DEF_ARCH);
    for all : BIDIR_LVDS_IO
	Use entity work.BIDIR_LVDS_IO(DEF_ARCH);
    for all : LVDS_BUFOUT
	Use entity work.LVDS_BUFOUT(DEF_ARCH);
    for all : ELINK_SLAVE_15_0
	Use entity work.ELINK_SLAVE_15_0(DEF_ARCH);
    for all : ELINK_SLAVE_15_5
	Use entity work.ELINK_SLAVE_15_5(DEF_ARCH);
begin 


    TFC_SYNC_DET : DFN1C0
      port map(D => \SYNC_STAT_DET.TFC_SYNC_DET_1\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_23, Q => 
        P_TFC_SYNC_DET_c);
    
    DEV_RST_B_pad : INBUF
      port map(PAD => DEV_RST_B, Y => DEV_RST_B_c);
    
    U_ELK1_CH : ELINK_SLAVE_INV_2
      port map(BIT_OS_SEL_0_d0 => \BIT_OS_SEL[2]\, BIT_OS_SEL_0_0
         => \BIT_OS_SEL_0[1]\, BIT_OS_SEL_1(2) => 
        \BIT_OS_SEL_1[2]\, BIT_OS_SEL_1(1) => \BIT_OS_SEL_1[1]\, 
        BIT_OS_SEL_1(0) => \BIT_OS_SEL_1[0]\, BIT_OS_SEL_2_0 => 
        \BIT_OS_SEL_2[0]\, ELK_RX_SER_WORD_1(7) => 
        \ELK_RX_SER_WORD_1[7]\, ELK_RX_SER_WORD_1(6) => 
        \ELK_RX_SER_WORD_1[6]\, ELK_RX_SER_WORD_1(5) => 
        \ELK_RX_SER_WORD_1[5]\, ELK_RX_SER_WORD_1(4) => 
        \ELK_RX_SER_WORD_1[4]\, ELK_RX_SER_WORD_1(3) => 
        \ELK_RX_SER_WORD_1[3]\, ELK_RX_SER_WORD_1(2) => 
        \ELK_RX_SER_WORD_1[2]\, ELK_RX_SER_WORD_1(1) => 
        \ELK_RX_SER_WORD_1[1]\, ELK_RX_SER_WORD_1(0) => 
        \ELK_RX_SER_WORD_1[0]\, OP_MODE_c_5_0 => \OP_MODE_c_5[1]\, 
        PATT_ELK_DAT_1(7) => \PATT_ELK_DAT_1[7]\, 
        PATT_ELK_DAT_1(6) => \PATT_ELK_DAT_1[6]\, 
        PATT_ELK_DAT_1(5) => \PATT_ELK_DAT_1[5]\, 
        PATT_ELK_DAT_1(4) => \PATT_ELK_DAT_1[4]\, 
        PATT_ELK_DAT_1(3) => \PATT_ELK_DAT_1[3]\, 
        PATT_ELK_DAT_1(2) => \PATT_ELK_DAT_1[2]\, 
        PATT_ELK_DAT_1(1) => \PATT_ELK_DAT_1[1]\, 
        PATT_ELK_DAT_1(0) => \PATT_ELK_DAT_1[0]\, 
        MASTER_DCB_POR_B_i_0_i => MASTER_DCB_POR_B_i_0_i, 
        ELK1_DAT_N => ELK1_DAT_N, ELK1_DAT_P => ELK1_DAT_P, 
        DCB_SALT_SEL_c_i => DCB_SALT_SEL_c_i, CCC_160M_FXD => 
        CCC_160M_FXD, MASTER_SALT_POR_B_i_0_i_14 => 
        MASTER_SALT_POR_B_i_0_i_14, MASTER_SALT_POR_B_i_0_i_7 => 
        MASTER_SALT_POR_B_i_0_i_7, MASTER_SALT_POR_B_i_0_i_1 => 
        MASTER_SALT_POR_B_i_0_i_1, MASTER_SALT_POR_B_i_0_i_16 => 
        MASTER_SALT_POR_B_i_0_i_16, MASTER_SALT_POR_B_i_0_i_4 => 
        MASTER_SALT_POR_B_i_0_i_4, CLK_40M_GL => CLK_40M_GL, 
        MASTER_SALT_POR_B_i_0_i_11 => MASTER_SALT_POR_B_i_0_i_11, 
        DEV_RST_B_c_0 => DEV_RST_B_c_0, CCC_160M_ADJ => 
        CCC_160M_ADJ);
    
    P_CCC_160M_ADJ_pad : OUTBUF
      port map(D => CCC_160M_ADJ, PAD => P_CCC_160M_ADJ);
    
    USBCLK60MHZ_pad : INBUF
      port map(PAD => USBCLK60MHZ, Y => USBCLK60MHZ_c);
    
    P_USB_RXF_B_pad : INBUF
      port map(PAD => P_USB_RXF_B, Y => P_USB_RXF_B_c);
    
    U_ELK3_CH : ELINK_SLAVE_INV_2_0
      port map(BIT_OS_SEL_7_0 => \BIT_OS_SEL_7[2]\, 
        BIT_OS_SEL_6_0 => \BIT_OS_SEL_6[1]\, BIT_OS_SEL_0_d0 => 
        \BIT_OS_SEL[1]\, BIT_OS_SEL_0(2) => \BIT_OS_SEL_0[2]\, 
        BIT_OS_SEL_0(1) => \BIT_OS_SEL_0[1]\, BIT_OS_SEL_1_0 => 
        \BIT_OS_SEL_1[0]\, ELK_RX_SER_WORD_3(7) => 
        \ELK_RX_SER_WORD_3[7]\, ELK_RX_SER_WORD_3(6) => 
        \ELK_RX_SER_WORD_3[6]\, ELK_RX_SER_WORD_3(5) => 
        \ELK_RX_SER_WORD_3[5]\, ELK_RX_SER_WORD_3(4) => 
        \ELK_RX_SER_WORD_3[4]\, ELK_RX_SER_WORD_3(3) => 
        \ELK_RX_SER_WORD_3[3]\, ELK_RX_SER_WORD_3(2) => 
        \ELK_RX_SER_WORD_3[2]\, ELK_RX_SER_WORD_3(1) => 
        \ELK_RX_SER_WORD_3[1]\, ELK_RX_SER_WORD_3(0) => 
        \ELK_RX_SER_WORD_3[0]\, OP_MODE_c_5_0 => \OP_MODE_c_5[1]\, 
        PATT_ELK_DAT_3(7) => \PATT_ELK_DAT_3[7]\, 
        PATT_ELK_DAT_3(6) => \PATT_ELK_DAT_3[6]\, 
        PATT_ELK_DAT_3(5) => \PATT_ELK_DAT_3[5]\, 
        PATT_ELK_DAT_3(4) => \PATT_ELK_DAT_3[4]\, 
        PATT_ELK_DAT_3(3) => \PATT_ELK_DAT_3[3]\, 
        PATT_ELK_DAT_3(2) => \PATT_ELK_DAT_3[2]\, 
        PATT_ELK_DAT_3(1) => \PATT_ELK_DAT_3[1]\, 
        PATT_ELK_DAT_3(0) => \PATT_ELK_DAT_3[0]\, 
        MASTER_DCB_POR_B_i_0_i => MASTER_DCB_POR_B_i_0_i, 
        ELK3_DAT_N => ELK3_DAT_N, ELK3_DAT_P => ELK3_DAT_P, 
        DCB_SALT_SEL_c_i => DCB_SALT_SEL_c_i, CCC_160M_FXD => 
        CCC_160M_FXD, MASTER_SALT_POR_B_i_0_i_8 => 
        MASTER_SALT_POR_B_i_0_i_8, MASTER_SALT_POR_B_i_0_i_5 => 
        MASTER_SALT_POR_B_i_0_i_5, MASTER_SALT_POR_B_i_0_i_2 => 
        MASTER_SALT_POR_B_i_0_i_2, MASTER_SALT_POR_B_i_0_i_3 => 
        MASTER_SALT_POR_B_i_0_i_3, MASTER_SALT_POR_B_i_0_i_16 => 
        MASTER_SALT_POR_B_i_0_i_16, MASTER_SALT_POR_B_i_0_i_12
         => MASTER_SALT_POR_B_i_0_i_12, CLK_40M_GL => CLK_40M_GL, 
        MASTER_SALT_POR_B_i_0_i_14 => MASTER_SALT_POR_B_i_0_i_14, 
        MASTER_SALT_POR_B_i_0_i_15 => MASTER_SALT_POR_B_i_0_i_15, 
        DEV_RST_B_c => DEV_RST_B_c, CCC_160M_ADJ => CCC_160M_ADJ);
    
    U50_PATTERNS : USB_INTERFACE
      port map(OP_MODE_c_6_0 => \OP_MODE_c_6[1]\, OP_MODE_c_5_0
         => \OP_MODE_c_5[1]\, OP_MODE_c_4_0 => \OP_MODE_c_4[1]\, 
        OP_MODE_c_3_0 => \OP_MODE_c_3[1]\, OP_MODE_c_2_0 => 
        \OP_MODE_c_2[1]\, OP_MODE_c_1_0 => \OP_MODE_c_1[1]\, 
        OP_MODE_c_0_0 => \OP_MODE_c_0[1]\, OP_MODE_c_1_d0 => 
        \OP_MODE_c[2]\, OP_MODE_c_5_d0 => \OP_MODE_c[6]\, 
        OP_MODE_c_4_d0 => \OP_MODE_c[5]\, OP_MODE_c_0_d0 => 
        \OP_MODE_c[1]\, OP_MODE_0_0 => \OP_MODE[0]\, OP_MODE_0_4
         => \OP_MODE[4]\, ELKS_STOP_ADDR(7) => 
        \ELKS_STOP_ADDR[7]\, ELKS_STOP_ADDR(6) => 
        \ELKS_STOP_ADDR[6]\, ELKS_STOP_ADDR(5) => 
        \ELKS_STOP_ADDR[5]\, ELKS_STOP_ADDR(4) => 
        \ELKS_STOP_ADDR[4]\, ELKS_STOP_ADDR(3) => 
        \ELKS_STOP_ADDR[3]\, ELKS_STOP_ADDR(2) => 
        \ELKS_STOP_ADDR[2]\, ELKS_STOP_ADDR(1) => 
        \ELKS_STOP_ADDR[1]\, ELKS_STOP_ADDR(0) => 
        \ELKS_STOP_ADDR[0]\, ELKS_STRT_ADDR(7) => 
        \ELKS_STRT_ADDR[7]\, ELKS_STRT_ADDR(6) => 
        \ELKS_STRT_ADDR[6]\, ELKS_STRT_ADDR(5) => 
        \ELKS_STRT_ADDR[5]\, ELKS_STRT_ADDR(4) => 
        \ELKS_STRT_ADDR[4]\, ELKS_STRT_ADDR(3) => 
        \ELKS_STRT_ADDR[3]\, ELKS_STRT_ADDR(2) => 
        \ELKS_STRT_ADDR[2]\, ELKS_STRT_ADDR(1) => 
        \ELKS_STRT_ADDR[1]\, ELKS_STRT_ADDR(0) => 
        \ELKS_STRT_ADDR[0]\, TFC_STOP_ADDR_0(7) => 
        \TFC_STOP_ADDR[7]\, TFC_STOP_ADDR_0(6) => 
        \TFC_STOP_ADDR[6]\, TFC_STOP_ADDR_0(5) => 
        \TFC_STOP_ADDR[5]\, TFC_STOP_ADDR_0(4) => 
        \TFC_STOP_ADDR[4]\, TFC_STOP_ADDR_0(3) => 
        \TFC_STOP_ADDR[3]\, TFC_STOP_ADDR_0(2) => 
        \TFC_STOP_ADDR[2]\, TFC_STOP_ADDR_0(1) => 
        \TFC_STOP_ADDR[1]\, TFC_STOP_ADDR_0(0) => 
        \TFC_STOP_ADDR[0]\, TFC_STRT_ADDR_0(7) => 
        \TFC_STRT_ADDR[7]\, TFC_STRT_ADDR_0(6) => 
        \TFC_STRT_ADDR[6]\, TFC_STRT_ADDR_0(5) => 
        \TFC_STRT_ADDR[5]\, TFC_STRT_ADDR_0(4) => 
        \TFC_STRT_ADDR[4]\, TFC_STRT_ADDR_0(3) => 
        \TFC_STRT_ADDR[3]\, TFC_STRT_ADDR_0(2) => 
        \TFC_STRT_ADDR[2]\, TFC_STRT_ADDR_0(1) => 
        \TFC_STRT_ADDR[1]\, TFC_STRT_ADDR_0(0) => 
        \TFC_STRT_ADDR[0]\, BIDIR_USB_ADBUS(7) => 
        BIDIR_USB_ADBUS(7), BIDIR_USB_ADBUS(6) => 
        BIDIR_USB_ADBUS(6), BIDIR_USB_ADBUS(5) => 
        BIDIR_USB_ADBUS(5), BIDIR_USB_ADBUS(4) => 
        BIDIR_USB_ADBUS(4), BIDIR_USB_ADBUS(3) => 
        BIDIR_USB_ADBUS(3), BIDIR_USB_ADBUS(2) => 
        BIDIR_USB_ADBUS(2), BIDIR_USB_ADBUS(1) => 
        BIDIR_USB_ADBUS(1), BIDIR_USB_ADBUS(0) => 
        BIDIR_USB_ADBUS(0), PATT_ELK_DAT_19(7) => 
        \PATT_ELK_DAT_19[7]\, PATT_ELK_DAT_19(6) => 
        \PATT_ELK_DAT_19[6]\, PATT_ELK_DAT_19(5) => 
        \PATT_ELK_DAT_19[5]\, PATT_ELK_DAT_19(4) => 
        \PATT_ELK_DAT_19[4]\, PATT_ELK_DAT_19(3) => 
        \PATT_ELK_DAT_19[3]\, PATT_ELK_DAT_19(2) => 
        \PATT_ELK_DAT_19[2]\, PATT_ELK_DAT_19(1) => 
        \PATT_ELK_DAT_19[1]\, PATT_ELK_DAT_19(0) => 
        \PATT_ELK_DAT_19[0]\, ELK_RX_SER_WORD_19(7) => 
        \ELK_RX_SER_WORD_19[7]\, ELK_RX_SER_WORD_19(6) => 
        \ELK_RX_SER_WORD_19[6]\, ELK_RX_SER_WORD_19(5) => 
        \ELK_RX_SER_WORD_19[5]\, ELK_RX_SER_WORD_19(4) => 
        \ELK_RX_SER_WORD_19[4]\, ELK_RX_SER_WORD_19(3) => 
        \ELK_RX_SER_WORD_19[3]\, ELK_RX_SER_WORD_19(2) => 
        \ELK_RX_SER_WORD_19[2]\, ELK_RX_SER_WORD_19(1) => 
        \ELK_RX_SER_WORD_19[1]\, ELK_RX_SER_WORD_19(0) => 
        \ELK_RX_SER_WORD_19[0]\, PATT_ELK_DAT_18(7) => 
        \PATT_ELK_DAT_18[7]\, PATT_ELK_DAT_18(6) => 
        \PATT_ELK_DAT_18[6]\, PATT_ELK_DAT_18(5) => 
        \PATT_ELK_DAT_18[5]\, PATT_ELK_DAT_18(4) => 
        \PATT_ELK_DAT_18[4]\, PATT_ELK_DAT_18(3) => 
        \PATT_ELK_DAT_18[3]\, PATT_ELK_DAT_18(2) => 
        \PATT_ELK_DAT_18[2]\, PATT_ELK_DAT_18(1) => 
        \PATT_ELK_DAT_18[1]\, PATT_ELK_DAT_18(0) => 
        \PATT_ELK_DAT_18[0]\, ELK_RX_SER_WORD_18(7) => 
        \ELK_RX_SER_WORD_18[7]\, ELK_RX_SER_WORD_18(6) => 
        \ELK_RX_SER_WORD_18[6]\, ELK_RX_SER_WORD_18(5) => 
        \ELK_RX_SER_WORD_18[5]\, ELK_RX_SER_WORD_18(4) => 
        \ELK_RX_SER_WORD_18[4]\, ELK_RX_SER_WORD_18(3) => 
        \ELK_RX_SER_WORD_18[3]\, ELK_RX_SER_WORD_18(2) => 
        \ELK_RX_SER_WORD_18[2]\, ELK_RX_SER_WORD_18(1) => 
        \ELK_RX_SER_WORD_18[1]\, ELK_RX_SER_WORD_18(0) => 
        \ELK_RX_SER_WORD_18[0]\, PATT_ELK_DAT_17(7) => 
        \PATT_ELK_DAT_17[7]\, PATT_ELK_DAT_17(6) => 
        \PATT_ELK_DAT_17[6]\, PATT_ELK_DAT_17(5) => 
        \PATT_ELK_DAT_17[5]\, PATT_ELK_DAT_17(4) => 
        \PATT_ELK_DAT_17[4]\, PATT_ELK_DAT_17(3) => 
        \PATT_ELK_DAT_17[3]\, PATT_ELK_DAT_17(2) => 
        \PATT_ELK_DAT_17[2]\, PATT_ELK_DAT_17(1) => 
        \PATT_ELK_DAT_17[1]\, PATT_ELK_DAT_17(0) => 
        \PATT_ELK_DAT_17[0]\, ELK_RX_SER_WORD_17(7) => 
        \ELK_RX_SER_WORD_17[7]\, ELK_RX_SER_WORD_17(6) => 
        \ELK_RX_SER_WORD_17[6]\, ELK_RX_SER_WORD_17(5) => 
        \ELK_RX_SER_WORD_17[5]\, ELK_RX_SER_WORD_17(4) => 
        \ELK_RX_SER_WORD_17[4]\, ELK_RX_SER_WORD_17(3) => 
        \ELK_RX_SER_WORD_17[3]\, ELK_RX_SER_WORD_17(2) => 
        \ELK_RX_SER_WORD_17[2]\, ELK_RX_SER_WORD_17(1) => 
        \ELK_RX_SER_WORD_17[1]\, ELK_RX_SER_WORD_17(0) => 
        \ELK_RX_SER_WORD_17[0]\, PATT_ELK_DAT_16(7) => 
        \PATT_ELK_DAT_16[7]\, PATT_ELK_DAT_16(6) => 
        \PATT_ELK_DAT_16[6]\, PATT_ELK_DAT_16(5) => 
        \PATT_ELK_DAT_16[5]\, PATT_ELK_DAT_16(4) => 
        \PATT_ELK_DAT_16[4]\, PATT_ELK_DAT_16(3) => 
        \PATT_ELK_DAT_16[3]\, PATT_ELK_DAT_16(2) => 
        \PATT_ELK_DAT_16[2]\, PATT_ELK_DAT_16(1) => 
        \PATT_ELK_DAT_16[1]\, PATT_ELK_DAT_16(0) => 
        \PATT_ELK_DAT_16[0]\, ELK_RX_SER_WORD_16(7) => 
        \ELK_RX_SER_WORD_16[7]\, ELK_RX_SER_WORD_16(6) => 
        \ELK_RX_SER_WORD_16[6]\, ELK_RX_SER_WORD_16(5) => 
        \ELK_RX_SER_WORD_16[5]\, ELK_RX_SER_WORD_16(4) => 
        \ELK_RX_SER_WORD_16[4]\, ELK_RX_SER_WORD_16(3) => 
        \ELK_RX_SER_WORD_16[3]\, ELK_RX_SER_WORD_16(2) => 
        \ELK_RX_SER_WORD_16[2]\, ELK_RX_SER_WORD_16(1) => 
        \ELK_RX_SER_WORD_16[1]\, ELK_RX_SER_WORD_16(0) => 
        \ELK_RX_SER_WORD_16[0]\, PATT_ELK_DAT_15(7) => 
        \PATT_ELK_DAT_15[7]\, PATT_ELK_DAT_15(6) => 
        \PATT_ELK_DAT_15[6]\, PATT_ELK_DAT_15(5) => 
        \PATT_ELK_DAT_15[5]\, PATT_ELK_DAT_15(4) => 
        \PATT_ELK_DAT_15[4]\, PATT_ELK_DAT_15(3) => 
        \PATT_ELK_DAT_15[3]\, PATT_ELK_DAT_15(2) => 
        \PATT_ELK_DAT_15[2]\, PATT_ELK_DAT_15(1) => 
        \PATT_ELK_DAT_15[1]\, PATT_ELK_DAT_15(0) => 
        \PATT_ELK_DAT_15[0]\, ELK_RX_SER_WORD_15(7) => 
        \ELK_RX_SER_WORD_15[7]\, ELK_RX_SER_WORD_15(6) => 
        \ELK_RX_SER_WORD_15[6]\, ELK_RX_SER_WORD_15(5) => 
        \ELK_RX_SER_WORD_15[5]\, ELK_RX_SER_WORD_15(4) => 
        \ELK_RX_SER_WORD_15[4]\, ELK_RX_SER_WORD_15(3) => 
        \ELK_RX_SER_WORD_15[3]\, ELK_RX_SER_WORD_15(2) => 
        \ELK_RX_SER_WORD_15[2]\, ELK_RX_SER_WORD_15(1) => 
        \ELK_RX_SER_WORD_15[1]\, ELK_RX_SER_WORD_15(0) => 
        \ELK_RX_SER_WORD_15[0]\, PATT_ELK_DAT_14(7) => 
        \PATT_ELK_DAT_14[7]\, PATT_ELK_DAT_14(6) => 
        \PATT_ELK_DAT_14[6]\, PATT_ELK_DAT_14(5) => 
        \PATT_ELK_DAT_14[5]\, PATT_ELK_DAT_14(4) => 
        \PATT_ELK_DAT_14[4]\, PATT_ELK_DAT_14(3) => 
        \PATT_ELK_DAT_14[3]\, PATT_ELK_DAT_14(2) => 
        \PATT_ELK_DAT_14[2]\, PATT_ELK_DAT_14(1) => 
        \PATT_ELK_DAT_14[1]\, PATT_ELK_DAT_14(0) => 
        \PATT_ELK_DAT_14[0]\, ELK_RX_SER_WORD_14(7) => 
        \ELK_RX_SER_WORD_14[7]\, ELK_RX_SER_WORD_14(6) => 
        \ELK_RX_SER_WORD_14[6]\, ELK_RX_SER_WORD_14(5) => 
        \ELK_RX_SER_WORD_14[5]\, ELK_RX_SER_WORD_14(4) => 
        \ELK_RX_SER_WORD_14[4]\, ELK_RX_SER_WORD_14(3) => 
        \ELK_RX_SER_WORD_14[3]\, ELK_RX_SER_WORD_14(2) => 
        \ELK_RX_SER_WORD_14[2]\, ELK_RX_SER_WORD_14(1) => 
        \ELK_RX_SER_WORD_14[1]\, ELK_RX_SER_WORD_14(0) => 
        \ELK_RX_SER_WORD_14[0]\, PATT_ELK_DAT_13(7) => 
        \PATT_ELK_DAT_13[7]\, PATT_ELK_DAT_13(6) => 
        \PATT_ELK_DAT_13[6]\, PATT_ELK_DAT_13(5) => 
        \PATT_ELK_DAT_13[5]\, PATT_ELK_DAT_13(4) => 
        \PATT_ELK_DAT_13[4]\, PATT_ELK_DAT_13(3) => 
        \PATT_ELK_DAT_13[3]\, PATT_ELK_DAT_13(2) => 
        \PATT_ELK_DAT_13[2]\, PATT_ELK_DAT_13(1) => 
        \PATT_ELK_DAT_13[1]\, PATT_ELK_DAT_13(0) => 
        \PATT_ELK_DAT_13[0]\, ELK_RX_SER_WORD_13(7) => 
        \ELK_RX_SER_WORD_13[7]\, ELK_RX_SER_WORD_13(6) => 
        \ELK_RX_SER_WORD_13[6]\, ELK_RX_SER_WORD_13(5) => 
        \ELK_RX_SER_WORD_13[5]\, ELK_RX_SER_WORD_13(4) => 
        \ELK_RX_SER_WORD_13[4]\, ELK_RX_SER_WORD_13(3) => 
        \ELK_RX_SER_WORD_13[3]\, ELK_RX_SER_WORD_13(2) => 
        \ELK_RX_SER_WORD_13[2]\, ELK_RX_SER_WORD_13(1) => 
        \ELK_RX_SER_WORD_13[1]\, ELK_RX_SER_WORD_13(0) => 
        \ELK_RX_SER_WORD_13[0]\, PATT_ELK_DAT_12(7) => 
        \PATT_ELK_DAT_12[7]\, PATT_ELK_DAT_12(6) => 
        \PATT_ELK_DAT_12[6]\, PATT_ELK_DAT_12(5) => 
        \PATT_ELK_DAT_12[5]\, PATT_ELK_DAT_12(4) => 
        \PATT_ELK_DAT_12[4]\, PATT_ELK_DAT_12(3) => 
        \PATT_ELK_DAT_12[3]\, PATT_ELK_DAT_12(2) => 
        \PATT_ELK_DAT_12[2]\, PATT_ELK_DAT_12(1) => 
        \PATT_ELK_DAT_12[1]\, PATT_ELK_DAT_12(0) => 
        \PATT_ELK_DAT_12[0]\, ELK_RX_SER_WORD_12(7) => 
        \ELK_RX_SER_WORD_12[7]\, ELK_RX_SER_WORD_12(6) => 
        \ELK_RX_SER_WORD_12[6]\, ELK_RX_SER_WORD_12(5) => 
        \ELK_RX_SER_WORD_12[5]\, ELK_RX_SER_WORD_12(4) => 
        \ELK_RX_SER_WORD_12[4]\, ELK_RX_SER_WORD_12(3) => 
        \ELK_RX_SER_WORD_12[3]\, ELK_RX_SER_WORD_12(2) => 
        \ELK_RX_SER_WORD_12[2]\, ELK_RX_SER_WORD_12(1) => 
        \ELK_RX_SER_WORD_12[1]\, ELK_RX_SER_WORD_12(0) => 
        \ELK_RX_SER_WORD_12[0]\, PATT_ELK_DAT_11(7) => 
        \PATT_ELK_DAT_11[7]\, PATT_ELK_DAT_11(6) => 
        \PATT_ELK_DAT_11[6]\, PATT_ELK_DAT_11(5) => 
        \PATT_ELK_DAT_11[5]\, PATT_ELK_DAT_11(4) => 
        \PATT_ELK_DAT_11[4]\, PATT_ELK_DAT_11(3) => 
        \PATT_ELK_DAT_11[3]\, PATT_ELK_DAT_11(2) => 
        \PATT_ELK_DAT_11[2]\, PATT_ELK_DAT_11(1) => 
        \PATT_ELK_DAT_11[1]\, PATT_ELK_DAT_11(0) => 
        \PATT_ELK_DAT_11[0]\, ELK_RX_SER_WORD_11(7) => 
        \ELK_RX_SER_WORD_11[7]\, ELK_RX_SER_WORD_11(6) => 
        \ELK_RX_SER_WORD_11[6]\, ELK_RX_SER_WORD_11(5) => 
        \ELK_RX_SER_WORD_11[5]\, ELK_RX_SER_WORD_11(4) => 
        \ELK_RX_SER_WORD_11[4]\, ELK_RX_SER_WORD_11(3) => 
        \ELK_RX_SER_WORD_11[3]\, ELK_RX_SER_WORD_11(2) => 
        \ELK_RX_SER_WORD_11[2]\, ELK_RX_SER_WORD_11(1) => 
        \ELK_RX_SER_WORD_11[1]\, ELK_RX_SER_WORD_11(0) => 
        \ELK_RX_SER_WORD_11[0]\, PATT_ELK_DAT_10(7) => 
        \PATT_ELK_DAT_10[7]\, PATT_ELK_DAT_10(6) => 
        \PATT_ELK_DAT_10[6]\, PATT_ELK_DAT_10(5) => 
        \PATT_ELK_DAT_10[5]\, PATT_ELK_DAT_10(4) => 
        \PATT_ELK_DAT_10[4]\, PATT_ELK_DAT_10(3) => 
        \PATT_ELK_DAT_10[3]\, PATT_ELK_DAT_10(2) => 
        \PATT_ELK_DAT_10[2]\, PATT_ELK_DAT_10(1) => 
        \PATT_ELK_DAT_10[1]\, PATT_ELK_DAT_10(0) => 
        \PATT_ELK_DAT_10[0]\, ELK_RX_SER_WORD_10(7) => 
        \ELK_RX_SER_WORD_10[7]\, ELK_RX_SER_WORD_10(6) => 
        \ELK_RX_SER_WORD_10[6]\, ELK_RX_SER_WORD_10(5) => 
        \ELK_RX_SER_WORD_10[5]\, ELK_RX_SER_WORD_10(4) => 
        \ELK_RX_SER_WORD_10[4]\, ELK_RX_SER_WORD_10(3) => 
        \ELK_RX_SER_WORD_10[3]\, ELK_RX_SER_WORD_10(2) => 
        \ELK_RX_SER_WORD_10[2]\, ELK_RX_SER_WORD_10(1) => 
        \ELK_RX_SER_WORD_10[1]\, ELK_RX_SER_WORD_10(0) => 
        \ELK_RX_SER_WORD_10[0]\, PATT_ELK_DAT_9(7) => 
        \PATT_ELK_DAT_9[7]\, PATT_ELK_DAT_9(6) => 
        \PATT_ELK_DAT_9[6]\, PATT_ELK_DAT_9(5) => 
        \PATT_ELK_DAT_9[5]\, PATT_ELK_DAT_9(4) => 
        \PATT_ELK_DAT_9[4]\, PATT_ELK_DAT_9(3) => 
        \PATT_ELK_DAT_9[3]\, PATT_ELK_DAT_9(2) => 
        \PATT_ELK_DAT_9[2]\, PATT_ELK_DAT_9(1) => 
        \PATT_ELK_DAT_9[1]\, PATT_ELK_DAT_9(0) => 
        \PATT_ELK_DAT_9[0]\, ELK_RX_SER_WORD_9(7) => 
        \ELK_RX_SER_WORD_9[7]\, ELK_RX_SER_WORD_9(6) => 
        \ELK_RX_SER_WORD_9[6]\, ELK_RX_SER_WORD_9(5) => 
        \ELK_RX_SER_WORD_9[5]\, ELK_RX_SER_WORD_9(4) => 
        \ELK_RX_SER_WORD_9[4]\, ELK_RX_SER_WORD_9(3) => 
        \ELK_RX_SER_WORD_9[3]\, ELK_RX_SER_WORD_9(2) => 
        \ELK_RX_SER_WORD_9[2]\, ELK_RX_SER_WORD_9(1) => 
        \ELK_RX_SER_WORD_9[1]\, ELK_RX_SER_WORD_9(0) => 
        \ELK_RX_SER_WORD_9[0]\, PATT_ELK_DAT_8(7) => 
        \PATT_ELK_DAT_8[7]\, PATT_ELK_DAT_8(6) => 
        \PATT_ELK_DAT_8[6]\, PATT_ELK_DAT_8(5) => 
        \PATT_ELK_DAT_8[5]\, PATT_ELK_DAT_8(4) => 
        \PATT_ELK_DAT_8[4]\, PATT_ELK_DAT_8(3) => 
        \PATT_ELK_DAT_8[3]\, PATT_ELK_DAT_8(2) => 
        \PATT_ELK_DAT_8[2]\, PATT_ELK_DAT_8(1) => 
        \PATT_ELK_DAT_8[1]\, PATT_ELK_DAT_8(0) => 
        \PATT_ELK_DAT_8[0]\, ELK_RX_SER_WORD_8(7) => 
        \ELK_RX_SER_WORD_8[7]\, ELK_RX_SER_WORD_8(6) => 
        \ELK_RX_SER_WORD_8[6]\, ELK_RX_SER_WORD_8(5) => 
        \ELK_RX_SER_WORD_8[5]\, ELK_RX_SER_WORD_8(4) => 
        \ELK_RX_SER_WORD_8[4]\, ELK_RX_SER_WORD_8(3) => 
        \ELK_RX_SER_WORD_8[3]\, ELK_RX_SER_WORD_8(2) => 
        \ELK_RX_SER_WORD_8[2]\, ELK_RX_SER_WORD_8(1) => 
        \ELK_RX_SER_WORD_8[1]\, ELK_RX_SER_WORD_8(0) => 
        \ELK_RX_SER_WORD_8[0]\, PATT_ELK_DAT_7(7) => 
        \PATT_ELK_DAT_7[7]\, PATT_ELK_DAT_7(6) => 
        \PATT_ELK_DAT_7[6]\, PATT_ELK_DAT_7(5) => 
        \PATT_ELK_DAT_7[5]\, PATT_ELK_DAT_7(4) => 
        \PATT_ELK_DAT_7[4]\, PATT_ELK_DAT_7(3) => 
        \PATT_ELK_DAT_7[3]\, PATT_ELK_DAT_7(2) => 
        \PATT_ELK_DAT_7[2]\, PATT_ELK_DAT_7(1) => 
        \PATT_ELK_DAT_7[1]\, PATT_ELK_DAT_7(0) => 
        \PATT_ELK_DAT_7[0]\, ELK_RX_SER_WORD_7(7) => 
        \ELK_RX_SER_WORD_7[7]\, ELK_RX_SER_WORD_7(6) => 
        \ELK_RX_SER_WORD_7[6]\, ELK_RX_SER_WORD_7(5) => 
        \ELK_RX_SER_WORD_7[5]\, ELK_RX_SER_WORD_7(4) => 
        \ELK_RX_SER_WORD_7[4]\, ELK_RX_SER_WORD_7(3) => 
        \ELK_RX_SER_WORD_7[3]\, ELK_RX_SER_WORD_7(2) => 
        \ELK_RX_SER_WORD_7[2]\, ELK_RX_SER_WORD_7(1) => 
        \ELK_RX_SER_WORD_7[1]\, ELK_RX_SER_WORD_7(0) => 
        \ELK_RX_SER_WORD_7[0]\, PATT_ELK_DAT_6(7) => 
        \PATT_ELK_DAT_6[7]\, PATT_ELK_DAT_6(6) => 
        \PATT_ELK_DAT_6[6]\, PATT_ELK_DAT_6(5) => 
        \PATT_ELK_DAT_6[5]\, PATT_ELK_DAT_6(4) => 
        \PATT_ELK_DAT_6[4]\, PATT_ELK_DAT_6(3) => 
        \PATT_ELK_DAT_6[3]\, PATT_ELK_DAT_6(2) => 
        \PATT_ELK_DAT_6[2]\, PATT_ELK_DAT_6(1) => 
        \PATT_ELK_DAT_6[1]\, PATT_ELK_DAT_6(0) => 
        \PATT_ELK_DAT_6[0]\, ELK_RX_SER_WORD_6(7) => 
        \ELK_RX_SER_WORD_6[7]\, ELK_RX_SER_WORD_6(6) => 
        \ELK_RX_SER_WORD_6[6]\, ELK_RX_SER_WORD_6(5) => 
        \ELK_RX_SER_WORD_6[5]\, ELK_RX_SER_WORD_6(4) => 
        \ELK_RX_SER_WORD_6[4]\, ELK_RX_SER_WORD_6(3) => 
        \ELK_RX_SER_WORD_6[3]\, ELK_RX_SER_WORD_6(2) => 
        \ELK_RX_SER_WORD_6[2]\, ELK_RX_SER_WORD_6(1) => 
        \ELK_RX_SER_WORD_6[1]\, ELK_RX_SER_WORD_6(0) => 
        \ELK_RX_SER_WORD_6[0]\, PATT_ELK_DAT_5(7) => 
        \PATT_ELK_DAT_5[7]\, PATT_ELK_DAT_5(6) => 
        \PATT_ELK_DAT_5[6]\, PATT_ELK_DAT_5(5) => 
        \PATT_ELK_DAT_5[5]\, PATT_ELK_DAT_5(4) => 
        \PATT_ELK_DAT_5[4]\, PATT_ELK_DAT_5(3) => 
        \PATT_ELK_DAT_5[3]\, PATT_ELK_DAT_5(2) => 
        \PATT_ELK_DAT_5[2]\, PATT_ELK_DAT_5(1) => 
        \PATT_ELK_DAT_5[1]\, PATT_ELK_DAT_5(0) => 
        \PATT_ELK_DAT_5[0]\, ELK_RX_SER_WORD_5(7) => 
        \ELK_RX_SER_WORD_5[7]\, ELK_RX_SER_WORD_5(6) => 
        \ELK_RX_SER_WORD_5[6]\, ELK_RX_SER_WORD_5(5) => 
        \ELK_RX_SER_WORD_5[5]\, ELK_RX_SER_WORD_5(4) => 
        \ELK_RX_SER_WORD_5[4]\, ELK_RX_SER_WORD_5(3) => 
        \ELK_RX_SER_WORD_5[3]\, ELK_RX_SER_WORD_5(2) => 
        \ELK_RX_SER_WORD_5[2]\, ELK_RX_SER_WORD_5(1) => 
        \ELK_RX_SER_WORD_5[1]\, ELK_RX_SER_WORD_5(0) => 
        \ELK_RX_SER_WORD_5[0]\, PATT_ELK_DAT_4(7) => 
        \PATT_ELK_DAT_4[7]\, PATT_ELK_DAT_4(6) => 
        \PATT_ELK_DAT_4[6]\, PATT_ELK_DAT_4(5) => 
        \PATT_ELK_DAT_4[5]\, PATT_ELK_DAT_4(4) => 
        \PATT_ELK_DAT_4[4]\, PATT_ELK_DAT_4(3) => 
        \PATT_ELK_DAT_4[3]\, PATT_ELK_DAT_4(2) => 
        \PATT_ELK_DAT_4[2]\, PATT_ELK_DAT_4(1) => 
        \PATT_ELK_DAT_4[1]\, PATT_ELK_DAT_4(0) => 
        \PATT_ELK_DAT_4[0]\, ELK_RX_SER_WORD_4(7) => 
        \ELK_RX_SER_WORD_4[7]\, ELK_RX_SER_WORD_4(6) => 
        \ELK_RX_SER_WORD_4[6]\, ELK_RX_SER_WORD_4(5) => 
        \ELK_RX_SER_WORD_4[5]\, ELK_RX_SER_WORD_4(4) => 
        \ELK_RX_SER_WORD_4[4]\, ELK_RX_SER_WORD_4(3) => 
        \ELK_RX_SER_WORD_4[3]\, ELK_RX_SER_WORD_4(2) => 
        \ELK_RX_SER_WORD_4[2]\, ELK_RX_SER_WORD_4(1) => 
        \ELK_RX_SER_WORD_4[1]\, ELK_RX_SER_WORD_4(0) => 
        \ELK_RX_SER_WORD_4[0]\, PATT_ELK_DAT_3(7) => 
        \PATT_ELK_DAT_3[7]\, PATT_ELK_DAT_3(6) => 
        \PATT_ELK_DAT_3[6]\, PATT_ELK_DAT_3(5) => 
        \PATT_ELK_DAT_3[5]\, PATT_ELK_DAT_3(4) => 
        \PATT_ELK_DAT_3[4]\, PATT_ELK_DAT_3(3) => 
        \PATT_ELK_DAT_3[3]\, PATT_ELK_DAT_3(2) => 
        \PATT_ELK_DAT_3[2]\, PATT_ELK_DAT_3(1) => 
        \PATT_ELK_DAT_3[1]\, PATT_ELK_DAT_3(0) => 
        \PATT_ELK_DAT_3[0]\, ELK_RX_SER_WORD_3(7) => 
        \ELK_RX_SER_WORD_3[7]\, ELK_RX_SER_WORD_3(6) => 
        \ELK_RX_SER_WORD_3[6]\, ELK_RX_SER_WORD_3(5) => 
        \ELK_RX_SER_WORD_3[5]\, ELK_RX_SER_WORD_3(4) => 
        \ELK_RX_SER_WORD_3[4]\, ELK_RX_SER_WORD_3(3) => 
        \ELK_RX_SER_WORD_3[3]\, ELK_RX_SER_WORD_3(2) => 
        \ELK_RX_SER_WORD_3[2]\, ELK_RX_SER_WORD_3(1) => 
        \ELK_RX_SER_WORD_3[1]\, ELK_RX_SER_WORD_3(0) => 
        \ELK_RX_SER_WORD_3[0]\, PATT_ELK_DAT_2(7) => 
        \PATT_ELK_DAT_2[7]\, PATT_ELK_DAT_2(6) => 
        \PATT_ELK_DAT_2[6]\, PATT_ELK_DAT_2(5) => 
        \PATT_ELK_DAT_2[5]\, PATT_ELK_DAT_2(4) => 
        \PATT_ELK_DAT_2[4]\, PATT_ELK_DAT_2(3) => 
        \PATT_ELK_DAT_2[3]\, PATT_ELK_DAT_2(2) => 
        \PATT_ELK_DAT_2[2]\, PATT_ELK_DAT_2(1) => 
        \PATT_ELK_DAT_2[1]\, PATT_ELK_DAT_2(0) => 
        \PATT_ELK_DAT_2[0]\, ELK_RX_SER_WORD_2(7) => 
        \ELK_RX_SER_WORD_2[7]\, ELK_RX_SER_WORD_2(6) => 
        \ELK_RX_SER_WORD_2[6]\, ELK_RX_SER_WORD_2(5) => 
        \ELK_RX_SER_WORD_2[5]\, ELK_RX_SER_WORD_2(4) => 
        \ELK_RX_SER_WORD_2[4]\, ELK_RX_SER_WORD_2(3) => 
        \ELK_RX_SER_WORD_2[3]\, ELK_RX_SER_WORD_2(2) => 
        \ELK_RX_SER_WORD_2[2]\, ELK_RX_SER_WORD_2(1) => 
        \ELK_RX_SER_WORD_2[1]\, ELK_RX_SER_WORD_2(0) => 
        \ELK_RX_SER_WORD_2[0]\, PATT_ELK_DAT_1(7) => 
        \PATT_ELK_DAT_1[7]\, PATT_ELK_DAT_1(6) => 
        \PATT_ELK_DAT_1[6]\, PATT_ELK_DAT_1(5) => 
        \PATT_ELK_DAT_1[5]\, PATT_ELK_DAT_1(4) => 
        \PATT_ELK_DAT_1[4]\, PATT_ELK_DAT_1(3) => 
        \PATT_ELK_DAT_1[3]\, PATT_ELK_DAT_1(2) => 
        \PATT_ELK_DAT_1[2]\, PATT_ELK_DAT_1(1) => 
        \PATT_ELK_DAT_1[1]\, PATT_ELK_DAT_1(0) => 
        \PATT_ELK_DAT_1[0]\, ELKS_ADDRB_0_0 => \ELKS_ADDRB_0[2]\, 
        ELKS_ADDRB_0_2 => \ELKS_ADDRB_0[4]\, ELKS_ADDRB_0_4 => 
        \ELKS_ADDRB_0[6]\, ELK_RX_SER_WORD_1(7) => 
        \ELK_RX_SER_WORD_1[7]\, ELK_RX_SER_WORD_1(6) => 
        \ELK_RX_SER_WORD_1[6]\, ELK_RX_SER_WORD_1(5) => 
        \ELK_RX_SER_WORD_1[5]\, ELK_RX_SER_WORD_1(4) => 
        \ELK_RX_SER_WORD_1[4]\, ELK_RX_SER_WORD_1(3) => 
        \ELK_RX_SER_WORD_1[3]\, ELK_RX_SER_WORD_1(2) => 
        \ELK_RX_SER_WORD_1[2]\, ELK_RX_SER_WORD_1(1) => 
        \ELK_RX_SER_WORD_1[1]\, ELK_RX_SER_WORD_1(0) => 
        \ELK_RX_SER_WORD_1[0]\, PATT_ELK_DAT_0(7) => 
        \PATT_ELK_DAT_0[7]\, PATT_ELK_DAT_0(6) => 
        \PATT_ELK_DAT_0[6]\, PATT_ELK_DAT_0(5) => 
        \PATT_ELK_DAT_0[5]\, PATT_ELK_DAT_0(4) => 
        \PATT_ELK_DAT_0[4]\, PATT_ELK_DAT_0(3) => 
        \PATT_ELK_DAT_0[3]\, PATT_ELK_DAT_0(2) => 
        \PATT_ELK_DAT_0[2]\, PATT_ELK_DAT_0(1) => 
        \PATT_ELK_DAT_0[1]\, PATT_ELK_DAT_0(0) => 
        \PATT_ELK_DAT_0[0]\, ELKS_ADDRB(7) => \ELKS_ADDRB[7]\, 
        ELKS_ADDRB(6) => \ELKS_ADDRB[6]\, ELKS_ADDRB(5) => 
        \ELKS_ADDRB[5]\, ELKS_ADDRB(4) => \ELKS_ADDRB[4]\, 
        ELKS_ADDRB(3) => \ELKS_ADDRB[3]\, ELKS_ADDRB(2) => 
        \ELKS_ADDRB[2]\, ELKS_ADDRB(1) => \ELKS_ADDRB[1]\, 
        ELKS_ADDRB(0) => \ELKS_ADDRB[0]\, ELK_RX_SER_WORD_0(7)
         => \ELK_RX_SER_WORD_0[7]\, ELK_RX_SER_WORD_0(6) => 
        \ELK_RX_SER_WORD_0[6]\, ELK_RX_SER_WORD_0(5) => 
        \ELK_RX_SER_WORD_0[5]\, ELK_RX_SER_WORD_0(4) => 
        \ELK_RX_SER_WORD_0[4]\, ELK_RX_SER_WORD_0(3) => 
        \ELK_RX_SER_WORD_0[3]\, ELK_RX_SER_WORD_0(2) => 
        \ELK_RX_SER_WORD_0[2]\, ELK_RX_SER_WORD_0(1) => 
        \ELK_RX_SER_WORD_0[1]\, ELK_RX_SER_WORD_0(0) => 
        \ELK_RX_SER_WORD_0[0]\, PATT_TFC_DAT(7) => 
        \PATT_TFC_DAT[7]\, PATT_TFC_DAT(6) => \PATT_TFC_DAT[6]\, 
        PATT_TFC_DAT(5) => \PATT_TFC_DAT[5]\, PATT_TFC_DAT(4) => 
        \PATT_TFC_DAT[4]\, PATT_TFC_DAT(3) => \PATT_TFC_DAT[3]\, 
        PATT_TFC_DAT(2) => \PATT_TFC_DAT[2]\, PATT_TFC_DAT(1) => 
        \PATT_TFC_DAT[1]\, PATT_TFC_DAT(0) => \PATT_TFC_DAT[0]\, 
        TFC_ADDRB(7) => \TFC_ADDRB[7]\, TFC_ADDRB(6) => 
        \TFC_ADDRB[6]\, TFC_ADDRB(5) => \TFC_ADDRB[5]\, 
        TFC_ADDRB(4) => \TFC_ADDRB[4]\, TFC_ADDRB(3) => 
        \TFC_ADDRB[3]\, TFC_ADDRB(2) => \TFC_ADDRB[2]\, 
        TFC_ADDRB(1) => \TFC_ADDRB[1]\, TFC_ADDRB(0) => 
        \TFC_ADDRB[0]\, TFC_RX_SER_WORD(7) => 
        \TFC_RX_SER_WORD[7]\, TFC_RX_SER_WORD(6) => 
        \TFC_RX_SER_WORD[6]\, TFC_RX_SER_WORD(5) => 
        \TFC_RX_SER_WORD[5]\, TFC_RX_SER_WORD(4) => 
        \TFC_RX_SER_WORD[4]\, TFC_RX_SER_WORD(3) => 
        \TFC_RX_SER_WORD[3]\, TFC_RX_SER_WORD(2) => 
        \TFC_RX_SER_WORD[2]\, TFC_RX_SER_WORD(1) => 
        \TFC_RX_SER_WORD[1]\, TFC_RX_SER_WORD(0) => 
        \TFC_RX_SER_WORD[0]\, P_MASTER_POR_B_c_0_0 => 
        P_MASTER_POR_B_c_0_0, P_MASTER_POR_B_c_1 => 
        P_MASTER_POR_B_c_1, P_MASTER_POR_B_c => P_MASTER_POR_B_c, 
        P_MASTER_POR_B_c_6 => P_MASTER_POR_B_c_6, 
        P_MASTER_POR_B_c_24 => P_MASTER_POR_B_c_24, 
        P_MASTER_POR_B_c_3 => P_MASTER_POR_B_c_3, 
        P_MASTER_POR_B_c_26 => P_MASTER_POR_B_c_26, 
        P_MASTER_POR_B_c_33 => P_MASTER_POR_B_c_33, 
        P_MASTER_POR_B_c_22_0 => P_MASTER_POR_B_c_22_0, 
        P_MASTER_POR_B_c_28 => P_MASTER_POR_B_c_28, 
        P_MASTER_POR_B_c_23 => P_MASTER_POR_B_c_23, 
        P_MASTER_POR_B_c_19 => P_MASTER_POR_B_c_19, 
        P_MASTER_POR_B_c_24_0 => P_MASTER_POR_B_c_24_0, 
        P_MASTER_POR_B_c_25 => P_MASTER_POR_B_c_25, 
        P_MASTER_POR_B_c_29 => P_MASTER_POR_B_c_29, 
        P_MASTER_POR_B_c_30 => P_MASTER_POR_B_c_30, 
        P_MASTER_POR_B_c_27 => P_MASTER_POR_B_c_27, 
        P_MASTER_POR_B_c_17 => P_MASTER_POR_B_c_17, 
        P_MASTER_POR_B_c_32 => P_MASTER_POR_B_c_32, 
        P_MASTER_POR_B_c_32_0 => P_MASTER_POR_B_c_32_0, 
        P_MASTER_POR_B_c_21 => P_MASTER_POR_B_c_21, 
        P_MASTER_POR_B_c_22 => P_MASTER_POR_B_c_22, 
        ELKS_RAM_BLKB_EN => ELKS_RAM_BLKB_EN, ELKS_RWB => 
        ELKS_RWB, TFC_RAM_BLKB_EN => TFC_RAM_BLKB_EN, CLK_40M_GL
         => CLK_40M_GL, TFC_RWB => TFC_RWB, P_USB_MASTER_EN_c_1
         => P_USB_MASTER_EN_c_1, P_USB_MASTER_EN_c_0 => 
        P_USB_MASTER_EN_c_0, P_USB_MASTER_EN_c_2 => 
        P_USB_MASTER_EN_c_2, P_USB_MASTER_EN_c_20 => 
        P_USB_MASTER_EN_c_20, P_USB_MASTER_EN_c_6 => 
        P_USB_MASTER_EN_c_6, P_USB_MASTER_EN_c_9 => 
        P_USB_MASTER_EN_c_9, P_USB_MASTER_EN_c_11 => 
        P_USB_MASTER_EN_c_11, P_USB_MASTER_EN_c_12 => 
        P_USB_MASTER_EN_c_12, P_USB_MASTER_EN_c_14 => 
        P_USB_MASTER_EN_c_14, P_USB_MASTER_EN_c_18 => 
        P_USB_MASTER_EN_c_18, P_USB_MASTER_EN_c_7 => 
        P_USB_MASTER_EN_c_7, P_USB_MASTER_EN_c_21 => 
        P_USB_MASTER_EN_c_21, P_USB_MASTER_EN_c_17 => 
        P_USB_MASTER_EN_c_17, P_USB_MASTER_EN_c_15 => 
        P_USB_MASTER_EN_c_15, P_USB_MASTER_EN_c_4 => 
        P_USB_MASTER_EN_c_4, USB_WR_BI => USB_WR_BI, 
        P_USB_MASTER_EN_c_3 => P_USB_MASTER_EN_c_3, 
        P_USB_MASTER_EN_c_8 => P_USB_MASTER_EN_c_8, USB_SIWU_BI
         => USB_SIWU_BI, P_USB_MASTER_EN_c_19 => 
        P_USB_MASTER_EN_c_19, USB_OE_BI => USB_OE_BI, USB_RD_BI
         => USB_RD_BI, P_USB_MASTER_EN_c_13 => 
        P_USB_MASTER_EN_c_13, P_USB_MASTER_EN_c_5 => 
        P_USB_MASTER_EN_c_5, P_USB_MASTER_EN_c_10 => 
        P_USB_MASTER_EN_c_10, P_USB_MASTER_EN_c_22 => 
        P_USB_MASTER_EN_c_22, P_USB_TXE_B_c => P_USB_TXE_B_c, 
        P_USB_MASTER_EN_c_16 => P_USB_MASTER_EN_c_16, 
        P_USB_MASTER_EN_c_22_0 => P_USB_MASTER_EN_c_22_0, 
        P_USB_MASTER_EN_c_2_0 => P_USB_MASTER_EN_c_2_0, 
        P_USB_MASTER_EN_c_1_0 => P_USB_MASTER_EN_c_1_0, 
        P_USB_MASTER_EN_c => P_USB_MASTER_EN_c, P_USB_RXF_B_c => 
        P_USB_RXF_B_c, CLK60MHZ => CLK60MHZ);
    
    P_OP_MODE6_EE_pad : OUTBUF
      port map(D => \OP_MODE_c[6]\, PAD => P_OP_MODE6_EE);
    
    P_USB_TXE_B_pad : INBUF
      port map(PAD => P_USB_TXE_B, Y => P_USB_TXE_B_c);
    
    ELK0_IN_F : DFN1C0
      port map(D => ELK0_IN_DDR_F_i, CLK => CCC_160M_ADJ, CLR => 
        DEV_RST_B_c, Q => \ELK0_IN_F\);
    
    U_TFC_SERDAT_SOURCE : SYNC_DAT_SEL
      port map(TFC_TX_DAT(7) => \TFC_TX_DAT[7]\, TFC_TX_DAT(6)
         => \TFC_TX_DAT[6]\, TFC_TX_DAT(5) => \TFC_TX_DAT[5]\, 
        TFC_TX_DAT(4) => \TFC_TX_DAT[4]\, TFC_TX_DAT(3) => 
        \TFC_TX_DAT[3]\, TFC_TX_DAT(2) => \TFC_TX_DAT[2]\, 
        TFC_TX_DAT(1) => \TFC_TX_DAT[1]\, TFC_TX_DAT(0) => 
        \TFC_TX_DAT[0]\, PATT_TFC_DAT(7) => \PATT_TFC_DAT[7]\, 
        PATT_TFC_DAT(6) => \PATT_TFC_DAT[6]\, PATT_TFC_DAT(5) => 
        \PATT_TFC_DAT[5]\, PATT_TFC_DAT(4) => \PATT_TFC_DAT[4]\, 
        PATT_TFC_DAT(3) => \PATT_TFC_DAT[3]\, PATT_TFC_DAT(2) => 
        \PATT_TFC_DAT[2]\, PATT_TFC_DAT(1) => \PATT_TFC_DAT[1]\, 
        PATT_TFC_DAT(0) => \PATT_TFC_DAT[0]\, OP_MODE_c_0_0 => 
        \OP_MODE_c_0[1]\, MASTER_DCB_POR_B_i_0_i => 
        MASTER_DCB_POR_B_i_0_i, CLK_40M_GL => CLK_40M_GL);
    
    U_MAINCLKGEN : CLK_FXD_40_160_A60M
      port map(USBCLK60MHZ_c => USBCLK60MHZ_c, CCC_MAIN_LOCK => 
        CCC_MAIN_LOCK, CLK60MHZ_1 => CLK60MHZ, CCC_160M_FXD_1 => 
        CCC_160M_FXD, CLK_40M_GL_1 => CLK_40M_GL, 
        CLK_40M_BUF_RECD => CLK_40M_BUF_RECD);
    
    U_ELK18_CH : ELINK_SLAVE_15_13
      port map(BIT_OS_SEL_0(2) => \BIT_OS_SEL_0[2]\, 
        BIT_OS_SEL_0(1) => \BIT_OS_SEL_0[1]\, BIT_OS_SEL_1(2) => 
        \BIT_OS_SEL_1[2]\, BIT_OS_SEL_1(1) => \BIT_OS_SEL_1[1]\, 
        BIT_OS_SEL_2(1) => \BIT_OS_SEL_2[1]\, BIT_OS_SEL_2(0) => 
        \BIT_OS_SEL_2[0]\, ELK_RX_SER_WORD_18(7) => 
        \ELK_RX_SER_WORD_18[7]\, ELK_RX_SER_WORD_18(6) => 
        \ELK_RX_SER_WORD_18[6]\, ELK_RX_SER_WORD_18(5) => 
        \ELK_RX_SER_WORD_18[5]\, ELK_RX_SER_WORD_18(4) => 
        \ELK_RX_SER_WORD_18[4]\, ELK_RX_SER_WORD_18(3) => 
        \ELK_RX_SER_WORD_18[3]\, ELK_RX_SER_WORD_18(2) => 
        \ELK_RX_SER_WORD_18[2]\, ELK_RX_SER_WORD_18(1) => 
        \ELK_RX_SER_WORD_18[1]\, ELK_RX_SER_WORD_18(0) => 
        \ELK_RX_SER_WORD_18[0]\, OP_MODE_c_1_0 => 
        \OP_MODE_c_1[1]\, OP_MODE_c_2_0 => \OP_MODE_c_2[1]\, 
        PATT_ELK_DAT_18(7) => \PATT_ELK_DAT_18[7]\, 
        PATT_ELK_DAT_18(6) => \PATT_ELK_DAT_18[6]\, 
        PATT_ELK_DAT_18(5) => \PATT_ELK_DAT_18[5]\, 
        PATT_ELK_DAT_18(4) => \PATT_ELK_DAT_18[4]\, 
        PATT_ELK_DAT_18(3) => \PATT_ELK_DAT_18[3]\, 
        PATT_ELK_DAT_18(2) => \PATT_ELK_DAT_18[2]\, 
        PATT_ELK_DAT_18(1) => \PATT_ELK_DAT_18[1]\, 
        PATT_ELK_DAT_18(0) => \PATT_ELK_DAT_18[0]\, 
        MASTER_DCB_POR_B_i_0_i => MASTER_DCB_POR_B_i_0_i, 
        ELK18_DAT_N => ELK18_DAT_N, ELK18_DAT_P => ELK18_DAT_P, 
        DCB_SALT_SEL_c_i => DCB_SALT_SEL_c_i, CCC_160M_FXD => 
        CCC_160M_FXD, MASTER_SALT_POR_B_i_0_i_9 => 
        MASTER_SALT_POR_B_i_0_i_9, MASTER_SALT_POR_B_i_0_i_4 => 
        MASTER_SALT_POR_B_i_0_i_4, MASTER_SALT_POR_B_i_0_i_1 => 
        MASTER_SALT_POR_B_i_0_i_1, MASTER_SALT_POR_B_i_0_i_17 => 
        MASTER_SALT_POR_B_i_0_i_17, MASTER_SALT_POR_B_i_0_i_3 => 
        MASTER_SALT_POR_B_i_0_i_3, MASTER_SALT_POR_B_i_0_i_0 => 
        MASTER_SALT_POR_B_i_0_i_0, CLK_40M_GL => CLK_40M_GL, 
        MASTER_SALT_POR_B_i_0_i_13 => MASTER_SALT_POR_B_i_0_i_13, 
        DEV_RST_B_c_0 => DEV_RST_B_c_0, CCC_160M_ADJ => 
        CCC_160M_ADJ);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    U62_TS_OE_BUF : tristate_buf_1
      port map(P_USB_MASTER_EN_c => P_USB_MASTER_EN_c, USB_OE_BI
         => USB_OE_BI, USB_OE_B => USB_OE_B);
    
    TFC_IN_R : DFN1C0
      port map(D => TFC_IN_DDR_R, CLK => CCC_160M_ADJ, CLR => 
        DEV_RST_B_c_0, Q => \TFC_IN_R\);
    
    P_MASTER_POR_B_pad : OUTBUF
      port map(D => P_MASTER_POR_B_c, PAD => P_MASTER_POR_B);
    
    U_REFCLKBUF : BIDIR_LVDS_IO_0
      port map(DCB_SALT_SEL_c => DCB_SALT_SEL_c, CLK_40M_GL => 
        CLK_40M_GL, EXTCLK_40MHZ_c => EXTCLK_40MHZ_c, REF_CLK_0P
         => REF_CLK_0P, REF_CLK_0N => REF_CLK_0N);
    
    U_ELK11_CH : ELINK_SLAVE_15_6
      port map(BIT_OS_SEL_4(2) => \BIT_OS_SEL_4[2]\, 
        BIT_OS_SEL_4(1) => \BIT_OS_SEL_4[1]\, BIT_OS_SEL_5(2) => 
        \BIT_OS_SEL_5[2]\, BIT_OS_SEL_5(1) => \BIT_OS_SEL_5[1]\, 
        BIT_OS_SEL_7_0 => \BIT_OS_SEL_7[2]\, BIT_OS_SEL_6_0 => 
        \BIT_OS_SEL_6[1]\, BIT_OS_SEL_0 => \BIT_OS_SEL[0]\, 
        ELK_RX_SER_WORD_11(7) => \ELK_RX_SER_WORD_11[7]\, 
        ELK_RX_SER_WORD_11(6) => \ELK_RX_SER_WORD_11[6]\, 
        ELK_RX_SER_WORD_11(5) => \ELK_RX_SER_WORD_11[5]\, 
        ELK_RX_SER_WORD_11(4) => \ELK_RX_SER_WORD_11[4]\, 
        ELK_RX_SER_WORD_11(3) => \ELK_RX_SER_WORD_11[3]\, 
        ELK_RX_SER_WORD_11(2) => \ELK_RX_SER_WORD_11[2]\, 
        ELK_RX_SER_WORD_11(1) => \ELK_RX_SER_WORD_11[1]\, 
        ELK_RX_SER_WORD_11(0) => \ELK_RX_SER_WORD_11[0]\, 
        OP_MODE_c_0 => \OP_MODE_c[1]\, PATT_ELK_DAT_11(7) => 
        \PATT_ELK_DAT_11[7]\, PATT_ELK_DAT_11(6) => 
        \PATT_ELK_DAT_11[6]\, PATT_ELK_DAT_11(5) => 
        \PATT_ELK_DAT_11[5]\, PATT_ELK_DAT_11(4) => 
        \PATT_ELK_DAT_11[4]\, PATT_ELK_DAT_11(3) => 
        \PATT_ELK_DAT_11[3]\, PATT_ELK_DAT_11(2) => 
        \PATT_ELK_DAT_11[2]\, PATT_ELK_DAT_11(1) => 
        \PATT_ELK_DAT_11[1]\, PATT_ELK_DAT_11(0) => 
        \PATT_ELK_DAT_11[0]\, MASTER_DCB_POR_B_i_0_i => 
        MASTER_DCB_POR_B_i_0_i, ELK11_DAT_N => ELK11_DAT_N, 
        ELK11_DAT_P => ELK11_DAT_P, DCB_SALT_SEL_c_i => 
        DCB_SALT_SEL_c_i, CCC_160M_FXD => CCC_160M_FXD, 
        MASTER_SALT_POR_B_i_0_i_5 => MASTER_SALT_POR_B_i_0_i_5, 
        MASTER_SALT_POR_B_i_0_i_16 => MASTER_SALT_POR_B_i_0_i_16, 
        MASTER_SALT_POR_B_i_0_i_10 => MASTER_SALT_POR_B_i_0_i_10, 
        MASTER_SALT_POR_B_i_0_i_2 => MASTER_SALT_POR_B_i_0_i_2, 
        MASTER_SALT_POR_B_i_0_i_11 => MASTER_SALT_POR_B_i_0_i_11, 
        MASTER_SALT_POR_B_i_0_i_7 => MASTER_SALT_POR_B_i_0_i_7, 
        CLK_40M_GL => CLK_40M_GL, MASTER_SALT_POR_B_i_0_i_0 => 
        MASTER_SALT_POR_B_i_0_i_0, DEV_RST_B_c_0 => DEV_RST_B_c_0, 
        CCC_160M_ADJ => CCC_160M_ADJ);
    
    U200B_ELINKS : GP_PATT_GEN_1_0
      port map(ELKS_ADDRB(7) => \ELKS_ADDRB[7]\, ELKS_ADDRB(6)
         => \ELKS_ADDRB[6]\, ELKS_ADDRB(5) => \ELKS_ADDRB[5]\, 
        ELKS_ADDRB(4) => \ELKS_ADDRB[4]\, ELKS_ADDRB(3) => 
        \ELKS_ADDRB[3]\, ELKS_ADDRB(2) => \ELKS_ADDRB[2]\, 
        ELKS_ADDRB(1) => \ELKS_ADDRB[1]\, ELKS_ADDRB(0) => 
        \ELKS_ADDRB[0]\, ELK_RX_SER_WORD_0(7) => 
        \ELK_RX_SER_WORD_0[7]\, ELK_RX_SER_WORD_0(6) => 
        \ELK_RX_SER_WORD_0[6]\, ELK_RX_SER_WORD_0(5) => 
        \ELK_RX_SER_WORD_0[5]\, ELK_RX_SER_WORD_0(4) => 
        \ELK_RX_SER_WORD_0[4]\, ELK_RX_SER_WORD_0(3) => 
        \ELK_RX_SER_WORD_0[3]\, ELK_RX_SER_WORD_0(2) => 
        \ELK_RX_SER_WORD_0[2]\, ELK_RX_SER_WORD_0(1) => 
        \ELK_RX_SER_WORD_0[1]\, ELK_RX_SER_WORD_0(0) => 
        \ELK_RX_SER_WORD_0[0]\, ELKS_STOP_ADDR(7) => 
        \ELKS_STOP_ADDR[7]\, ELKS_STOP_ADDR(6) => 
        \ELKS_STOP_ADDR[6]\, ELKS_STOP_ADDR(5) => 
        \ELKS_STOP_ADDR[5]\, ELKS_STOP_ADDR(4) => 
        \ELKS_STOP_ADDR[4]\, ELKS_STOP_ADDR(3) => 
        \ELKS_STOP_ADDR[3]\, ELKS_STOP_ADDR(2) => 
        \ELKS_STOP_ADDR[2]\, ELKS_STOP_ADDR(1) => 
        \ELKS_STOP_ADDR[1]\, ELKS_STOP_ADDR(0) => 
        \ELKS_STOP_ADDR[0]\, ELKS_STRT_ADDR(7) => 
        \ELKS_STRT_ADDR[7]\, ELKS_STRT_ADDR(6) => 
        \ELKS_STRT_ADDR[6]\, ELKS_STRT_ADDR(5) => 
        \ELKS_STRT_ADDR[5]\, ELKS_STRT_ADDR(4) => 
        \ELKS_STRT_ADDR[4]\, ELKS_STRT_ADDR(3) => 
        \ELKS_STRT_ADDR[3]\, ELKS_STRT_ADDR(2) => 
        \ELKS_STRT_ADDR[2]\, ELKS_STRT_ADDR(1) => 
        \ELKS_STRT_ADDR[1]\, ELKS_STRT_ADDR(0) => 
        \ELKS_STRT_ADDR[0]\, OP_MODE_0 => \OP_MODE[4]\, 
        OP_MODE_c_0 => \OP_MODE_c[6]\, ELKS_ADDRB_0_0 => 
        \ELKS_ADDRB_0[2]\, ELKS_ADDRB_0_2 => \ELKS_ADDRB_0[4]\, 
        ELKS_ADDRB_0_4 => \ELKS_ADDRB_0[6]\, P_MASTER_POR_B_c_32
         => P_MASTER_POR_B_c_32, P_MASTER_POR_B_c_26 => 
        P_MASTER_POR_B_c_26, P_MASTER_POR_B_c_25 => 
        P_MASTER_POR_B_c_25, P_MASTER_POR_B_c_23 => 
        P_MASTER_POR_B_c_23, P_MASTER_POR_B_c_7 => 
        P_MASTER_POR_B_c_7, P_MASTER_POR_B_c_11 => 
        P_MASTER_POR_B_c_11, P_MASTER_POR_B_c_29 => 
        P_MASTER_POR_B_c_29, DCB_SALT_SEL_c_i => DCB_SALT_SEL_c_i, 
        P_MASTER_POR_B_c_2 => P_MASTER_POR_B_c_2, 
        P_MASTER_POR_B_c_12 => P_MASTER_POR_B_c_12, ELKS_RWB => 
        ELKS_RWB, P_MASTER_POR_B_c_13 => P_MASTER_POR_B_c_13, 
        ELKS_RAM_BLKB_EN => ELKS_RAM_BLKB_EN, P_USB_MASTER_EN_c
         => P_USB_MASTER_EN_c, ALIGN_ACTIVE => ALIGN_ACTIVE, 
        P_MASTER_POR_B_c_34_0 => P_MASTER_POR_B_c_34_0, 
        P_MASTER_POR_B_c_32_0 => P_MASTER_POR_B_c_32_0, 
        P_MASTER_POR_B_c_31_0 => P_MASTER_POR_B_c_31_0, 
        CLK_40M_GL => CLK_40M_GL);
    
    DEV_RST_B_pad_RNICBV3 : BUFF
      port map(A => DEV_RST_B_c, Y => DEV_RST_B_c_0);
    
    ALL_PLL_LOCK_pad : OUTBUF
      port map(D => ALL_PLL_LOCK_c, PAD => ALL_PLL_LOCK);
    
    P_CCC_160M_FXD_pad : OUTBUF
      port map(D => CCC_160M_FXD, PAD => P_CCC_160M_FXD);
    
    DEV_RST_B_pad_RNICBV3_0 : BUFF
      port map(A => DEV_RST_B_c, Y => DEV_RST_B_c_1);
    
    U_TFC_CMD_TX : SER320M_3_34
      port map(TFC_TX_DAT(7) => \TFC_TX_DAT[7]\, TFC_TX_DAT(6)
         => \TFC_TX_DAT[6]\, TFC_TX_DAT(5) => \TFC_TX_DAT[5]\, 
        TFC_TX_DAT(4) => \TFC_TX_DAT[4]\, TFC_TX_DAT(3) => 
        \TFC_TX_DAT[3]\, TFC_TX_DAT(2) => \TFC_TX_DAT[2]\, 
        TFC_TX_DAT(1) => \TFC_TX_DAT[1]\, TFC_TX_DAT(0) => 
        \TFC_TX_DAT[0]\, TFC_OUT_R => TFC_OUT_R, TFC_OUT_F => 
        TFC_OUT_F, MASTER_DCB_POR_B_i_0_i => 
        MASTER_DCB_POR_B_i_0_i, CCC_160M_FXD => CCC_160M_FXD, 
        CLK_40M_GL => CLK_40M_GL);
    
    U_ELK0_CMD_TX : SER320M_3_34_0
      port map(ELK0_TX_DAT(7) => \ELK0_TX_DAT[7]\, ELK0_TX_DAT(6)
         => \ELK0_TX_DAT[6]\, ELK0_TX_DAT(5) => \ELK0_TX_DAT[5]\, 
        ELK0_TX_DAT(4) => \ELK0_TX_DAT[4]\, ELK0_TX_DAT(3) => 
        \ELK0_TX_DAT[3]\, ELK0_TX_DAT(2) => \ELK0_TX_DAT[2]\, 
        ELK0_TX_DAT(1) => \ELK0_TX_DAT[1]\, ELK0_TX_DAT(0) => 
        \ELK0_TX_DAT[0]\, MASTER_SALT_POR_B_i_0_i_17 => 
        MASTER_SALT_POR_B_i_0_i_17, MASTER_SALT_POR_B_i_0_i_3 => 
        MASTER_SALT_POR_B_i_0_i_3, MASTER_SALT_POR_B_i_0_i_7 => 
        MASTER_SALT_POR_B_i_0_i_7, ELK0_OUT_R_i_0 => 
        ELK0_OUT_R_i_0, MASTER_SALT_POR_B_i_0_i_10 => 
        MASTER_SALT_POR_B_i_0_i_10, ELK0_OUT_F_i_0 => 
        ELK0_OUT_F_i_0, MASTER_SALT_POR_B_i_0_i_5 => 
        MASTER_SALT_POR_B_i_0_i_5, CLK_40M_GL => CLK_40M_GL, 
        MASTER_SALT_POR_B_i_0_i_13 => MASTER_SALT_POR_B_i_0_i_13, 
        MASTER_SALT_POR_B_i_0_i_14 => MASTER_SALT_POR_B_i_0_i_14, 
        CCC_160M_FXD => CCC_160M_FXD);
    
    EXT_INT_REF_SEL_pad : INBUF
      port map(PAD => EXT_INT_REF_SEL, Y => EXT_INT_REF_SEL_c);
    
    U_ELK12_CH : ELINK_SLAVE_15_7
      port map(BIT_OS_SEL_3_0 => \BIT_OS_SEL_3[2]\, 
        BIT_OS_SEL_4(2) => \BIT_OS_SEL_4[2]\, BIT_OS_SEL_4(1) => 
        \BIT_OS_SEL_4[1]\, BIT_OS_SEL_6(2) => \BIT_OS_SEL_6[2]\, 
        BIT_OS_SEL_6(1) => \BIT_OS_SEL_6[1]\, BIT_OS_SEL_5_0 => 
        \BIT_OS_SEL_5[0]\, ELK_RX_SER_WORD_12(7) => 
        \ELK_RX_SER_WORD_12[7]\, ELK_RX_SER_WORD_12(6) => 
        \ELK_RX_SER_WORD_12[6]\, ELK_RX_SER_WORD_12(5) => 
        \ELK_RX_SER_WORD_12[5]\, ELK_RX_SER_WORD_12(4) => 
        \ELK_RX_SER_WORD_12[4]\, ELK_RX_SER_WORD_12(3) => 
        \ELK_RX_SER_WORD_12[3]\, ELK_RX_SER_WORD_12(2) => 
        \ELK_RX_SER_WORD_12[2]\, ELK_RX_SER_WORD_12(1) => 
        \ELK_RX_SER_WORD_12[1]\, ELK_RX_SER_WORD_12(0) => 
        \ELK_RX_SER_WORD_12[0]\, OP_MODE_c_2_0 => 
        \OP_MODE_c_2[1]\, OP_MODE_c_3_0 => \OP_MODE_c_3[1]\, 
        PATT_ELK_DAT_12(7) => \PATT_ELK_DAT_12[7]\, 
        PATT_ELK_DAT_12(6) => \PATT_ELK_DAT_12[6]\, 
        PATT_ELK_DAT_12(5) => \PATT_ELK_DAT_12[5]\, 
        PATT_ELK_DAT_12(4) => \PATT_ELK_DAT_12[4]\, 
        PATT_ELK_DAT_12(3) => \PATT_ELK_DAT_12[3]\, 
        PATT_ELK_DAT_12(2) => \PATT_ELK_DAT_12[2]\, 
        PATT_ELK_DAT_12(1) => \PATT_ELK_DAT_12[1]\, 
        PATT_ELK_DAT_12(0) => \PATT_ELK_DAT_12[0]\, 
        MASTER_DCB_POR_B_i_0_i => MASTER_DCB_POR_B_i_0_i, 
        ELK12_DAT_N => ELK12_DAT_N, ELK12_DAT_P => ELK12_DAT_P, 
        DCB_SALT_SEL_c_i => DCB_SALT_SEL_c_i, CCC_160M_FXD => 
        CCC_160M_FXD, MASTER_SALT_POR_B_i_0_i_6 => 
        MASTER_SALT_POR_B_i_0_i_6, MASTER_SALT_POR_B_i_0_i_12 => 
        MASTER_SALT_POR_B_i_0_i_12, MASTER_SALT_POR_B_i_0_i_8 => 
        MASTER_SALT_POR_B_i_0_i_8, MASTER_SALT_POR_B_i_0_i_0 => 
        MASTER_SALT_POR_B_i_0_i_0, MASTER_SALT_POR_B_i_0_i_10 => 
        MASTER_SALT_POR_B_i_0_i_10, MASTER_SALT_POR_B_i_0_i_15
         => MASTER_SALT_POR_B_i_0_i_15, CLK_40M_GL => CLK_40M_GL, 
        MASTER_SALT_POR_B_i_0_i_2 => MASTER_SALT_POR_B_i_0_i_2, 
        DEV_RST_B_c => DEV_RST_B_c, CCC_160M_ADJ => CCC_160M_ADJ);
    
    U_ELK13_CH : ELINK_SLAVE_15_8
      port map(BIT_OS_SEL_2_0 => \BIT_OS_SEL_2[2]\, 
        BIT_OS_SEL_3(2) => \BIT_OS_SEL_3[2]\, BIT_OS_SEL_3(1) => 
        \BIT_OS_SEL_3[1]\, BIT_OS_SEL_6_0 => \BIT_OS_SEL_6[2]\, 
        BIT_OS_SEL_5_0 => \BIT_OS_SEL_5[1]\, BIT_OS_SEL_4_0 => 
        \BIT_OS_SEL_4[0]\, ELK_RX_SER_WORD_13(7) => 
        \ELK_RX_SER_WORD_13[7]\, ELK_RX_SER_WORD_13(6) => 
        \ELK_RX_SER_WORD_13[6]\, ELK_RX_SER_WORD_13(5) => 
        \ELK_RX_SER_WORD_13[5]\, ELK_RX_SER_WORD_13(4) => 
        \ELK_RX_SER_WORD_13[4]\, ELK_RX_SER_WORD_13(3) => 
        \ELK_RX_SER_WORD_13[3]\, ELK_RX_SER_WORD_13(2) => 
        \ELK_RX_SER_WORD_13[2]\, ELK_RX_SER_WORD_13(1) => 
        \ELK_RX_SER_WORD_13[1]\, ELK_RX_SER_WORD_13(0) => 
        \ELK_RX_SER_WORD_13[0]\, OP_MODE_c_6_0 => 
        \OP_MODE_c_6[1]\, OP_MODE_c_0 => \OP_MODE_c[1]\, 
        PATT_ELK_DAT_13(7) => \PATT_ELK_DAT_13[7]\, 
        PATT_ELK_DAT_13(6) => \PATT_ELK_DAT_13[6]\, 
        PATT_ELK_DAT_13(5) => \PATT_ELK_DAT_13[5]\, 
        PATT_ELK_DAT_13(4) => \PATT_ELK_DAT_13[4]\, 
        PATT_ELK_DAT_13(3) => \PATT_ELK_DAT_13[3]\, 
        PATT_ELK_DAT_13(2) => \PATT_ELK_DAT_13[2]\, 
        PATT_ELK_DAT_13(1) => \PATT_ELK_DAT_13[1]\, 
        PATT_ELK_DAT_13(0) => \PATT_ELK_DAT_13[0]\, 
        MASTER_DCB_POR_B_i_0_i => MASTER_DCB_POR_B_i_0_i, 
        ELK13_DAT_N => ELK13_DAT_N, ELK13_DAT_P => ELK13_DAT_P, 
        DCB_SALT_SEL_c_i => DCB_SALT_SEL_c_i, CCC_160M_FXD => 
        CCC_160M_FXD, MASTER_SALT_POR_B_i_0_i_6 => 
        MASTER_SALT_POR_B_i_0_i_6, MASTER_SALT_POR_B_i_0_i_1 => 
        MASTER_SALT_POR_B_i_0_i_1, MASTER_SALT_POR_B_i_0_i_9 => 
        MASTER_SALT_POR_B_i_0_i_9, MASTER_SALT_POR_B_i_0_i_16 => 
        MASTER_SALT_POR_B_i_0_i_16, CLK_40M_GL => CLK_40M_GL, 
        MASTER_SALT_POR_B_i_0_i_4 => MASTER_SALT_POR_B_i_0_i_4, 
        DEV_RST_B_c => DEV_RST_B_c, CCC_160M_ADJ => CCC_160M_ADJ);
    
    U_ELK0_SERDAT_SOURCE : SYNC_DAT_SEL_0
      port map(ELK0_TX_DAT(7) => \ELK0_TX_DAT[7]\, ELK0_TX_DAT(6)
         => \ELK0_TX_DAT[6]\, ELK0_TX_DAT(5) => \ELK0_TX_DAT[5]\, 
        ELK0_TX_DAT(4) => \ELK0_TX_DAT[4]\, ELK0_TX_DAT(3) => 
        \ELK0_TX_DAT[3]\, ELK0_TX_DAT(2) => \ELK0_TX_DAT[2]\, 
        ELK0_TX_DAT(1) => \ELK0_TX_DAT[1]\, ELK0_TX_DAT(0) => 
        \ELK0_TX_DAT[0]\, PATT_ELK_DAT_0(7) => 
        \PATT_ELK_DAT_0[7]\, PATT_ELK_DAT_0(6) => 
        \PATT_ELK_DAT_0[6]\, PATT_ELK_DAT_0(5) => 
        \PATT_ELK_DAT_0[5]\, PATT_ELK_DAT_0(4) => 
        \PATT_ELK_DAT_0[4]\, PATT_ELK_DAT_0(3) => 
        \PATT_ELK_DAT_0[3]\, PATT_ELK_DAT_0(2) => 
        \PATT_ELK_DAT_0[2]\, PATT_ELK_DAT_0(1) => 
        \PATT_ELK_DAT_0[1]\, PATT_ELK_DAT_0(0) => 
        \PATT_ELK_DAT_0[0]\, OP_MODE_c_4_0 => \OP_MODE_c_4[1]\, 
        MASTER_SALT_POR_B_i_0_i_10 => MASTER_SALT_POR_B_i_0_i_10, 
        CLK_40M_GL => CLK_40M_GL);
    
    GND_i : GND
      port map(Y => \GND\);
    
    U_EXEC_MASTER : EXEC_MODE_CNTL
      port map(CLK60MHZ => CLK60MHZ, P_USB_MASTER_EN_c_1_0 => 
        P_USB_MASTER_EN_c_1_0, P_USB_MASTER_EN_c_2_0 => 
        P_USB_MASTER_EN_c_2_0, P_USB_MASTER_EN_c_22_0 => 
        P_USB_MASTER_EN_c_22_0, P_USB_MASTER_EN_c_22 => 
        P_USB_MASTER_EN_c_22, P_USB_MASTER_EN_c_21 => 
        P_USB_MASTER_EN_c_21, P_USB_MASTER_EN_c_20 => 
        P_USB_MASTER_EN_c_20, P_USB_MASTER_EN_c_19 => 
        P_USB_MASTER_EN_c_19, P_USB_MASTER_EN_c_18 => 
        P_USB_MASTER_EN_c_18, P_USB_MASTER_EN_c_17 => 
        P_USB_MASTER_EN_c_17, P_USB_MASTER_EN_c_16 => 
        P_USB_MASTER_EN_c_16, P_USB_MASTER_EN_c_15 => 
        P_USB_MASTER_EN_c_15, P_USB_MASTER_EN_c_14 => 
        P_USB_MASTER_EN_c_14, P_USB_MASTER_EN_c_13 => 
        P_USB_MASTER_EN_c_13, P_USB_MASTER_EN_c_12 => 
        P_USB_MASTER_EN_c_12, P_USB_MASTER_EN_c_11 => 
        P_USB_MASTER_EN_c_11, P_USB_MASTER_EN_c_10 => 
        P_USB_MASTER_EN_c_10, P_USB_MASTER_EN_c_9 => 
        P_USB_MASTER_EN_c_9, P_USB_MASTER_EN_c_8 => 
        P_USB_MASTER_EN_c_8, P_USB_MASTER_EN_c_7 => 
        P_USB_MASTER_EN_c_7, P_USB_MASTER_EN_c_6 => 
        P_USB_MASTER_EN_c_6, P_USB_MASTER_EN_c_5 => 
        P_USB_MASTER_EN_c_5, P_USB_MASTER_EN_c_4 => 
        P_USB_MASTER_EN_c_4, P_USB_MASTER_EN_c_3 => 
        P_USB_MASTER_EN_c_3, P_USB_MASTER_EN_c_2 => 
        P_USB_MASTER_EN_c_2, P_USB_MASTER_EN_c_1 => 
        P_USB_MASTER_EN_c_1, P_USB_MASTER_EN_c_0 => 
        P_USB_MASTER_EN_c_0, P_USB_MASTER_EN_c => 
        P_USB_MASTER_EN_c, P_MASTER_POR_B_c => P_MASTER_POR_B_c, 
        CCC_MAIN_LOCK => CCC_MAIN_LOCK, DCB_SALT_SEL_c => 
        DCB_SALT_SEL_c, DEV_RST_B_c_1 => DEV_RST_B_c_1, 
        MASTER_SALT_POR_B_i_0_i => MASTER_SALT_POR_B_i_0_i, 
        MASTER_DCB_POR_B_i_0_i => MASTER_DCB_POR_B_i_0_i, 
        MASTER_SALT_POR_B_i_0_i_0 => MASTER_SALT_POR_B_i_0_i_0, 
        MASTER_SALT_POR_B_i_0_i_1 => MASTER_SALT_POR_B_i_0_i_1, 
        MASTER_SALT_POR_B_i_0_i_2 => MASTER_SALT_POR_B_i_0_i_2, 
        MASTER_SALT_POR_B_i_0_i_3 => MASTER_SALT_POR_B_i_0_i_3, 
        MASTER_SALT_POR_B_i_0_i_4 => MASTER_SALT_POR_B_i_0_i_4, 
        MASTER_SALT_POR_B_i_0_i_5 => MASTER_SALT_POR_B_i_0_i_5, 
        MASTER_SALT_POR_B_i_0_i_6 => MASTER_SALT_POR_B_i_0_i_6, 
        MASTER_SALT_POR_B_i_0_i_7 => MASTER_SALT_POR_B_i_0_i_7, 
        MASTER_SALT_POR_B_i_0_i_8 => MASTER_SALT_POR_B_i_0_i_8, 
        MASTER_SALT_POR_B_i_0_i_9 => MASTER_SALT_POR_B_i_0_i_9, 
        MASTER_SALT_POR_B_i_0_i_10 => MASTER_SALT_POR_B_i_0_i_10, 
        MASTER_SALT_POR_B_i_0_i_11 => MASTER_SALT_POR_B_i_0_i_11, 
        MASTER_SALT_POR_B_i_0_i_12 => MASTER_SALT_POR_B_i_0_i_12, 
        MASTER_SALT_POR_B_i_0_i_13 => MASTER_SALT_POR_B_i_0_i_13, 
        MASTER_SALT_POR_B_i_0_i_14 => MASTER_SALT_POR_B_i_0_i_14, 
        MASTER_SALT_POR_B_i_0_i_15 => MASTER_SALT_POR_B_i_0_i_15, 
        MASTER_SALT_POR_B_i_0_i_16 => MASTER_SALT_POR_B_i_0_i_16, 
        MASTER_SALT_POR_B_i_0_i_17 => MASTER_SALT_POR_B_i_0_i_17, 
        P_MASTER_POR_B_c_1 => P_MASTER_POR_B_c_1, 
        P_MASTER_POR_B_c_2 => P_MASTER_POR_B_c_2, 
        P_MASTER_POR_B_c_3 => P_MASTER_POR_B_c_3, 
        P_MASTER_POR_B_c_4 => P_MASTER_POR_B_c_4, 
        P_MASTER_POR_B_c_5 => P_MASTER_POR_B_c_5, 
        P_MASTER_POR_B_c_6 => P_MASTER_POR_B_c_6, 
        P_MASTER_POR_B_c_7 => P_MASTER_POR_B_c_7, 
        P_MASTER_POR_B_c_8 => P_MASTER_POR_B_c_8, 
        P_MASTER_POR_B_c_9 => P_MASTER_POR_B_c_9, 
        P_MASTER_POR_B_c_10 => P_MASTER_POR_B_c_10, 
        P_MASTER_POR_B_c_11 => P_MASTER_POR_B_c_11, 
        P_MASTER_POR_B_c_12 => P_MASTER_POR_B_c_12, 
        P_MASTER_POR_B_c_13 => P_MASTER_POR_B_c_13, 
        P_MASTER_POR_B_c_14 => P_MASTER_POR_B_c_14, 
        P_MASTER_POR_B_c_15 => P_MASTER_POR_B_c_15, 
        P_MASTER_POR_B_c_16 => P_MASTER_POR_B_c_16, 
        P_MASTER_POR_B_c_17 => P_MASTER_POR_B_c_17, 
        P_MASTER_POR_B_c_18 => P_MASTER_POR_B_c_18, 
        P_MASTER_POR_B_c_19 => P_MASTER_POR_B_c_19, 
        P_MASTER_POR_B_c_20 => P_MASTER_POR_B_c_20, 
        P_MASTER_POR_B_c_21 => P_MASTER_POR_B_c_21, 
        P_MASTER_POR_B_c_22 => P_MASTER_POR_B_c_22, 
        P_MASTER_POR_B_c_23 => P_MASTER_POR_B_c_23, 
        P_MASTER_POR_B_c_24 => P_MASTER_POR_B_c_24, 
        P_MASTER_POR_B_c_25 => P_MASTER_POR_B_c_25, 
        P_MASTER_POR_B_c_26 => P_MASTER_POR_B_c_26, 
        P_MASTER_POR_B_c_27 => P_MASTER_POR_B_c_27, 
        P_MASTER_POR_B_c_28 => P_MASTER_POR_B_c_28, 
        P_MASTER_POR_B_c_29 => P_MASTER_POR_B_c_29, 
        P_MASTER_POR_B_c_30 => P_MASTER_POR_B_c_30, 
        P_MASTER_POR_B_c_31 => P_MASTER_POR_B_c_31, 
        P_MASTER_POR_B_c_32 => P_MASTER_POR_B_c_32, 
        P_MASTER_POR_B_c_33 => P_MASTER_POR_B_c_33, 
        P_MASTER_POR_B_c_34 => P_MASTER_POR_B_c_34, 
        P_MASTER_POR_B_c_34_0 => P_MASTER_POR_B_c_34_0, 
        P_MASTER_POR_B_c_32_0 => P_MASTER_POR_B_c_32_0, 
        P_MASTER_POR_B_c_31_0 => P_MASTER_POR_B_c_31_0, 
        P_MASTER_POR_B_c_27_0 => P_MASTER_POR_B_c_27_0, 
        P_MASTER_POR_B_c_27_1 => P_MASTER_POR_B_c_27_1, 
        P_MASTER_POR_B_c_24_0 => P_MASTER_POR_B_c_24_0, 
        P_MASTER_POR_B_c_22_0 => P_MASTER_POR_B_c_22_0, 
        P_MASTER_POR_B_c_17_0 => P_MASTER_POR_B_c_17_0, 
        P_MASTER_POR_B_c_16_0 => P_MASTER_POR_B_c_16_0, 
        DEV_RST_B_c => DEV_RST_B_c, CCC_160M_FXD => CCC_160M_FXD, 
        CLK_40M_GL => CLK_40M_GL, P_MASTER_POR_B_c_0_0 => 
        P_MASTER_POR_B_c_0_0);
    
    U_ELK7_CH : ELINK_SLAVE_15_2
      port map(BIT_OS_SEL_4(2) => \BIT_OS_SEL_4[2]\, 
        BIT_OS_SEL_4(1) => \BIT_OS_SEL_4[1]\, BIT_OS_SEL_6(2) => 
        \BIT_OS_SEL_6[2]\, BIT_OS_SEL_6(1) => \BIT_OS_SEL_6[1]\, 
        BIT_OS_SEL_5_2 => \BIT_OS_SEL_5[2]\, BIT_OS_SEL_5_0 => 
        \BIT_OS_SEL_5[0]\, BIT_OS_SEL_0 => \BIT_OS_SEL[0]\, 
        ELK_RX_SER_WORD_7(7) => \ELK_RX_SER_WORD_7[7]\, 
        ELK_RX_SER_WORD_7(6) => \ELK_RX_SER_WORD_7[6]\, 
        ELK_RX_SER_WORD_7(5) => \ELK_RX_SER_WORD_7[5]\, 
        ELK_RX_SER_WORD_7(4) => \ELK_RX_SER_WORD_7[4]\, 
        ELK_RX_SER_WORD_7(3) => \ELK_RX_SER_WORD_7[3]\, 
        ELK_RX_SER_WORD_7(2) => \ELK_RX_SER_WORD_7[2]\, 
        ELK_RX_SER_WORD_7(1) => \ELK_RX_SER_WORD_7[1]\, 
        ELK_RX_SER_WORD_7(0) => \ELK_RX_SER_WORD_7[0]\, 
        OP_MODE_c_4_0 => \OP_MODE_c_4[1]\, PATT_ELK_DAT_7(7) => 
        \PATT_ELK_DAT_7[7]\, PATT_ELK_DAT_7(6) => 
        \PATT_ELK_DAT_7[6]\, PATT_ELK_DAT_7(5) => 
        \PATT_ELK_DAT_7[5]\, PATT_ELK_DAT_7(4) => 
        \PATT_ELK_DAT_7[4]\, PATT_ELK_DAT_7(3) => 
        \PATT_ELK_DAT_7[3]\, PATT_ELK_DAT_7(2) => 
        \PATT_ELK_DAT_7[2]\, PATT_ELK_DAT_7(1) => 
        \PATT_ELK_DAT_7[1]\, PATT_ELK_DAT_7(0) => 
        \PATT_ELK_DAT_7[0]\, MASTER_DCB_POR_B_i_0_i => 
        MASTER_DCB_POR_B_i_0_i, ELK7_DAT_N => ELK7_DAT_N, 
        ELK7_DAT_P => ELK7_DAT_P, DCB_SALT_SEL_c_i => 
        DCB_SALT_SEL_c_i, CCC_160M_FXD => CCC_160M_FXD, 
        MASTER_SALT_POR_B_i_0_i_11 => MASTER_SALT_POR_B_i_0_i_11, 
        MASTER_SALT_POR_B_i_0_i_12 => MASTER_SALT_POR_B_i_0_i_12, 
        MASTER_SALT_POR_B_i_0_i_8 => MASTER_SALT_POR_B_i_0_i_8, 
        MASTER_SALT_POR_B_i_0_i_2 => MASTER_SALT_POR_B_i_0_i_2, 
        MASTER_SALT_POR_B_i_0_i_13 => MASTER_SALT_POR_B_i_0_i_13, 
        MASTER_SALT_POR_B_i_0_i_14 => MASTER_SALT_POR_B_i_0_i_14, 
        MASTER_SALT_POR_B_i_0_i_10 => MASTER_SALT_POR_B_i_0_i_10, 
        CLK_40M_GL => CLK_40M_GL, MASTER_SALT_POR_B_i_0_i_3 => 
        MASTER_SALT_POR_B_i_0_i_3, DEV_RST_B_c_1 => DEV_RST_B_c_1, 
        CCC_160M_ADJ => CCC_160M_ADJ);
    
    U_ELK14_CH : ELINK_SLAVE_15_9
      port map(BIT_OS_SEL_2(2) => \BIT_OS_SEL_2[2]\, 
        BIT_OS_SEL_2(1) => \BIT_OS_SEL_2[1]\, BIT_OS_SEL_5_0 => 
        \BIT_OS_SEL_5[2]\, BIT_OS_SEL_3_0 => \BIT_OS_SEL_3[0]\, 
        BIT_OS_SEL_4(1) => \BIT_OS_SEL_4[1]\, BIT_OS_SEL_4(0) => 
        \BIT_OS_SEL_4[0]\, ELK_RX_SER_WORD_14(7) => 
        \ELK_RX_SER_WORD_14[7]\, ELK_RX_SER_WORD_14(6) => 
        \ELK_RX_SER_WORD_14[6]\, ELK_RX_SER_WORD_14(5) => 
        \ELK_RX_SER_WORD_14[5]\, ELK_RX_SER_WORD_14(4) => 
        \ELK_RX_SER_WORD_14[4]\, ELK_RX_SER_WORD_14(3) => 
        \ELK_RX_SER_WORD_14[3]\, ELK_RX_SER_WORD_14(2) => 
        \ELK_RX_SER_WORD_14[2]\, ELK_RX_SER_WORD_14(1) => 
        \ELK_RX_SER_WORD_14[1]\, ELK_RX_SER_WORD_14(0) => 
        \ELK_RX_SER_WORD_14[0]\, OP_MODE_c_2_0 => 
        \OP_MODE_c_2[1]\, PATT_ELK_DAT_14(7) => 
        \PATT_ELK_DAT_14[7]\, PATT_ELK_DAT_14(6) => 
        \PATT_ELK_DAT_14[6]\, PATT_ELK_DAT_14(5) => 
        \PATT_ELK_DAT_14[5]\, PATT_ELK_DAT_14(4) => 
        \PATT_ELK_DAT_14[4]\, PATT_ELK_DAT_14(3) => 
        \PATT_ELK_DAT_14[3]\, PATT_ELK_DAT_14(2) => 
        \PATT_ELK_DAT_14[2]\, PATT_ELK_DAT_14(1) => 
        \PATT_ELK_DAT_14[1]\, PATT_ELK_DAT_14(0) => 
        \PATT_ELK_DAT_14[0]\, MASTER_DCB_POR_B_i_0_i => 
        MASTER_DCB_POR_B_i_0_i, ELK14_DAT_N => ELK14_DAT_N, 
        ELK14_DAT_P => ELK14_DAT_P, DCB_SALT_SEL_c_i => 
        DCB_SALT_SEL_c_i, CCC_160M_FXD => CCC_160M_FXD, 
        MASTER_SALT_POR_B_i_0_i_7 => MASTER_SALT_POR_B_i_0_i_7, 
        MASTER_SALT_POR_B_i_0_i_15 => MASTER_SALT_POR_B_i_0_i_15, 
        MASTER_SALT_POR_B_i_0_i_12 => MASTER_SALT_POR_B_i_0_i_12, 
        MASTER_SALT_POR_B_i_0_i_0 => MASTER_SALT_POR_B_i_0_i_0, 
        MASTER_SALT_POR_B_i_0_i_10 => MASTER_SALT_POR_B_i_0_i_10, 
        MASTER_SALT_POR_B_i_0_i_5 => MASTER_SALT_POR_B_i_0_i_5, 
        MASTER_SALT_POR_B_i_0_i_2 => MASTER_SALT_POR_B_i_0_i_2, 
        CLK_40M_GL => CLK_40M_GL, MASTER_SALT_POR_B_i_0_i_6 => 
        MASTER_SALT_POR_B_i_0_i_6, DEV_RST_B_c => DEV_RST_B_c, 
        CCC_160M_ADJ => CCC_160M_ADJ);
    
    U61_TS_WR_BUF : tristate_buf_0
      port map(P_USB_MASTER_EN_c => P_USB_MASTER_EN_c, USB_WR_BI
         => USB_WR_BI, USB_WR_B => USB_WR_B);
    
    P_ELK0_SYNC_DET_pad : OUTBUF
      port map(D => P_ELK0_SYNC_DET_c, PAD => P_ELK0_SYNC_DET);
    
    U_ELK2_CH : ELINK_SLAVE_15
      port map(BIT_OS_SEL_7_0 => \BIT_OS_SEL_7[2]\, BIT_OS_SEL(2)
         => \BIT_OS_SEL[2]\, BIT_OS_SEL(1) => \BIT_OS_SEL[1]\, 
        BIT_OS_SEL_0_0 => \BIT_OS_SEL_0[2]\, BIT_OS_SEL_1(1) => 
        \BIT_OS_SEL_1[1]\, BIT_OS_SEL_1(0) => \BIT_OS_SEL_1[0]\, 
        ELK_RX_SER_WORD_2(7) => \ELK_RX_SER_WORD_2[7]\, 
        ELK_RX_SER_WORD_2(6) => \ELK_RX_SER_WORD_2[6]\, 
        ELK_RX_SER_WORD_2(5) => \ELK_RX_SER_WORD_2[5]\, 
        ELK_RX_SER_WORD_2(4) => \ELK_RX_SER_WORD_2[4]\, 
        ELK_RX_SER_WORD_2(3) => \ELK_RX_SER_WORD_2[3]\, 
        ELK_RX_SER_WORD_2(2) => \ELK_RX_SER_WORD_2[2]\, 
        ELK_RX_SER_WORD_2(1) => \ELK_RX_SER_WORD_2[1]\, 
        ELK_RX_SER_WORD_2(0) => \ELK_RX_SER_WORD_2[0]\, 
        OP_MODE_c_1_0 => \OP_MODE_c_1[1]\, PATT_ELK_DAT_2(7) => 
        \PATT_ELK_DAT_2[7]\, PATT_ELK_DAT_2(6) => 
        \PATT_ELK_DAT_2[6]\, PATT_ELK_DAT_2(5) => 
        \PATT_ELK_DAT_2[5]\, PATT_ELK_DAT_2(4) => 
        \PATT_ELK_DAT_2[4]\, PATT_ELK_DAT_2(3) => 
        \PATT_ELK_DAT_2[3]\, PATT_ELK_DAT_2(2) => 
        \PATT_ELK_DAT_2[2]\, PATT_ELK_DAT_2(1) => 
        \PATT_ELK_DAT_2[1]\, PATT_ELK_DAT_2(0) => 
        \PATT_ELK_DAT_2[0]\, MASTER_DCB_POR_B_i_0_i => 
        MASTER_DCB_POR_B_i_0_i, ELK2_DAT_N => ELK2_DAT_N, 
        ELK2_DAT_P => ELK2_DAT_P, DCB_SALT_SEL_c_i => 
        DCB_SALT_SEL_c_i, CCC_160M_FXD => CCC_160M_FXD, 
        MASTER_SALT_POR_B_i_0_i_8 => MASTER_SALT_POR_B_i_0_i_8, 
        MASTER_SALT_POR_B_i_0_i_12 => MASTER_SALT_POR_B_i_0_i_12, 
        MASTER_SALT_POR_B_i_0_i_5 => MASTER_SALT_POR_B_i_0_i_5, 
        CLK_40M_GL => CLK_40M_GL, MASTER_SALT_POR_B_i_0_i_13 => 
        MASTER_SALT_POR_B_i_0_i_13, DEV_RST_B_c_0 => 
        DEV_RST_B_c_0, CCC_160M_ADJ => CCC_160M_ADJ);
    
    P_CLK_40M_GL_pad : OUTBUF
      port map(D => CLK_40M_GL, PAD => P_CLK_40M_GL);
    
    U_ELK4_CH : ELINK_SLAVE_INV_2_1
      port map(BIT_OS_SEL_7_0 => \BIT_OS_SEL_7[2]\, 
        BIT_OS_SEL_6(2) => \BIT_OS_SEL_6[2]\, BIT_OS_SEL_6(1) => 
        \BIT_OS_SEL_6[1]\, BIT_OS_SEL_0_d0 => \BIT_OS_SEL[2]\, 
        BIT_OS_SEL_0(1) => \BIT_OS_SEL_0[1]\, BIT_OS_SEL_0(0) => 
        \BIT_OS_SEL_0[0]\, BIT_OS_SEL_1_0 => \BIT_OS_SEL_1[0]\, 
        ELK_RX_SER_WORD_4(7) => \ELK_RX_SER_WORD_4[7]\, 
        ELK_RX_SER_WORD_4(6) => \ELK_RX_SER_WORD_4[6]\, 
        ELK_RX_SER_WORD_4(5) => \ELK_RX_SER_WORD_4[5]\, 
        ELK_RX_SER_WORD_4(4) => \ELK_RX_SER_WORD_4[4]\, 
        ELK_RX_SER_WORD_4(3) => \ELK_RX_SER_WORD_4[3]\, 
        ELK_RX_SER_WORD_4(2) => \ELK_RX_SER_WORD_4[2]\, 
        ELK_RX_SER_WORD_4(1) => \ELK_RX_SER_WORD_4[1]\, 
        ELK_RX_SER_WORD_4(0) => \ELK_RX_SER_WORD_4[0]\, 
        OP_MODE_c_1_0 => \OP_MODE_c_1[1]\, PATT_ELK_DAT_4(7) => 
        \PATT_ELK_DAT_4[7]\, PATT_ELK_DAT_4(6) => 
        \PATT_ELK_DAT_4[6]\, PATT_ELK_DAT_4(5) => 
        \PATT_ELK_DAT_4[5]\, PATT_ELK_DAT_4(4) => 
        \PATT_ELK_DAT_4[4]\, PATT_ELK_DAT_4(3) => 
        \PATT_ELK_DAT_4[3]\, PATT_ELK_DAT_4(2) => 
        \PATT_ELK_DAT_4[2]\, PATT_ELK_DAT_4(1) => 
        \PATT_ELK_DAT_4[1]\, PATT_ELK_DAT_4(0) => 
        \PATT_ELK_DAT_4[0]\, MASTER_DCB_POR_B_i_0_i => 
        MASTER_DCB_POR_B_i_0_i, ELK4_DAT_N => ELK4_DAT_N, 
        ELK4_DAT_P => ELK4_DAT_P, DCB_SALT_SEL_c_i => 
        DCB_SALT_SEL_c_i, CCC_160M_FXD => CCC_160M_FXD, 
        MASTER_SALT_POR_B_i_0_i_4 => MASTER_SALT_POR_B_i_0_i_4, 
        MASTER_SALT_POR_B_i_0_i_9 => MASTER_SALT_POR_B_i_0_i_9, 
        MASTER_SALT_POR_B_i_0_i_13 => MASTER_SALT_POR_B_i_0_i_13, 
        MASTER_SALT_POR_B_i_0_i_1 => MASTER_SALT_POR_B_i_0_i_1, 
        MASTER_SALT_POR_B_i_0_i_17 => MASTER_SALT_POR_B_i_0_i_17, 
        CLK_40M_GL => CLK_40M_GL, MASTER_SALT_POR_B_i_0_i_16 => 
        MASTER_SALT_POR_B_i_0_i_16, DEV_RST_B_c => DEV_RST_B_c, 
        CCC_160M_ADJ => CCC_160M_ADJ);
    
    U_DDR_TFC : DDR_BIDIR_LVDS_DUAL_CLK
      port map(DCB_SALT_SEL_c => DCB_SALT_SEL_c, TFC_DAT_0P => 
        TFC_DAT_0P, TFC_DAT_0N => TFC_DAT_0N, TFC_OUT_R => 
        TFC_OUT_R, TFC_OUT_F => TFC_OUT_F, CCC_160M_FXD => 
        CCC_160M_FXD, CCC_160M_ADJ => CCC_160M_ADJ, TFC_IN_DDR_R
         => TFC_IN_DDR_R, TFC_IN_DDR_F => TFC_IN_DDR_F);
    
    U60_TS_RD_BUF : tristate_buf
      port map(P_USB_MASTER_EN_c => P_USB_MASTER_EN_c, USB_RD_BI
         => USB_RD_BI, USB_RD_B => USB_RD_B);
    
    TFC_IN_F : DFN1C0
      port map(D => TFC_IN_DDR_F, CLK => CCC_160M_ADJ, CLR => 
        DEV_RST_B_c_0, Q => \TFC_IN_F\);
    
    U_GEN_REF_CLK : REF_CLK_DIV_GEN
      port map(DEV_RST_B_c_1 => DEV_RST_B_c_1, Y => Y, 
        CLK40M_10NS_REF => CLK40M_10NS_REF);
    
    U_ELK6_CH : ELINK_SLAVE_15_1
      port map(BIT_OS_SEL_5(2) => \BIT_OS_SEL_5[2]\, 
        BIT_OS_SEL_5(1) => \BIT_OS_SEL_5[1]\, BIT_OS_SEL_7_0 => 
        \BIT_OS_SEL_7[2]\, BIT_OS_SEL_6_0 => \BIT_OS_SEL_6[1]\, 
        BIT_OS_SEL_0 => \BIT_OS_SEL[0]\, ELK_RX_SER_WORD_6(7) => 
        \ELK_RX_SER_WORD_6[7]\, ELK_RX_SER_WORD_6(6) => 
        \ELK_RX_SER_WORD_6[6]\, ELK_RX_SER_WORD_6(5) => 
        \ELK_RX_SER_WORD_6[5]\, ELK_RX_SER_WORD_6(4) => 
        \ELK_RX_SER_WORD_6[4]\, ELK_RX_SER_WORD_6(3) => 
        \ELK_RX_SER_WORD_6[3]\, ELK_RX_SER_WORD_6(2) => 
        \ELK_RX_SER_WORD_6[2]\, ELK_RX_SER_WORD_6(1) => 
        \ELK_RX_SER_WORD_6[1]\, ELK_RX_SER_WORD_6(0) => 
        \ELK_RX_SER_WORD_6[0]\, OP_MODE_c_0_0 => \OP_MODE_c_0[1]\, 
        OP_MODE_c_1_0 => \OP_MODE_c_1[1]\, PATT_ELK_DAT_6(7) => 
        \PATT_ELK_DAT_6[7]\, PATT_ELK_DAT_6(6) => 
        \PATT_ELK_DAT_6[6]\, PATT_ELK_DAT_6(5) => 
        \PATT_ELK_DAT_6[5]\, PATT_ELK_DAT_6(4) => 
        \PATT_ELK_DAT_6[4]\, PATT_ELK_DAT_6(3) => 
        \PATT_ELK_DAT_6[3]\, PATT_ELK_DAT_6(2) => 
        \PATT_ELK_DAT_6[2]\, PATT_ELK_DAT_6(1) => 
        \PATT_ELK_DAT_6[1]\, PATT_ELK_DAT_6(0) => 
        \PATT_ELK_DAT_6[0]\, MASTER_DCB_POR_B_i_0_i => 
        MASTER_DCB_POR_B_i_0_i, ELK6_DAT_N => ELK6_DAT_N, 
        ELK6_DAT_P => ELK6_DAT_P, DCB_SALT_SEL_c_i => 
        DCB_SALT_SEL_c_i, CCC_160M_FXD => CCC_160M_FXD, 
        MASTER_SALT_POR_B_i_0_i_10 => MASTER_SALT_POR_B_i_0_i_10, 
        MASTER_SALT_POR_B_i_0_i_16 => MASTER_SALT_POR_B_i_0_i_16, 
        MASTER_SALT_POR_B_i_0_i_12 => MASTER_SALT_POR_B_i_0_i_12, 
        MASTER_SALT_POR_B_i_0_i_3 => MASTER_SALT_POR_B_i_0_i_3, 
        MASTER_SALT_POR_B_i_0_i_9 => MASTER_SALT_POR_B_i_0_i_9, 
        MASTER_SALT_POR_B_i_0_i_6 => MASTER_SALT_POR_B_i_0_i_6, 
        CLK_40M_GL => CLK_40M_GL, MASTER_SALT_POR_B_i_0_i_1 => 
        MASTER_SALT_POR_B_i_0_i_1, MASTER_SALT_POR_B_i_0_i_2 => 
        MASTER_SALT_POR_B_i_0_i_2, DEV_RST_B_c_1 => DEV_RST_B_c_1, 
        CCC_160M_ADJ => CCC_160M_ADJ);
    
    U_MASTER_DES : TOP_MASTER_DES320M
      port map(BIT_OS_SEL_7_0 => \BIT_OS_SEL_7[2]\, 
        BIT_OS_SEL_6(2) => \BIT_OS_SEL_6[2]\, BIT_OS_SEL_6(1) => 
        \BIT_OS_SEL_6[1]\, BIT_OS_SEL_5(2) => \BIT_OS_SEL_5[2]\, 
        BIT_OS_SEL_5(1) => \BIT_OS_SEL_5[1]\, BIT_OS_SEL_5(0) => 
        \BIT_OS_SEL_5[0]\, BIT_OS_SEL_4(2) => \BIT_OS_SEL_4[2]\, 
        BIT_OS_SEL_4(1) => \BIT_OS_SEL_4[1]\, BIT_OS_SEL_4(0) => 
        \BIT_OS_SEL_4[0]\, BIT_OS_SEL_3(2) => \BIT_OS_SEL_3[2]\, 
        BIT_OS_SEL_3(1) => \BIT_OS_SEL_3[1]\, BIT_OS_SEL_3(0) => 
        \BIT_OS_SEL_3[0]\, BIT_OS_SEL_2(2) => \BIT_OS_SEL_2[2]\, 
        BIT_OS_SEL_2(1) => \BIT_OS_SEL_2[1]\, BIT_OS_SEL_2(0) => 
        \BIT_OS_SEL_2[0]\, BIT_OS_SEL_1(2) => \BIT_OS_SEL_1[2]\, 
        BIT_OS_SEL_1(1) => \BIT_OS_SEL_1[1]\, BIT_OS_SEL_1(0) => 
        \BIT_OS_SEL_1[0]\, BIT_OS_SEL_0(2) => \BIT_OS_SEL_0[2]\, 
        BIT_OS_SEL_0(1) => \BIT_OS_SEL_0[1]\, BIT_OS_SEL_0(0) => 
        \BIT_OS_SEL_0[0]\, OP_MODE_c_0 => \OP_MODE_c[5]\, 
        BIT_OS_SEL(2) => \BIT_OS_SEL[2]\, BIT_OS_SEL(1) => 
        \BIT_OS_SEL[1]\, BIT_OS_SEL(0) => \BIT_OS_SEL[0]\, 
        TFC_RX_SER_WORD(7) => \TFC_RX_SER_WORD[7]\, 
        TFC_RX_SER_WORD(6) => \TFC_RX_SER_WORD[6]\, 
        TFC_RX_SER_WORD(5) => \TFC_RX_SER_WORD[5]\, 
        TFC_RX_SER_WORD(4) => \TFC_RX_SER_WORD[4]\, 
        TFC_RX_SER_WORD(3) => \TFC_RX_SER_WORD[3]\, 
        TFC_RX_SER_WORD(2) => \TFC_RX_SER_WORD[2]\, 
        TFC_RX_SER_WORD(1) => \TFC_RX_SER_WORD[1]\, 
        TFC_RX_SER_WORD(0) => \TFC_RX_SER_WORD[0]\, 
        ELK_RX_SER_WORD_0(7) => \ELK_RX_SER_WORD_0[7]\, 
        ELK_RX_SER_WORD_0(6) => \ELK_RX_SER_WORD_0[6]\, 
        ELK_RX_SER_WORD_0(5) => \ELK_RX_SER_WORD_0[5]\, 
        ELK_RX_SER_WORD_0(4) => \ELK_RX_SER_WORD_0[4]\, 
        ELK_RX_SER_WORD_0(3) => \ELK_RX_SER_WORD_0[3]\, 
        ELK_RX_SER_WORD_0(2) => \ELK_RX_SER_WORD_0[2]\, 
        ELK_RX_SER_WORD_0(1) => \ELK_RX_SER_WORD_0[1]\, 
        ELK_RX_SER_WORD_0(0) => \ELK_RX_SER_WORD_0[0]\, 
        P_MASTER_POR_B_c_27_0 => P_MASTER_POR_B_c_27_0, 
        P_MASTER_POR_B_c_27_1 => P_MASTER_POR_B_c_27_1, 
        P_MASTER_POR_B_c_16_0 => P_MASTER_POR_B_c_16_0, 
        P_MASTER_POR_B_c_17_0 => P_MASTER_POR_B_c_17_0, 
        P_MASTER_POR_B_c_24_0 => P_MASTER_POR_B_c_24_0, 
        TFC_SYNC_DET_1 => \SYNC_STAT_DET.TFC_SYNC_DET_1\, 
        ELK0_SYNC_DET_1 => \SYNC_STAT_DET.ELK0_SYNC_DET_1\, 
        DCB_SALT_SEL_c => DCB_SALT_SEL_c, TFC_IN_R => \TFC_IN_R\, 
        ELK0_IN_R => \ELK0_IN_R\, TFC_IN_F => \TFC_IN_F\, 
        ELK0_IN_F => \ELK0_IN_F\, ALL_PLL_LOCK_c => 
        ALL_PLL_LOCK_c, CCC_MAIN_LOCK => CCC_MAIN_LOCK, 
        P_MASTER_POR_B_c_31_0 => P_MASTER_POR_B_c_31_0, 
        P_MASTER_POR_B_c_26 => P_MASTER_POR_B_c_26, 
        P_MASTER_POR_B_c_32 => P_MASTER_POR_B_c_32, 
        P_MASTER_POR_B_c_24 => P_MASTER_POR_B_c_24, 
        P_MASTER_POR_B_c_5 => P_MASTER_POR_B_c_5, 
        P_MASTER_POR_B_c_4 => P_MASTER_POR_B_c_4, 
        P_MASTER_POR_B_c_2 => P_MASTER_POR_B_c_2, 
        P_MASTER_POR_B_c_3 => P_MASTER_POR_B_c_3, 
        P_MASTER_POR_B_c_9 => P_MASTER_POR_B_c_9, 
        P_MASTER_POR_B_c_21 => P_MASTER_POR_B_c_21, 
        P_MASTER_POR_B_c_15 => P_MASTER_POR_B_c_15, 
        P_MASTER_POR_B_c_16 => P_MASTER_POR_B_c_16, 
        P_MASTER_POR_B_c_12 => P_MASTER_POR_B_c_12, 
        P_MASTER_POR_B_c_11 => P_MASTER_POR_B_c_11, 
        P_MASTER_POR_B_c_7 => P_MASTER_POR_B_c_7, ALIGN_ACTIVE
         => ALIGN_ACTIVE, P_MASTER_POR_B_c_27 => 
        P_MASTER_POR_B_c_27, P_MASTER_POR_B_c_10 => 
        P_MASTER_POR_B_c_10, P_MASTER_POR_B_c_17 => 
        P_MASTER_POR_B_c_17, P_MASTER_POR_B_c_1 => 
        P_MASTER_POR_B_c_1, P_MASTER_POR_B_c_20 => 
        P_MASTER_POR_B_c_20, P_MASTER_POR_B_c_8 => 
        P_MASTER_POR_B_c_8, P_MASTER_POR_B_c_29 => 
        P_MASTER_POR_B_c_29, P_MASTER_POR_B_c_30 => 
        P_MASTER_POR_B_c_30, P_MASTER_POR_B_c_28 => 
        P_MASTER_POR_B_c_28, P_MASTER_POR_B_c_34_0 => 
        P_MASTER_POR_B_c_34_0, P_MASTER_POR_B_c_32_0 => 
        P_MASTER_POR_B_c_32_0, CCC_160M_FXD => CCC_160M_FXD, 
        P_MASTER_POR_B_c_23 => P_MASTER_POR_B_c_23, 
        P_MASTER_POR_B_c => P_MASTER_POR_B_c, CLK_40M_BUF_RECD
         => CLK_40M_BUF_RECD, CLK_40M_GL => CLK_40M_GL, 
        P_MASTER_POR_B_c_22_0 => P_MASTER_POR_B_c_22_0, 
        P_MASTER_POR_B_c_14 => P_MASTER_POR_B_c_14, 
        P_MASTER_POR_B_c_6 => P_MASTER_POR_B_c_6, 
        P_MASTER_POR_B_c_25 => P_MASTER_POR_B_c_25, 
        P_MASTER_POR_B_c_13 => P_MASTER_POR_B_c_13, 
        P_MASTER_POR_B_c_22 => P_MASTER_POR_B_c_22, 
        P_MASTER_POR_B_c_31 => P_MASTER_POR_B_c_31, 
        P_MASTER_POR_B_c_33 => P_MASTER_POR_B_c_33, 
        P_MASTER_POR_B_c_18 => P_MASTER_POR_B_c_18, 
        P_MASTER_POR_B_c_19 => P_MASTER_POR_B_c_19, 
        P_MASTER_POR_B_c_34 => P_MASTER_POR_B_c_34, CCC_160M_ADJ
         => CCC_160M_ADJ);
    
    U_ELK16_CH : ELINK_SLAVE_15_11
      port map(BIT_OS_SEL_1(2) => \BIT_OS_SEL_1[2]\, 
        BIT_OS_SEL_1(1) => \BIT_OS_SEL_1[1]\, BIT_OS_SEL_2_0 => 
        \BIT_OS_SEL_2[1]\, BIT_OS_SEL_3(2) => \BIT_OS_SEL_3[2]\, 
        BIT_OS_SEL_3(1) => \BIT_OS_SEL_3[1]\, BIT_OS_SEL_3(0) => 
        \BIT_OS_SEL_3[0]\, ELK_RX_SER_WORD_16(7) => 
        \ELK_RX_SER_WORD_16[7]\, ELK_RX_SER_WORD_16(6) => 
        \ELK_RX_SER_WORD_16[6]\, ELK_RX_SER_WORD_16(5) => 
        \ELK_RX_SER_WORD_16[5]\, ELK_RX_SER_WORD_16(4) => 
        \ELK_RX_SER_WORD_16[4]\, ELK_RX_SER_WORD_16(3) => 
        \ELK_RX_SER_WORD_16[3]\, ELK_RX_SER_WORD_16(2) => 
        \ELK_RX_SER_WORD_16[2]\, ELK_RX_SER_WORD_16(1) => 
        \ELK_RX_SER_WORD_16[1]\, ELK_RX_SER_WORD_16(0) => 
        \ELK_RX_SER_WORD_16[0]\, OP_MODE_c_2_0 => 
        \OP_MODE_c_2[1]\, PATT_ELK_DAT_16(7) => 
        \PATT_ELK_DAT_16[7]\, PATT_ELK_DAT_16(6) => 
        \PATT_ELK_DAT_16[6]\, PATT_ELK_DAT_16(5) => 
        \PATT_ELK_DAT_16[5]\, PATT_ELK_DAT_16(4) => 
        \PATT_ELK_DAT_16[4]\, PATT_ELK_DAT_16(3) => 
        \PATT_ELK_DAT_16[3]\, PATT_ELK_DAT_16(2) => 
        \PATT_ELK_DAT_16[2]\, PATT_ELK_DAT_16(1) => 
        \PATT_ELK_DAT_16[1]\, PATT_ELK_DAT_16(0) => 
        \PATT_ELK_DAT_16[0]\, MASTER_DCB_POR_B_i_0_i => 
        MASTER_DCB_POR_B_i_0_i, ELK16_DAT_N => ELK16_DAT_N, 
        ELK16_DAT_P => ELK16_DAT_P, DCB_SALT_SEL_c_i => 
        DCB_SALT_SEL_c_i, CCC_160M_FXD => CCC_160M_FXD, 
        MASTER_SALT_POR_B_i_0_i_8 => MASTER_SALT_POR_B_i_0_i_8, 
        MASTER_SALT_POR_B_i_0_i_1 => MASTER_SALT_POR_B_i_0_i_1, 
        MASTER_SALT_POR_B_i_0_i_16 => MASTER_SALT_POR_B_i_0_i_16, 
        MASTER_SALT_POR_B_i_0_i_0 => MASTER_SALT_POR_B_i_0_i_0, 
        MASTER_SALT_POR_B_i_0_i_10 => MASTER_SALT_POR_B_i_0_i_10, 
        MASTER_SALT_POR_B_i_0_i_14 => MASTER_SALT_POR_B_i_0_i_14, 
        CLK_40M_GL => CLK_40M_GL, MASTER_SALT_POR_B_i_0_i_9 => 
        MASTER_SALT_POR_B_i_0_i_9, DEV_RST_B_c_1 => DEV_RST_B_c_1, 
        CCC_160M_ADJ => CCC_160M_ADJ);
    
    U63_TS_SIWU_BUF : tristate_buf_2
      port map(P_USB_MASTER_EN_c => P_USB_MASTER_EN_c, 
        USB_SIWU_BI => USB_SIWU_BI, USB_SIWU_B => USB_SIWU_B);
    
    P_OP_MODE2_TE_pad : OUTBUF
      port map(D => \OP_MODE_c[2]\, PAD => P_OP_MODE2_TE);
    
    P_OP_MODE5_AAE_pad : OUTBUF
      port map(D => \OP_MODE_c[5]\, PAD => P_OP_MODE5_AAE);
    
    ELK0_IN_R : DFN1C0
      port map(D => ELK0_IN_DDR_R_i, CLK => CCC_160M_ADJ, CLR => 
        DEV_RST_B_c, Q => \ELK0_IN_R\);
    
    DCB_SALT_SEL_pad_RNIJM3B : INV
      port map(A => DCB_SALT_SEL_c, Y => DCB_SALT_SEL_c_i);
    
    U_DDR_ELK0 : DDR_BIDIR_LVDS_DUAL_CLK_0
      port map(DCB_SALT_SEL_c_i => DCB_SALT_SEL_c_i, ELK0_DAT_P
         => ELK0_DAT_P, ELK0_DAT_N => ELK0_DAT_N, ELK0_OUT_R_i_0
         => ELK0_OUT_R_i_0, ELK0_OUT_F_i_0 => ELK0_OUT_F_i_0, 
        CCC_160M_FXD => CCC_160M_FXD, CCC_160M_ADJ => 
        CCC_160M_ADJ, ELK0_IN_DDR_F_i => ELK0_IN_DDR_F_i, 
        ELK0_IN_DDR_R_i => ELK0_IN_DDR_R_i);
    
    P_USB_MASTER_EN_pad : OUTBUF
      port map(D => P_USB_MASTER_EN_c, PAD => P_USB_MASTER_EN);
    
    U0_200M_BUF : LVDS_CLK_IN
      port map(CLK200_N => CLK200_N, CLK200_P => CLK200_P, Y => Y);
    
    ELK0_SYNC_DET : DFN1C0
      port map(D => \SYNC_STAT_DET.ELK0_SYNC_DET_1\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_25, Q => 
        P_ELK0_SYNC_DET_c);
    
    U_ELK19_CH : ELINK_SLAVE_15_14
      port map(BIT_OS_SEL_0_d0 => \BIT_OS_SEL[2]\, 
        BIT_OS_SEL_0(2) => \BIT_OS_SEL_0[2]\, BIT_OS_SEL_0(1) => 
        \BIT_OS_SEL_0[1]\, BIT_OS_SEL_1(2) => \BIT_OS_SEL_1[2]\, 
        BIT_OS_SEL_1(1) => \BIT_OS_SEL_1[1]\, BIT_OS_SEL_2_0 => 
        \BIT_OS_SEL_2[0]\, ELK_RX_SER_WORD_19(7) => 
        \ELK_RX_SER_WORD_19[7]\, ELK_RX_SER_WORD_19(6) => 
        \ELK_RX_SER_WORD_19[6]\, ELK_RX_SER_WORD_19(5) => 
        \ELK_RX_SER_WORD_19[5]\, ELK_RX_SER_WORD_19(4) => 
        \ELK_RX_SER_WORD_19[4]\, ELK_RX_SER_WORD_19(3) => 
        \ELK_RX_SER_WORD_19[3]\, ELK_RX_SER_WORD_19(2) => 
        \ELK_RX_SER_WORD_19[2]\, ELK_RX_SER_WORD_19(1) => 
        \ELK_RX_SER_WORD_19[1]\, ELK_RX_SER_WORD_19(0) => 
        \ELK_RX_SER_WORD_19[0]\, OP_MODE_c_5_0 => 
        \OP_MODE_c_5[1]\, OP_MODE_c_6_0 => \OP_MODE_c_6[1]\, 
        PATT_ELK_DAT_19(7) => \PATT_ELK_DAT_19[7]\, 
        PATT_ELK_DAT_19(6) => \PATT_ELK_DAT_19[6]\, 
        PATT_ELK_DAT_19(5) => \PATT_ELK_DAT_19[5]\, 
        PATT_ELK_DAT_19(4) => \PATT_ELK_DAT_19[4]\, 
        PATT_ELK_DAT_19(3) => \PATT_ELK_DAT_19[3]\, 
        PATT_ELK_DAT_19(2) => \PATT_ELK_DAT_19[2]\, 
        PATT_ELK_DAT_19(1) => \PATT_ELK_DAT_19[1]\, 
        PATT_ELK_DAT_19(0) => \PATT_ELK_DAT_19[0]\, 
        MASTER_DCB_POR_B_i_0_i => MASTER_DCB_POR_B_i_0_i, 
        ELK19_DAT_N => ELK19_DAT_N, ELK19_DAT_P => ELK19_DAT_P, 
        DCB_SALT_SEL_c_i => DCB_SALT_SEL_c_i, CCC_160M_FXD => 
        CCC_160M_FXD, MASTER_SALT_POR_B_i_0_i_10 => 
        MASTER_SALT_POR_B_i_0_i_10, MASTER_SALT_POR_B_i_0_i_16
         => MASTER_SALT_POR_B_i_0_i_16, 
        MASTER_SALT_POR_B_i_0_i_12 => MASTER_SALT_POR_B_i_0_i_12, 
        MASTER_SALT_POR_B_i_0_i_8 => MASTER_SALT_POR_B_i_0_i_8, 
        MASTER_SALT_POR_B_i_0_i_0 => MASTER_SALT_POR_B_i_0_i_0, 
        MASTER_SALT_POR_B_i_0_i_7 => MASTER_SALT_POR_B_i_0_i_7, 
        MASTER_SALT_POR_B_i_0_i_4 => MASTER_SALT_POR_B_i_0_i_4, 
        CLK_40M_GL => CLK_40M_GL, MASTER_SALT_POR_B_i_0_i_15 => 
        MASTER_SALT_POR_B_i_0_i_15, DEV_RST_B_c_0 => 
        DEV_RST_B_c_0, CCC_160M_ADJ => CCC_160M_ADJ);
    
    U_ELK9_CH : ELINK_SLAVE_15_4
      port map(BIT_OS_SEL_2(2) => \BIT_OS_SEL_2[2]\, 
        BIT_OS_SEL_2(1) => \BIT_OS_SEL_2[1]\, BIT_OS_SEL_3(2) => 
        \BIT_OS_SEL_3[2]\, BIT_OS_SEL_3(1) => \BIT_OS_SEL_3[1]\, 
        BIT_OS_SEL_5(2) => \BIT_OS_SEL_5[2]\, BIT_OS_SEL_5(1) => 
        \BIT_OS_SEL_5[1]\, BIT_OS_SEL_4_0 => \BIT_OS_SEL_4[0]\, 
        ELK_RX_SER_WORD_9(7) => \ELK_RX_SER_WORD_9[7]\, 
        ELK_RX_SER_WORD_9(6) => \ELK_RX_SER_WORD_9[6]\, 
        ELK_RX_SER_WORD_9(5) => \ELK_RX_SER_WORD_9[5]\, 
        ELK_RX_SER_WORD_9(4) => \ELK_RX_SER_WORD_9[4]\, 
        ELK_RX_SER_WORD_9(3) => \ELK_RX_SER_WORD_9[3]\, 
        ELK_RX_SER_WORD_9(2) => \ELK_RX_SER_WORD_9[2]\, 
        ELK_RX_SER_WORD_9(1) => \ELK_RX_SER_WORD_9[1]\, 
        ELK_RX_SER_WORD_9(0) => \ELK_RX_SER_WORD_9[0]\, 
        OP_MODE_c_3_0 => \OP_MODE_c_3[1]\, PATT_ELK_DAT_9(7) => 
        \PATT_ELK_DAT_9[7]\, PATT_ELK_DAT_9(6) => 
        \PATT_ELK_DAT_9[6]\, PATT_ELK_DAT_9(5) => 
        \PATT_ELK_DAT_9[5]\, PATT_ELK_DAT_9(4) => 
        \PATT_ELK_DAT_9[4]\, PATT_ELK_DAT_9(3) => 
        \PATT_ELK_DAT_9[3]\, PATT_ELK_DAT_9(2) => 
        \PATT_ELK_DAT_9[2]\, PATT_ELK_DAT_9(1) => 
        \PATT_ELK_DAT_9[1]\, PATT_ELK_DAT_9(0) => 
        \PATT_ELK_DAT_9[0]\, MASTER_DCB_POR_B_i_0_i => 
        MASTER_DCB_POR_B_i_0_i, ELK9_DAT_N => ELK9_DAT_N, 
        ELK9_DAT_P => ELK9_DAT_P, DCB_SALT_SEL_c_i => 
        DCB_SALT_SEL_c_i, CCC_160M_FXD => CCC_160M_FXD, 
        MASTER_SALT_POR_B_i_0_i_12 => MASTER_SALT_POR_B_i_0_i_12, 
        MASTER_SALT_POR_B_i_0_i_16 => MASTER_SALT_POR_B_i_0_i_16, 
        MASTER_SALT_POR_B_i_0_i_13 => MASTER_SALT_POR_B_i_0_i_13, 
        MASTER_SALT_POR_B_i_0_i_2 => MASTER_SALT_POR_B_i_0_i_2, 
        MASTER_SALT_POR_B_i_0_i_3 => MASTER_SALT_POR_B_i_0_i_3, 
        MASTER_SALT_POR_B_i_0_i_4 => MASTER_SALT_POR_B_i_0_i_4, 
        MASTER_SALT_POR_B_i_0_i_0 => MASTER_SALT_POR_B_i_0_i_0, 
        CLK_40M_GL => CLK_40M_GL, MASTER_SALT_POR_B_i_0_i_7 => 
        MASTER_SALT_POR_B_i_0_i_7, DEV_RST_B_c_0 => DEV_RST_B_c_0, 
        CCC_160M_ADJ => CCC_160M_ADJ);
    
    DCB_SALT_SEL_pad : INBUF
      port map(PAD => DCB_SALT_SEL, Y => DCB_SALT_SEL_c);
    
    P_TFC_SYNC_DET_pad : OUTBUF
      port map(D => P_TFC_SYNC_DET_c, PAD => P_TFC_SYNC_DET);
    
    U200A_TFC : GP_PATT_GEN_1
      port map(TFC_ADDRB(7) => \TFC_ADDRB[7]\, TFC_ADDRB(6) => 
        \TFC_ADDRB[6]\, TFC_ADDRB(5) => \TFC_ADDRB[5]\, 
        TFC_ADDRB(4) => \TFC_ADDRB[4]\, TFC_ADDRB(3) => 
        \TFC_ADDRB[3]\, TFC_ADDRB(2) => \TFC_ADDRB[2]\, 
        TFC_ADDRB(1) => \TFC_ADDRB[1]\, TFC_ADDRB(0) => 
        \TFC_ADDRB[0]\, TFC_RX_SER_WORD(7) => 
        \TFC_RX_SER_WORD[7]\, TFC_RX_SER_WORD(6) => 
        \TFC_RX_SER_WORD[6]\, TFC_RX_SER_WORD(5) => 
        \TFC_RX_SER_WORD[5]\, TFC_RX_SER_WORD(4) => 
        \TFC_RX_SER_WORD[4]\, TFC_RX_SER_WORD(3) => 
        \TFC_RX_SER_WORD[3]\, TFC_RX_SER_WORD(2) => 
        \TFC_RX_SER_WORD[2]\, TFC_RX_SER_WORD(1) => 
        \TFC_RX_SER_WORD[1]\, TFC_RX_SER_WORD(0) => 
        \TFC_RX_SER_WORD[0]\, TFC_STOP_ADDR(7) => 
        \TFC_STOP_ADDR[7]\, TFC_STOP_ADDR(6) => 
        \TFC_STOP_ADDR[6]\, TFC_STOP_ADDR(5) => 
        \TFC_STOP_ADDR[5]\, TFC_STOP_ADDR(4) => 
        \TFC_STOP_ADDR[4]\, TFC_STOP_ADDR(3) => 
        \TFC_STOP_ADDR[3]\, TFC_STOP_ADDR(2) => 
        \TFC_STOP_ADDR[2]\, TFC_STOP_ADDR(1) => 
        \TFC_STOP_ADDR[1]\, TFC_STOP_ADDR(0) => 
        \TFC_STOP_ADDR[0]\, TFC_STRT_ADDR(7) => 
        \TFC_STRT_ADDR[7]\, TFC_STRT_ADDR(6) => 
        \TFC_STRT_ADDR[6]\, TFC_STRT_ADDR(5) => 
        \TFC_STRT_ADDR[5]\, TFC_STRT_ADDR(4) => 
        \TFC_STRT_ADDR[4]\, TFC_STRT_ADDR(3) => 
        \TFC_STRT_ADDR[3]\, TFC_STRT_ADDR(2) => 
        \TFC_STRT_ADDR[2]\, TFC_STRT_ADDR(1) => 
        \TFC_STRT_ADDR[1]\, TFC_STRT_ADDR(0) => 
        \TFC_STRT_ADDR[0]\, OP_MODE_0 => \OP_MODE[0]\, 
        OP_MODE_c_0 => \OP_MODE_c[2]\, P_MASTER_POR_B_c_24 => 
        P_MASTER_POR_B_c_24, P_MASTER_POR_B_c => P_MASTER_POR_B_c, 
        P_MASTER_POR_B_c_31 => P_MASTER_POR_B_c_31, 
        P_MASTER_POR_B_c_30 => P_MASTER_POR_B_c_30, 
        P_MASTER_POR_B_c_1 => P_MASTER_POR_B_c_1, 
        P_MASTER_POR_B_c_5 => P_MASTER_POR_B_c_5, 
        P_MASTER_POR_B_c_4 => P_MASTER_POR_B_c_4, 
        P_MASTER_POR_B_c_28 => P_MASTER_POR_B_c_28, 
        DCB_SALT_SEL_c => DCB_SALT_SEL_c, P_MASTER_POR_B_c_15 => 
        P_MASTER_POR_B_c_15, P_MASTER_POR_B_c_16_0 => 
        P_MASTER_POR_B_c_16_0, TFC_RWB => TFC_RWB, 
        P_MASTER_POR_B_c_9 => P_MASTER_POR_B_c_9, TFC_RAM_BLKB_EN
         => TFC_RAM_BLKB_EN, P_USB_MASTER_EN_c_22_0 => 
        P_USB_MASTER_EN_c_22_0, ALIGN_ACTIVE => ALIGN_ACTIVE, 
        P_MASTER_POR_B_c_27_1 => P_MASTER_POR_B_c_27_1, 
        CLK_40M_GL => CLK_40M_GL);
    
    U_ELK8_CH : ELINK_SLAVE_15_3
      port map(BIT_OS_SEL_4_0 => \BIT_OS_SEL_4[2]\, 
        BIT_OS_SEL_3(2) => \BIT_OS_SEL_3[2]\, BIT_OS_SEL_3(1) => 
        \BIT_OS_SEL_3[1]\, BIT_OS_SEL_6_0 => \BIT_OS_SEL_6[2]\, 
        BIT_OS_SEL_5(1) => \BIT_OS_SEL_5[1]\, BIT_OS_SEL_5(0) => 
        \BIT_OS_SEL_5[0]\, ELK_RX_SER_WORD_8(7) => 
        \ELK_RX_SER_WORD_8[7]\, ELK_RX_SER_WORD_8(6) => 
        \ELK_RX_SER_WORD_8[6]\, ELK_RX_SER_WORD_8(5) => 
        \ELK_RX_SER_WORD_8[5]\, ELK_RX_SER_WORD_8(4) => 
        \ELK_RX_SER_WORD_8[4]\, ELK_RX_SER_WORD_8(3) => 
        \ELK_RX_SER_WORD_8[3]\, ELK_RX_SER_WORD_8(2) => 
        \ELK_RX_SER_WORD_8[2]\, ELK_RX_SER_WORD_8(1) => 
        \ELK_RX_SER_WORD_8[1]\, ELK_RX_SER_WORD_8(0) => 
        \ELK_RX_SER_WORD_8[0]\, OP_MODE_c_0_0 => \OP_MODE_c_0[1]\, 
        PATT_ELK_DAT_8(7) => \PATT_ELK_DAT_8[7]\, 
        PATT_ELK_DAT_8(6) => \PATT_ELK_DAT_8[6]\, 
        PATT_ELK_DAT_8(5) => \PATT_ELK_DAT_8[5]\, 
        PATT_ELK_DAT_8(4) => \PATT_ELK_DAT_8[4]\, 
        PATT_ELK_DAT_8(3) => \PATT_ELK_DAT_8[3]\, 
        PATT_ELK_DAT_8(2) => \PATT_ELK_DAT_8[2]\, 
        PATT_ELK_DAT_8(1) => \PATT_ELK_DAT_8[1]\, 
        PATT_ELK_DAT_8(0) => \PATT_ELK_DAT_8[0]\, 
        MASTER_DCB_POR_B_i_0_i => MASTER_DCB_POR_B_i_0_i, 
        ELK8_DAT_N => ELK8_DAT_N, ELK8_DAT_P => ELK8_DAT_P, 
        DCB_SALT_SEL_c_i => DCB_SALT_SEL_c_i, CCC_160M_FXD => 
        CCC_160M_FXD, MASTER_SALT_POR_B_i_0_i_12 => 
        MASTER_SALT_POR_B_i_0_i_12, MASTER_SALT_POR_B_i_0_i_2 => 
        MASTER_SALT_POR_B_i_0_i_2, MASTER_SALT_POR_B_i_0_i_3 => 
        MASTER_SALT_POR_B_i_0_i_3, MASTER_SALT_POR_B_i_0_i => 
        MASTER_SALT_POR_B_i_0_i, MASTER_SALT_POR_B_i_0_i_15 => 
        MASTER_SALT_POR_B_i_0_i_15, CLK_40M_GL => CLK_40M_GL, 
        MASTER_SALT_POR_B_i_0_i_5 => MASTER_SALT_POR_B_i_0_i_5, 
        DEV_RST_B_c_1 => DEV_RST_B_c_1, DEV_RST_B_c_0 => 
        DEV_RST_B_c_0, CCC_160M_ADJ => CCC_160M_ADJ);
    
    U_ELK17_CH : ELINK_SLAVE_15_12
      port map(BIT_OS_SEL_0_0 => \BIT_OS_SEL_0[2]\, 
        BIT_OS_SEL_1_0 => \BIT_OS_SEL_1[1]\, BIT_OS_SEL_2(2) => 
        \BIT_OS_SEL_2[2]\, BIT_OS_SEL_2(1) => \BIT_OS_SEL_2[1]\, 
        BIT_OS_SEL_2(0) => \BIT_OS_SEL_2[0]\, BIT_OS_SEL_3_0 => 
        \BIT_OS_SEL_3[0]\, ELK_RX_SER_WORD_17(7) => 
        \ELK_RX_SER_WORD_17[7]\, ELK_RX_SER_WORD_17(6) => 
        \ELK_RX_SER_WORD_17[6]\, ELK_RX_SER_WORD_17(5) => 
        \ELK_RX_SER_WORD_17[5]\, ELK_RX_SER_WORD_17(4) => 
        \ELK_RX_SER_WORD_17[4]\, ELK_RX_SER_WORD_17(3) => 
        \ELK_RX_SER_WORD_17[3]\, ELK_RX_SER_WORD_17(2) => 
        \ELK_RX_SER_WORD_17[2]\, ELK_RX_SER_WORD_17(1) => 
        \ELK_RX_SER_WORD_17[1]\, ELK_RX_SER_WORD_17(0) => 
        \ELK_RX_SER_WORD_17[0]\, OP_MODE_c_6_0 => 
        \OP_MODE_c_6[1]\, PATT_ELK_DAT_17(7) => 
        \PATT_ELK_DAT_17[7]\, PATT_ELK_DAT_17(6) => 
        \PATT_ELK_DAT_17[6]\, PATT_ELK_DAT_17(5) => 
        \PATT_ELK_DAT_17[5]\, PATT_ELK_DAT_17(4) => 
        \PATT_ELK_DAT_17[4]\, PATT_ELK_DAT_17(3) => 
        \PATT_ELK_DAT_17[3]\, PATT_ELK_DAT_17(2) => 
        \PATT_ELK_DAT_17[2]\, PATT_ELK_DAT_17(1) => 
        \PATT_ELK_DAT_17[1]\, PATT_ELK_DAT_17(0) => 
        \PATT_ELK_DAT_17[0]\, MASTER_DCB_POR_B_i_0_i => 
        MASTER_DCB_POR_B_i_0_i, ELK17_DAT_N => ELK17_DAT_N, 
        ELK17_DAT_P => ELK17_DAT_P, DCB_SALT_SEL_c_i => 
        DCB_SALT_SEL_c_i, CCC_160M_FXD => CCC_160M_FXD, 
        MASTER_SALT_POR_B_i_0_i_9 => MASTER_SALT_POR_B_i_0_i_9, 
        MASTER_SALT_POR_B_i_0_i_8 => MASTER_SALT_POR_B_i_0_i_8, 
        MASTER_SALT_POR_B_i_0_i_0 => MASTER_SALT_POR_B_i_0_i_0, 
        MASTER_SALT_POR_B_i_0_i_17 => MASTER_SALT_POR_B_i_0_i_17, 
        MASTER_SALT_POR_B_i_0_i_14 => MASTER_SALT_POR_B_i_0_i_14, 
        CLK_40M_GL => CLK_40M_GL, MASTER_SALT_POR_B_i_0_i_11 => 
        MASTER_SALT_POR_B_i_0_i_11, MASTER_SALT_POR_B_i_0_i_12
         => MASTER_SALT_POR_B_i_0_i_12, DEV_RST_B_c_1 => 
        DEV_RST_B_c_1, CCC_160M_ADJ => CCC_160M_ADJ);
    
    U_ELK15_CH : ELINK_SLAVE_15_10
      port map(BIT_OS_SEL_1_0 => \BIT_OS_SEL_1[2]\, 
        BIT_OS_SEL_2(2) => \BIT_OS_SEL_2[2]\, BIT_OS_SEL_2(1) => 
        \BIT_OS_SEL_2[1]\, BIT_OS_SEL_4_0 => \BIT_OS_SEL_4[2]\, 
        BIT_OS_SEL_3(1) => \BIT_OS_SEL_3[1]\, BIT_OS_SEL_3(0) => 
        \BIT_OS_SEL_3[0]\, ELK_RX_SER_WORD_15(7) => 
        \ELK_RX_SER_WORD_15[7]\, ELK_RX_SER_WORD_15(6) => 
        \ELK_RX_SER_WORD_15[6]\, ELK_RX_SER_WORD_15(5) => 
        \ELK_RX_SER_WORD_15[5]\, ELK_RX_SER_WORD_15(4) => 
        \ELK_RX_SER_WORD_15[4]\, ELK_RX_SER_WORD_15(3) => 
        \ELK_RX_SER_WORD_15[3]\, ELK_RX_SER_WORD_15(2) => 
        \ELK_RX_SER_WORD_15[2]\, ELK_RX_SER_WORD_15(1) => 
        \ELK_RX_SER_WORD_15[1]\, ELK_RX_SER_WORD_15(0) => 
        \ELK_RX_SER_WORD_15[0]\, OP_MODE_c_6_0 => 
        \OP_MODE_c_6[1]\, PATT_ELK_DAT_15(7) => 
        \PATT_ELK_DAT_15[7]\, PATT_ELK_DAT_15(6) => 
        \PATT_ELK_DAT_15[6]\, PATT_ELK_DAT_15(5) => 
        \PATT_ELK_DAT_15[5]\, PATT_ELK_DAT_15(4) => 
        \PATT_ELK_DAT_15[4]\, PATT_ELK_DAT_15(3) => 
        \PATT_ELK_DAT_15[3]\, PATT_ELK_DAT_15(2) => 
        \PATT_ELK_DAT_15[2]\, PATT_ELK_DAT_15(1) => 
        \PATT_ELK_DAT_15[1]\, PATT_ELK_DAT_15(0) => 
        \PATT_ELK_DAT_15[0]\, MASTER_DCB_POR_B_i_0_i => 
        MASTER_DCB_POR_B_i_0_i, ELK15_DAT_N => ELK15_DAT_N, 
        ELK15_DAT_P => ELK15_DAT_P, DCB_SALT_SEL_c_i => 
        DCB_SALT_SEL_c_i, CCC_160M_FXD => CCC_160M_FXD, 
        MASTER_SALT_POR_B_i_0_i_5 => MASTER_SALT_POR_B_i_0_i_5, 
        MASTER_SALT_POR_B_i_0_i_9 => MASTER_SALT_POR_B_i_0_i_9, 
        MASTER_SALT_POR_B_i_0_i_1 => MASTER_SALT_POR_B_i_0_i_1, 
        MASTER_SALT_POR_B_i_0_i_6 => MASTER_SALT_POR_B_i_0_i_6, 
        CLK_40M_GL => CLK_40M_GL, MASTER_SALT_POR_B_i_0_i_7 => 
        MASTER_SALT_POR_B_i_0_i_7, MASTER_SALT_POR_B_i_0_i_8 => 
        MASTER_SALT_POR_B_i_0_i_8, DEV_RST_B_c_1 => DEV_RST_B_c_1, 
        CCC_160M_ADJ => CCC_160M_ADJ);
    
    U0A_40M_REFCLK : BIDIR_LVDS_IO
      port map(EXT_INT_REF_SEL_c => EXT_INT_REF_SEL_c, 
        CLK40M_10NS_REF => CLK40M_10NS_REF, CLK_40M_BUF_RECD => 
        CLK_40M_BUF_RECD, BIDIR_CLK40M_P => BIDIR_CLK40M_P, 
        BIDIR_CLK40M_N => BIDIR_CLK40M_N);
    
    U0B_TX40M_REFCLK : LVDS_BUFOUT
      port map(CLK_40M_BUF_RECD => CLK_40M_BUF_RECD, TX_CLK40M_P
         => TX_CLK40M_P, TX_CLK40M_N => TX_CLK40M_N);
    
    P_OP_MODE1_SPE_pad : OUTBUF
      port map(D => \OP_MODE_c[1]\, PAD => P_OP_MODE1_SPE);
    
    U_ELK5_CH : ELINK_SLAVE_15_0
      port map(BIT_OS_SEL_5(2) => \BIT_OS_SEL_5[2]\, 
        BIT_OS_SEL_5(1) => \BIT_OS_SEL_5[1]\, BIT_OS_SEL_6(2) => 
        \BIT_OS_SEL_6[2]\, BIT_OS_SEL_6(1) => \BIT_OS_SEL_6[1]\, 
        BIT_OS_SEL_7_0 => \BIT_OS_SEL_7[2]\, BIT_OS_SEL_0_d0 => 
        \BIT_OS_SEL[1]\, BIT_OS_SEL_0_0 => \BIT_OS_SEL_0[0]\, 
        ELK_RX_SER_WORD_5(7) => \ELK_RX_SER_WORD_5[7]\, 
        ELK_RX_SER_WORD_5(6) => \ELK_RX_SER_WORD_5[6]\, 
        ELK_RX_SER_WORD_5(5) => \ELK_RX_SER_WORD_5[5]\, 
        ELK_RX_SER_WORD_5(4) => \ELK_RX_SER_WORD_5[4]\, 
        ELK_RX_SER_WORD_5(3) => \ELK_RX_SER_WORD_5[3]\, 
        ELK_RX_SER_WORD_5(2) => \ELK_RX_SER_WORD_5[2]\, 
        ELK_RX_SER_WORD_5(1) => \ELK_RX_SER_WORD_5[1]\, 
        ELK_RX_SER_WORD_5(0) => \ELK_RX_SER_WORD_5[0]\, 
        OP_MODE_c_4_0 => \OP_MODE_c_4[1]\, OP_MODE_c_5_0 => 
        \OP_MODE_c_5[1]\, PATT_ELK_DAT_5(7) => 
        \PATT_ELK_DAT_5[7]\, PATT_ELK_DAT_5(6) => 
        \PATT_ELK_DAT_5[6]\, PATT_ELK_DAT_5(5) => 
        \PATT_ELK_DAT_5[5]\, PATT_ELK_DAT_5(4) => 
        \PATT_ELK_DAT_5[4]\, PATT_ELK_DAT_5(3) => 
        \PATT_ELK_DAT_5[3]\, PATT_ELK_DAT_5(2) => 
        \PATT_ELK_DAT_5[2]\, PATT_ELK_DAT_5(1) => 
        \PATT_ELK_DAT_5[1]\, PATT_ELK_DAT_5(0) => 
        \PATT_ELK_DAT_5[0]\, MASTER_DCB_POR_B_i_0_i => 
        MASTER_DCB_POR_B_i_0_i, ELK5_DAT_N => ELK5_DAT_N, 
        ELK5_DAT_P => ELK5_DAT_P, DCB_SALT_SEL_c_i => 
        DCB_SALT_SEL_c_i, CCC_160M_FXD => CCC_160M_FXD, 
        MASTER_SALT_POR_B_i_0_i_9 => MASTER_SALT_POR_B_i_0_i_9, 
        MASTER_SALT_POR_B_i_0_i_8 => MASTER_SALT_POR_B_i_0_i_8, 
        MASTER_SALT_POR_B_i_0_i_5 => MASTER_SALT_POR_B_i_0_i_5, 
        MASTER_SALT_POR_B_i_0_i_3 => MASTER_SALT_POR_B_i_0_i_3, 
        MASTER_SALT_POR_B_i_0_i_14 => MASTER_SALT_POR_B_i_0_i_14, 
        MASTER_SALT_POR_B_i_0_i_6 => MASTER_SALT_POR_B_i_0_i_6, 
        MASTER_SALT_POR_B_i_0_i_2 => MASTER_SALT_POR_B_i_0_i_2, 
        CLK_40M_GL => CLK_40M_GL, MASTER_SALT_POR_B_i_0_i_17 => 
        MASTER_SALT_POR_B_i_0_i_17, MASTER_SALT_POR_B_i_0_i => 
        MASTER_SALT_POR_B_i_0_i, DEV_RST_B_c => DEV_RST_B_c, 
        CCC_160M_ADJ => CCC_160M_ADJ);
    
    U_ELK10_CH : ELINK_SLAVE_15_5
      port map(BIT_OS_SEL_6_0 => \BIT_OS_SEL_6[2]\, 
        BIT_OS_SEL_5(2) => \BIT_OS_SEL_5[2]\, BIT_OS_SEL_5(1) => 
        \BIT_OS_SEL_5[1]\, BIT_OS_SEL_7_0 => \BIT_OS_SEL_7[2]\, 
        BIT_OS_SEL_0_d0 => \BIT_OS_SEL[1]\, BIT_OS_SEL_0_0 => 
        \BIT_OS_SEL_0[0]\, ELK_RX_SER_WORD_10(7) => 
        \ELK_RX_SER_WORD_10[7]\, ELK_RX_SER_WORD_10(6) => 
        \ELK_RX_SER_WORD_10[6]\, ELK_RX_SER_WORD_10(5) => 
        \ELK_RX_SER_WORD_10[5]\, ELK_RX_SER_WORD_10(4) => 
        \ELK_RX_SER_WORD_10[4]\, ELK_RX_SER_WORD_10(3) => 
        \ELK_RX_SER_WORD_10[3]\, ELK_RX_SER_WORD_10(2) => 
        \ELK_RX_SER_WORD_10[2]\, ELK_RX_SER_WORD_10(1) => 
        \ELK_RX_SER_WORD_10[1]\, ELK_RX_SER_WORD_10(0) => 
        \ELK_RX_SER_WORD_10[0]\, OP_MODE_c_3_0 => 
        \OP_MODE_c_3[1]\, PATT_ELK_DAT_10(7) => 
        \PATT_ELK_DAT_10[7]\, PATT_ELK_DAT_10(6) => 
        \PATT_ELK_DAT_10[6]\, PATT_ELK_DAT_10(5) => 
        \PATT_ELK_DAT_10[5]\, PATT_ELK_DAT_10(4) => 
        \PATT_ELK_DAT_10[4]\, PATT_ELK_DAT_10(3) => 
        \PATT_ELK_DAT_10[3]\, PATT_ELK_DAT_10(2) => 
        \PATT_ELK_DAT_10[2]\, PATT_ELK_DAT_10(1) => 
        \PATT_ELK_DAT_10[1]\, PATT_ELK_DAT_10(0) => 
        \PATT_ELK_DAT_10[0]\, MASTER_DCB_POR_B_i_0_i => 
        MASTER_DCB_POR_B_i_0_i, ELK10_DAT_N => ELK10_DAT_N, 
        ELK10_DAT_P => ELK10_DAT_P, DCB_SALT_SEL_c_i => 
        DCB_SALT_SEL_c_i, CCC_160M_FXD => CCC_160M_FXD, 
        MASTER_SALT_POR_B_i_0_i_5 => MASTER_SALT_POR_B_i_0_i_5, 
        MASTER_SALT_POR_B_i_0_i_8 => MASTER_SALT_POR_B_i_0_i_8, 
        MASTER_SALT_POR_B_i_0_i_1 => MASTER_SALT_POR_B_i_0_i_1, 
        MASTER_SALT_POR_B_i_0_i_11 => MASTER_SALT_POR_B_i_0_i_11, 
        MASTER_SALT_POR_B_i_0_i_6 => MASTER_SALT_POR_B_i_0_i_6, 
        MASTER_SALT_POR_B_i_0_i_3 => MASTER_SALT_POR_B_i_0_i_3, 
        CLK_40M_GL => CLK_40M_GL, MASTER_SALT_POR_B_i_0_i_17 => 
        MASTER_SALT_POR_B_i_0_i_17, DEV_RST_B_c_0 => 
        DEV_RST_B_c_0, CCC_160M_ADJ => CCC_160M_ADJ);
    
    EXTCLK_40MHZ_pad : OUTBUF
      port map(D => EXTCLK_40MHZ_c, PAD => EXTCLK_40MHZ);
    

end DEF_ARCH; 
