-- Version: v11.7 11.7.0.119
-- File used only for Simulation

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity TOP_COMET is

    port( CLK200_P        : in    std_logic;
          CLK200_N        : in    std_logic;
          DEV_RST_B       : in    std_logic;
          DCB_SALT_SEL    : in    std_logic;
          EXTCLK_40MHZ    : out   std_logic;
          EXT_INT_REF_SEL : in    std_logic;
          ALL_PLL_LOCK    : out   std_logic;
          P_MASTER_POR_B  : out   std_logic;
          P_USB_MASTER_EN : out   std_logic;
          P_CLK_40M_GL    : out   std_logic;
          P_CCC_160M_FXD  : out   std_logic;
          P_CCC_160M_ADJ  : out   std_logic;
          P_ELK0_SYNC_DET : out   std_logic;
          P_TFC_SYNC_DET  : out   std_logic;
          P_OP_MODE1_SPE  : out   std_logic;
          P_OP_MODE2_TE   : out   std_logic;
          P_OP_MODE5_AAE  : out   std_logic;
          P_OP_MODE6_EE   : out   std_logic;
          BIDIR_CLK40M_P  : inout std_logic := 'Z';
          BIDIR_CLK40M_N  : inout std_logic := 'Z';
          TX_CLK40M_P     : out   std_logic;
          TX_CLK40M_N     : out   std_logic;
          USBCLK60MHZ     : in    std_logic;
          BIDIR_USB_ADBUS : inout std_logic_vector(7 downto 0) := (others => 'Z');
          USB_OE_B        : out   std_logic;
          P_USB_RXF_B     : in    std_logic;
          USB_RD_B        : out   std_logic;
          P_USB_TXE_B     : in    std_logic;
          USB_WR_B        : out   std_logic;
          USB_SIWU_B      : out   std_logic;
          TFC_DAT_0P      : inout std_logic := 'Z';
          TFC_DAT_0N      : inout std_logic := 'Z';
          REF_CLK_0P      : inout std_logic := 'Z';
          REF_CLK_0N      : inout std_logic := 'Z';
          ELK0_DAT_P      : inout std_logic := 'Z';
          ELK0_DAT_N      : inout std_logic := 'Z';
          ELK1_DAT_P      : inout std_logic := 'Z';
          ELK1_DAT_N      : inout std_logic := 'Z';
          ELK2_DAT_P      : inout std_logic := 'Z';
          ELK2_DAT_N      : inout std_logic := 'Z';
          ELK3_DAT_P      : inout std_logic := 'Z';
          ELK3_DAT_N      : inout std_logic := 'Z';
          ELK4_DAT_P      : inout std_logic := 'Z';
          ELK4_DAT_N      : inout std_logic := 'Z';
          ELK5_DAT_P      : inout std_logic := 'Z';
          ELK5_DAT_N      : inout std_logic := 'Z';
          ELK6_DAT_P      : inout std_logic := 'Z';
          ELK6_DAT_N      : inout std_logic := 'Z';
          ELK7_DAT_P      : inout std_logic := 'Z';
          ELK7_DAT_N      : inout std_logic := 'Z';
          ELK8_DAT_P      : inout std_logic := 'Z';
          ELK8_DAT_N      : inout std_logic := 'Z';
          ELK9_DAT_P      : inout std_logic := 'Z';
          ELK9_DAT_N      : inout std_logic := 'Z';
          ELK10_DAT_P     : inout std_logic := 'Z';
          ELK10_DAT_N     : inout std_logic := 'Z';
          ELK11_DAT_P     : inout std_logic := 'Z';
          ELK11_DAT_N     : inout std_logic := 'Z';
          ELK12_DAT_P     : inout std_logic := 'Z';
          ELK12_DAT_N     : inout std_logic := 'Z';
          ELK13_DAT_P     : inout std_logic := 'Z';
          ELK13_DAT_N     : inout std_logic := 'Z';
          ELK14_DAT_P     : inout std_logic := 'Z';
          ELK14_DAT_N     : inout std_logic := 'Z';
          ELK15_DAT_P     : inout std_logic := 'Z';
          ELK15_DAT_N     : inout std_logic := 'Z';
          ELK16_DAT_P     : inout std_logic := 'Z';
          ELK16_DAT_N     : inout std_logic := 'Z';
          ELK17_DAT_P     : inout std_logic := 'Z';
          ELK17_DAT_N     : inout std_logic := 'Z';
          ELK18_DAT_P     : inout std_logic := 'Z';
          ELK18_DAT_N     : inout std_logic := 'Z';
          ELK19_DAT_P     : inout std_logic := 'Z';
          ELK19_DAT_N     : inout std_logic := 'Z'
        );

end TOP_COMET;

architecture DEF_ARCH of TOP_COMET is 

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component IOIN_IB
    port( YIN : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component AND3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1D
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NAND2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component IOBI_ID_OD_EB
    port( DR   : in    std_logic := 'U';
          DF   : in    std_logic := 'U';
          CLR  : in    std_logic := 'U';
          E    : in    std_logic := 'U';
          ICLK : in    std_logic := 'U';
          OCLK : in    std_logic := 'U';
          YIN  : in    std_logic := 'U';
          DOUT : out   std_logic;
          EOUT : out   std_logic;
          YR   : out   std_logic;
          YF   : out   std_logic
        );
  end component;

  component AOI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component INV
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XNOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XO1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NAND2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component IOBI_IRC_OB_EB
    port( D    : in    std_logic := 'U';
          CLR  : in    std_logic := 'U';
          E    : in    std_logic := 'U';
          ICLK : in    std_logic := 'U';
          YIN  : in    std_logic := 'U';
          DOUT : out   std_logic;
          EOUT : out   std_logic;
          Y    : out   std_logic
        );
  end component;

  component AO1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component IOPAD_TRI_U
    port( D   : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          PAD : out   std_logic
        );
  end component;

  component NAND3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NAND2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFI1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          QN  : out   std_logic
        );
  end component;

  component DFN1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component XA1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NAND3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1D
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NAND3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XO1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component IOPADP_BI
    port( N2PIN : in    std_logic := 'U';
          D     : in    std_logic := 'U';
          E     : in    std_logic := 'U';
          PAD   : inout   std_logic;
          Y     : out   std_logic
        );
  end component;

  component NAND3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component IOTRI_OB_EB
    port( D    : in    std_logic := 'U';
          E    : in    std_logic := 'U';
          DOUT : out   std_logic;
          EOUT : out   std_logic
        );
  end component;

  component XA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component RAM4K9
    generic (MEMORYFILE:string := "");

    port( ADDRA11 : in    std_logic := 'U';
          ADDRA10 : in    std_logic := 'U';
          ADDRA9  : in    std_logic := 'U';
          ADDRA8  : in    std_logic := 'U';
          ADDRA7  : in    std_logic := 'U';
          ADDRA6  : in    std_logic := 'U';
          ADDRA5  : in    std_logic := 'U';
          ADDRA4  : in    std_logic := 'U';
          ADDRA3  : in    std_logic := 'U';
          ADDRA2  : in    std_logic := 'U';
          ADDRA1  : in    std_logic := 'U';
          ADDRA0  : in    std_logic := 'U';
          ADDRB11 : in    std_logic := 'U';
          ADDRB10 : in    std_logic := 'U';
          ADDRB9  : in    std_logic := 'U';
          ADDRB8  : in    std_logic := 'U';
          ADDRB7  : in    std_logic := 'U';
          ADDRB6  : in    std_logic := 'U';
          ADDRB5  : in    std_logic := 'U';
          ADDRB4  : in    std_logic := 'U';
          ADDRB3  : in    std_logic := 'U';
          ADDRB2  : in    std_logic := 'U';
          ADDRB1  : in    std_logic := 'U';
          ADDRB0  : in    std_logic := 'U';
          DINA8   : in    std_logic := 'U';
          DINA7   : in    std_logic := 'U';
          DINA6   : in    std_logic := 'U';
          DINA5   : in    std_logic := 'U';
          DINA4   : in    std_logic := 'U';
          DINA3   : in    std_logic := 'U';
          DINA2   : in    std_logic := 'U';
          DINA1   : in    std_logic := 'U';
          DINA0   : in    std_logic := 'U';
          DINB8   : in    std_logic := 'U';
          DINB7   : in    std_logic := 'U';
          DINB6   : in    std_logic := 'U';
          DINB5   : in    std_logic := 'U';
          DINB4   : in    std_logic := 'U';
          DINB3   : in    std_logic := 'U';
          DINB2   : in    std_logic := 'U';
          DINB1   : in    std_logic := 'U';
          DINB0   : in    std_logic := 'U';
          WIDTHA0 : in    std_logic := 'U';
          WIDTHA1 : in    std_logic := 'U';
          WIDTHB0 : in    std_logic := 'U';
          WIDTHB1 : in    std_logic := 'U';
          PIPEA   : in    std_logic := 'U';
          PIPEB   : in    std_logic := 'U';
          WMODEA  : in    std_logic := 'U';
          WMODEB  : in    std_logic := 'U';
          BLKA    : in    std_logic := 'U';
          BLKB    : in    std_logic := 'U';
          WENA    : in    std_logic := 'U';
          WENB    : in    std_logic := 'U';
          CLKA    : in    std_logic := 'U';
          CLKB    : in    std_logic := 'U';
          RESET   : in    std_logic := 'U';
          DOUTA8  : out   std_logic;
          DOUTA7  : out   std_logic;
          DOUTA6  : out   std_logic;
          DOUTA5  : out   std_logic;
          DOUTA4  : out   std_logic;
          DOUTA3  : out   std_logic;
          DOUTA2  : out   std_logic;
          DOUTA1  : out   std_logic;
          DOUTA0  : out   std_logic;
          DOUTB8  : out   std_logic;
          DOUTB7  : out   std_logic;
          DOUTB6  : out   std_logic;
          DOUTB5  : out   std_logic;
          DOUTB4  : out   std_logic;
          DOUTB3  : out   std_logic;
          DOUTB2  : out   std_logic;
          DOUTB1  : out   std_logic;
          DOUTB0  : out   std_logic
        );
  end component;

  component AO18
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component IOPADN_BI
    port( DB     : in    std_logic := 'U';
          E      : in    std_logic := 'U';
          PAD    : inout   std_logic;
          N2POUT : out   std_logic
        );
  end component;

  component NOR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DYNCCC
    generic (VCOFREQUENCY:real := 0.0);

    port( CLKA      : in    std_logic := 'U';
          EXTFB     : in    std_logic := 'U';
          POWERDOWN : in    std_logic := 'U';
          GLA       : out   std_logic;
          LOCK      : out   std_logic;
          CLKB      : in    std_logic := 'U';
          GLB       : out   std_logic;
          YB        : out   std_logic;
          CLKC      : in    std_logic := 'U';
          GLC       : out   std_logic;
          YC        : out   std_logic;
          SDIN      : in    std_logic := 'U';
          SCLK      : in    std_logic := 'U';
          SSHIFT    : in    std_logic := 'U';
          SUPDATE   : in    std_logic := 'U';
          MODE      : in    std_logic := 'U';
          SDOUT     : out   std_logic;
          OADIV0    : in    std_logic := 'U';
          OADIV1    : in    std_logic := 'U';
          OADIV2    : in    std_logic := 'U';
          OADIV3    : in    std_logic := 'U';
          OADIV4    : in    std_logic := 'U';
          OAMUX0    : in    std_logic := 'U';
          OAMUX1    : in    std_logic := 'U';
          OAMUX2    : in    std_logic := 'U';
          DLYGLA0   : in    std_logic := 'U';
          DLYGLA1   : in    std_logic := 'U';
          DLYGLA2   : in    std_logic := 'U';
          DLYGLA3   : in    std_logic := 'U';
          DLYGLA4   : in    std_logic := 'U';
          OBDIV0    : in    std_logic := 'U';
          OBDIV1    : in    std_logic := 'U';
          OBDIV2    : in    std_logic := 'U';
          OBDIV3    : in    std_logic := 'U';
          OBDIV4    : in    std_logic := 'U';
          OBMUX0    : in    std_logic := 'U';
          OBMUX1    : in    std_logic := 'U';
          OBMUX2    : in    std_logic := 'U';
          DLYYB0    : in    std_logic := 'U';
          DLYYB1    : in    std_logic := 'U';
          DLYYB2    : in    std_logic := 'U';
          DLYYB3    : in    std_logic := 'U';
          DLYYB4    : in    std_logic := 'U';
          DLYGLB0   : in    std_logic := 'U';
          DLYGLB1   : in    std_logic := 'U';
          DLYGLB2   : in    std_logic := 'U';
          DLYGLB3   : in    std_logic := 'U';
          DLYGLB4   : in    std_logic := 'U';
          OCDIV0    : in    std_logic := 'U';
          OCDIV1    : in    std_logic := 'U';
          OCDIV2    : in    std_logic := 'U';
          OCDIV3    : in    std_logic := 'U';
          OCDIV4    : in    std_logic := 'U';
          OCMUX0    : in    std_logic := 'U';
          OCMUX1    : in    std_logic := 'U';
          OCMUX2    : in    std_logic := 'U';
          DLYYC0    : in    std_logic := 'U';
          DLYYC1    : in    std_logic := 'U';
          DLYYC2    : in    std_logic := 'U';
          DLYYC3    : in    std_logic := 'U';
          DLYYC4    : in    std_logic := 'U';
          DLYGLC0   : in    std_logic := 'U';
          DLYGLC1   : in    std_logic := 'U';
          DLYGLC2   : in    std_logic := 'U';
          DLYGLC3   : in    std_logic := 'U';
          DLYGLC4   : in    std_logic := 'U';
          FINDIV0   : in    std_logic := 'U';
          FINDIV1   : in    std_logic := 'U';
          FINDIV2   : in    std_logic := 'U';
          FINDIV3   : in    std_logic := 'U';
          FINDIV4   : in    std_logic := 'U';
          FINDIV5   : in    std_logic := 'U';
          FINDIV6   : in    std_logic := 'U';
          FBDIV0    : in    std_logic := 'U';
          FBDIV1    : in    std_logic := 'U';
          FBDIV2    : in    std_logic := 'U';
          FBDIV3    : in    std_logic := 'U';
          FBDIV4    : in    std_logic := 'U';
          FBDIV5    : in    std_logic := 'U';
          FBDIV6    : in    std_logic := 'U';
          FBDLY0    : in    std_logic := 'U';
          FBDLY1    : in    std_logic := 'U';
          FBDLY2    : in    std_logic := 'U';
          FBDLY3    : in    std_logic := 'U';
          FBDLY4    : in    std_logic := 'U';
          FBSEL0    : in    std_logic := 'U';
          FBSEL1    : in    std_logic := 'U';
          XDLYSEL   : in    std_logic := 'U';
          VCOSEL0   : in    std_logic := 'U';
          VCOSEL1   : in    std_logic := 'U';
          VCOSEL2   : in    std_logic := 'U'
        );
  end component;

  component IOPAD_BI_U
    port( D   : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Y   : out   std_logic;
          PAD : inout   std_logic
        );
  end component;

  component IOPAD_IN_U
    port( PAD : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component AX1E
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO13
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component IOBI_IB_OB_EB
    port( D    : in    std_logic := 'U';
          E    : in    std_logic := 'U';
          YIN  : in    std_logic := 'U';
          DOUT : out   std_logic;
          EOUT : out   std_logic;
          Y    : out   std_logic
        );
  end component;

  component DFI1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          QN  : out   std_logic
        );
  end component;

  component AO1E
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AXOI4
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AXOI3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component IOPADP_TRI
    port( D   : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          PAD : out   std_logic
        );
  end component;

  component AX1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component IOPADN_IN
    port( PAD    : in    std_logic := 'U';
          N2POUT : out   std_logic
        );
  end component;

  component AXOI7
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AXOI5
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XNOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component IOIN_IRP
    port( PRE  : in    std_logic := 'U';
          ICLK : in    std_logic := 'U';
          YIN  : in    std_logic := 'U';
          Y    : out   std_logic
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component IOPAD_IN
    port( PAD : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component IOPADN_OUT
    port( DB  : in    std_logic := 'U';
          PAD : out   std_logic
        );
  end component;

  component IOPADP_IN
    port( N2PIN : in    std_logic := 'U';
          PAD   : in    std_logic := 'U';
          Y     : out   std_logic
        );
  end component;

  component GND
    port(Y : out std_logic); 
  end component;

  component VCC
    port(Y : out std_logic); 
  end component;

    signal Y, CLK40M_10NS_REF, CLK_40M_BUF_RECD, CCC_MAIN_LOCK, 
        CLK60MHZ, \PATT_TFC_DAT[0]\, \PATT_TFC_DAT[1]\, 
        \PATT_TFC_DAT[2]\, \PATT_TFC_DAT[3]\, \PATT_TFC_DAT[4]\, 
        \PATT_TFC_DAT[5]\, \PATT_TFC_DAT[6]\, \PATT_TFC_DAT[7]\, 
        \TFC_TX_DAT[0]\, \TFC_TX_DAT[1]\, \TFC_TX_DAT[2]\, 
        \TFC_TX_DAT[3]\, \TFC_TX_DAT[4]\, \TFC_TX_DAT[5]\, 
        \TFC_TX_DAT[6]\, \TFC_TX_DAT[7]\, TFC_OUT_R, TFC_OUT_F, 
        TFC_IN_DDR_R, TFC_IN_DDR_F, \PATT_ELK_DAT_0[0]\, 
        \PATT_ELK_DAT_0[1]\, \PATT_ELK_DAT_0[2]\, 
        \PATT_ELK_DAT_0[3]\, \PATT_ELK_DAT_0[4]\, 
        \PATT_ELK_DAT_0[5]\, \PATT_ELK_DAT_0[6]\, 
        \PATT_ELK_DAT_0[7]\, \TFC_RX_SER_WORD[0]\, 
        \TFC_RX_SER_WORD[1]\, \TFC_RX_SER_WORD[2]\, 
        \TFC_RX_SER_WORD[3]\, \TFC_RX_SER_WORD[4]\, 
        \TFC_RX_SER_WORD[5]\, \TFC_RX_SER_WORD[6]\, 
        \TFC_RX_SER_WORD[7]\, \ELK_RX_SER_WORD_0[0]\, 
        \ELK_RX_SER_WORD_0[1]\, \ELK_RX_SER_WORD_0[2]\, 
        \ELK_RX_SER_WORD_0[3]\, \ELK_RX_SER_WORD_0[4]\, 
        \ELK_RX_SER_WORD_0[5]\, \ELK_RX_SER_WORD_0[6]\, 
        \ELK_RX_SER_WORD_0[7]\, \PATT_ELK_DAT_1[0]\, 
        \PATT_ELK_DAT_1[1]\, \PATT_ELK_DAT_1[2]\, 
        \PATT_ELK_DAT_1[3]\, \PATT_ELK_DAT_1[4]\, 
        \PATT_ELK_DAT_1[5]\, \PATT_ELK_DAT_1[6]\, 
        \PATT_ELK_DAT_1[7]\, \ELK_RX_SER_WORD_1[0]\, 
        \ELK_RX_SER_WORD_1[1]\, \ELK_RX_SER_WORD_1[2]\, 
        \ELK_RX_SER_WORD_1[3]\, \ELK_RX_SER_WORD_1[4]\, 
        \ELK_RX_SER_WORD_1[5]\, \ELK_RX_SER_WORD_1[6]\, 
        \ELK_RX_SER_WORD_1[7]\, \PATT_ELK_DAT_2[0]\, 
        \PATT_ELK_DAT_2[1]\, \PATT_ELK_DAT_2[2]\, 
        \PATT_ELK_DAT_2[3]\, \PATT_ELK_DAT_2[4]\, 
        \PATT_ELK_DAT_2[5]\, \PATT_ELK_DAT_2[6]\, 
        \PATT_ELK_DAT_2[7]\, \ELK_RX_SER_WORD_2[0]\, 
        \ELK_RX_SER_WORD_2[1]\, \ELK_RX_SER_WORD_2[2]\, 
        \ELK_RX_SER_WORD_2[3]\, \ELK_RX_SER_WORD_2[4]\, 
        \ELK_RX_SER_WORD_2[5]\, \ELK_RX_SER_WORD_2[6]\, 
        \ELK_RX_SER_WORD_2[7]\, \PATT_ELK_DAT_3[0]\, 
        \PATT_ELK_DAT_3[1]\, \PATT_ELK_DAT_3[2]\, 
        \PATT_ELK_DAT_3[3]\, \PATT_ELK_DAT_3[4]\, 
        \PATT_ELK_DAT_3[5]\, \PATT_ELK_DAT_3[6]\, 
        \PATT_ELK_DAT_3[7]\, \ELK_RX_SER_WORD_3[0]\, 
        \ELK_RX_SER_WORD_3[1]\, \ELK_RX_SER_WORD_3[2]\, 
        \ELK_RX_SER_WORD_3[3]\, \ELK_RX_SER_WORD_3[4]\, 
        \ELK_RX_SER_WORD_3[5]\, \ELK_RX_SER_WORD_3[6]\, 
        \ELK_RX_SER_WORD_3[7]\, \PATT_ELK_DAT_4[0]\, 
        \PATT_ELK_DAT_4[1]\, \PATT_ELK_DAT_4[2]\, 
        \PATT_ELK_DAT_4[3]\, \PATT_ELK_DAT_4[4]\, 
        \PATT_ELK_DAT_4[5]\, \PATT_ELK_DAT_4[6]\, 
        \PATT_ELK_DAT_4[7]\, \ELK_RX_SER_WORD_4[0]\, 
        \ELK_RX_SER_WORD_4[1]\, \ELK_RX_SER_WORD_4[2]\, 
        \ELK_RX_SER_WORD_4[3]\, \ELK_RX_SER_WORD_4[4]\, 
        \ELK_RX_SER_WORD_4[5]\, \ELK_RX_SER_WORD_4[6]\, 
        \ELK_RX_SER_WORD_4[7]\, \PATT_ELK_DAT_5[0]\, 
        \PATT_ELK_DAT_5[1]\, \PATT_ELK_DAT_5[2]\, 
        \PATT_ELK_DAT_5[3]\, \PATT_ELK_DAT_5[4]\, 
        \PATT_ELK_DAT_5[5]\, \PATT_ELK_DAT_5[6]\, 
        \PATT_ELK_DAT_5[7]\, \ELK_RX_SER_WORD_5[0]\, 
        \ELK_RX_SER_WORD_5[1]\, \ELK_RX_SER_WORD_5[2]\, 
        \ELK_RX_SER_WORD_5[3]\, \ELK_RX_SER_WORD_5[4]\, 
        \ELK_RX_SER_WORD_5[5]\, \ELK_RX_SER_WORD_5[6]\, 
        \ELK_RX_SER_WORD_5[7]\, \PATT_ELK_DAT_6[0]\, 
        \PATT_ELK_DAT_6[1]\, \PATT_ELK_DAT_6[2]\, 
        \PATT_ELK_DAT_6[3]\, \PATT_ELK_DAT_6[4]\, 
        \PATT_ELK_DAT_6[5]\, \PATT_ELK_DAT_6[6]\, 
        \PATT_ELK_DAT_6[7]\, \ELK_RX_SER_WORD_6[0]\, 
        \ELK_RX_SER_WORD_6[1]\, \ELK_RX_SER_WORD_6[2]\, 
        \ELK_RX_SER_WORD_6[3]\, \ELK_RX_SER_WORD_6[4]\, 
        \ELK_RX_SER_WORD_6[5]\, \ELK_RX_SER_WORD_6[6]\, 
        \ELK_RX_SER_WORD_6[7]\, \PATT_ELK_DAT_7[0]\, 
        \PATT_ELK_DAT_7[1]\, \PATT_ELK_DAT_7[2]\, 
        \PATT_ELK_DAT_7[3]\, \PATT_ELK_DAT_7[4]\, 
        \PATT_ELK_DAT_7[5]\, \PATT_ELK_DAT_7[6]\, 
        \PATT_ELK_DAT_7[7]\, \ELK_RX_SER_WORD_7[0]\, 
        \ELK_RX_SER_WORD_7[1]\, \ELK_RX_SER_WORD_7[2]\, 
        \ELK_RX_SER_WORD_7[3]\, \ELK_RX_SER_WORD_7[4]\, 
        \ELK_RX_SER_WORD_7[5]\, \ELK_RX_SER_WORD_7[6]\, 
        \ELK_RX_SER_WORD_7[7]\, \PATT_ELK_DAT_8[0]\, 
        \PATT_ELK_DAT_8[1]\, \PATT_ELK_DAT_8[2]\, 
        \PATT_ELK_DAT_8[3]\, \PATT_ELK_DAT_8[4]\, 
        \PATT_ELK_DAT_8[5]\, \PATT_ELK_DAT_8[6]\, 
        \PATT_ELK_DAT_8[7]\, \ELK_RX_SER_WORD_8[0]\, 
        \ELK_RX_SER_WORD_8[1]\, \ELK_RX_SER_WORD_8[2]\, 
        \ELK_RX_SER_WORD_8[3]\, \ELK_RX_SER_WORD_8[4]\, 
        \ELK_RX_SER_WORD_8[5]\, \ELK_RX_SER_WORD_8[6]\, 
        \ELK_RX_SER_WORD_8[7]\, \PATT_ELK_DAT_9[0]\, 
        \PATT_ELK_DAT_9[1]\, \PATT_ELK_DAT_9[2]\, 
        \PATT_ELK_DAT_9[3]\, \PATT_ELK_DAT_9[4]\, 
        \PATT_ELK_DAT_9[5]\, \PATT_ELK_DAT_9[6]\, 
        \PATT_ELK_DAT_9[7]\, \ELK_RX_SER_WORD_9[0]\, 
        \ELK_RX_SER_WORD_9[1]\, \ELK_RX_SER_WORD_9[2]\, 
        \ELK_RX_SER_WORD_9[3]\, \ELK_RX_SER_WORD_9[4]\, 
        \ELK_RX_SER_WORD_9[5]\, \ELK_RX_SER_WORD_9[6]\, 
        \ELK_RX_SER_WORD_9[7]\, \PATT_ELK_DAT_10[0]\, 
        \PATT_ELK_DAT_10[1]\, \PATT_ELK_DAT_10[2]\, 
        \PATT_ELK_DAT_10[3]\, \PATT_ELK_DAT_10[4]\, 
        \PATT_ELK_DAT_10[5]\, \PATT_ELK_DAT_10[6]\, 
        \PATT_ELK_DAT_10[7]\, \ELK_RX_SER_WORD_10[0]\, 
        \ELK_RX_SER_WORD_10[1]\, \ELK_RX_SER_WORD_10[2]\, 
        \ELK_RX_SER_WORD_10[3]\, \ELK_RX_SER_WORD_10[4]\, 
        \ELK_RX_SER_WORD_10[5]\, \ELK_RX_SER_WORD_10[6]\, 
        \ELK_RX_SER_WORD_10[7]\, \PATT_ELK_DAT_11[0]\, 
        \PATT_ELK_DAT_11[1]\, \PATT_ELK_DAT_11[2]\, 
        \PATT_ELK_DAT_11[3]\, \PATT_ELK_DAT_11[4]\, 
        \PATT_ELK_DAT_11[5]\, \PATT_ELK_DAT_11[6]\, 
        \PATT_ELK_DAT_11[7]\, \ELK_RX_SER_WORD_11[0]\, 
        \ELK_RX_SER_WORD_11[1]\, \ELK_RX_SER_WORD_11[2]\, 
        \ELK_RX_SER_WORD_11[3]\, \ELK_RX_SER_WORD_11[4]\, 
        \ELK_RX_SER_WORD_11[5]\, \ELK_RX_SER_WORD_11[6]\, 
        \ELK_RX_SER_WORD_11[7]\, \PATT_ELK_DAT_12[0]\, 
        \PATT_ELK_DAT_12[1]\, \PATT_ELK_DAT_12[2]\, 
        \PATT_ELK_DAT_12[3]\, \PATT_ELK_DAT_12[4]\, 
        \PATT_ELK_DAT_12[5]\, \PATT_ELK_DAT_12[6]\, 
        \PATT_ELK_DAT_12[7]\, \ELK_RX_SER_WORD_12[0]\, 
        \ELK_RX_SER_WORD_12[1]\, \ELK_RX_SER_WORD_12[2]\, 
        \ELK_RX_SER_WORD_12[3]\, \ELK_RX_SER_WORD_12[4]\, 
        \ELK_RX_SER_WORD_12[5]\, \ELK_RX_SER_WORD_12[6]\, 
        \ELK_RX_SER_WORD_12[7]\, \PATT_ELK_DAT_13[0]\, 
        \PATT_ELK_DAT_13[1]\, \PATT_ELK_DAT_13[2]\, 
        \PATT_ELK_DAT_13[3]\, \PATT_ELK_DAT_13[4]\, 
        \PATT_ELK_DAT_13[5]\, \PATT_ELK_DAT_13[6]\, 
        \PATT_ELK_DAT_13[7]\, \ELK_RX_SER_WORD_13[0]\, 
        \ELK_RX_SER_WORD_13[1]\, \ELK_RX_SER_WORD_13[2]\, 
        \ELK_RX_SER_WORD_13[3]\, \ELK_RX_SER_WORD_13[4]\, 
        \ELK_RX_SER_WORD_13[5]\, \ELK_RX_SER_WORD_13[6]\, 
        \ELK_RX_SER_WORD_13[7]\, \PATT_ELK_DAT_14[0]\, 
        \PATT_ELK_DAT_14[1]\, \PATT_ELK_DAT_14[2]\, 
        \PATT_ELK_DAT_14[3]\, \PATT_ELK_DAT_14[4]\, 
        \PATT_ELK_DAT_14[5]\, \PATT_ELK_DAT_14[6]\, 
        \PATT_ELK_DAT_14[7]\, \ELK_RX_SER_WORD_14[0]\, 
        \ELK_RX_SER_WORD_14[1]\, \ELK_RX_SER_WORD_14[2]\, 
        \ELK_RX_SER_WORD_14[3]\, \ELK_RX_SER_WORD_14[4]\, 
        \ELK_RX_SER_WORD_14[5]\, \ELK_RX_SER_WORD_14[6]\, 
        \ELK_RX_SER_WORD_14[7]\, \PATT_ELK_DAT_15[0]\, 
        \PATT_ELK_DAT_15[1]\, \PATT_ELK_DAT_15[2]\, 
        \PATT_ELK_DAT_15[3]\, \PATT_ELK_DAT_15[4]\, 
        \PATT_ELK_DAT_15[5]\, \PATT_ELK_DAT_15[6]\, 
        \PATT_ELK_DAT_15[7]\, \ELK_RX_SER_WORD_15[0]\, 
        \ELK_RX_SER_WORD_15[1]\, \ELK_RX_SER_WORD_15[2]\, 
        \ELK_RX_SER_WORD_15[3]\, \ELK_RX_SER_WORD_15[4]\, 
        \ELK_RX_SER_WORD_15[5]\, \ELK_RX_SER_WORD_15[6]\, 
        \ELK_RX_SER_WORD_15[7]\, \PATT_ELK_DAT_16[0]\, 
        \PATT_ELK_DAT_16[1]\, \PATT_ELK_DAT_16[2]\, 
        \PATT_ELK_DAT_16[3]\, \PATT_ELK_DAT_16[4]\, 
        \PATT_ELK_DAT_16[5]\, \PATT_ELK_DAT_16[6]\, 
        \PATT_ELK_DAT_16[7]\, \ELK_RX_SER_WORD_16[0]\, 
        \ELK_RX_SER_WORD_16[1]\, \ELK_RX_SER_WORD_16[2]\, 
        \ELK_RX_SER_WORD_16[3]\, \ELK_RX_SER_WORD_16[4]\, 
        \ELK_RX_SER_WORD_16[5]\, \ELK_RX_SER_WORD_16[6]\, 
        \ELK_RX_SER_WORD_16[7]\, \PATT_ELK_DAT_17[0]\, 
        \PATT_ELK_DAT_17[1]\, \PATT_ELK_DAT_17[2]\, 
        \PATT_ELK_DAT_17[3]\, \PATT_ELK_DAT_17[4]\, 
        \PATT_ELK_DAT_17[5]\, \PATT_ELK_DAT_17[6]\, 
        \PATT_ELK_DAT_17[7]\, \ELK_RX_SER_WORD_17[0]\, 
        \ELK_RX_SER_WORD_17[1]\, \ELK_RX_SER_WORD_17[2]\, 
        \ELK_RX_SER_WORD_17[3]\, \ELK_RX_SER_WORD_17[4]\, 
        \ELK_RX_SER_WORD_17[5]\, \ELK_RX_SER_WORD_17[6]\, 
        \ELK_RX_SER_WORD_17[7]\, \PATT_ELK_DAT_18[0]\, 
        \PATT_ELK_DAT_18[1]\, \PATT_ELK_DAT_18[2]\, 
        \PATT_ELK_DAT_18[3]\, \PATT_ELK_DAT_18[4]\, 
        \PATT_ELK_DAT_18[5]\, \PATT_ELK_DAT_18[6]\, 
        \PATT_ELK_DAT_18[7]\, \ELK_RX_SER_WORD_18[0]\, 
        \ELK_RX_SER_WORD_18[1]\, \ELK_RX_SER_WORD_18[2]\, 
        \ELK_RX_SER_WORD_18[3]\, \ELK_RX_SER_WORD_18[4]\, 
        \ELK_RX_SER_WORD_18[5]\, \ELK_RX_SER_WORD_18[6]\, 
        \ELK_RX_SER_WORD_18[7]\, \PATT_ELK_DAT_19[0]\, 
        \PATT_ELK_DAT_19[1]\, \PATT_ELK_DAT_19[2]\, 
        \PATT_ELK_DAT_19[3]\, \PATT_ELK_DAT_19[4]\, 
        \PATT_ELK_DAT_19[5]\, \PATT_ELK_DAT_19[6]\, 
        \PATT_ELK_DAT_19[7]\, \ELK_RX_SER_WORD_19[0]\, 
        \ELK_RX_SER_WORD_19[1]\, \ELK_RX_SER_WORD_19[2]\, 
        \ELK_RX_SER_WORD_19[3]\, \ELK_RX_SER_WORD_19[4]\, 
        \ELK_RX_SER_WORD_19[5]\, \ELK_RX_SER_WORD_19[6]\, 
        \ELK_RX_SER_WORD_19[7]\, USB_OE_BI, USB_RD_BI, USB_WR_BI, 
        USB_SIWU_BI, \TFC_ADDRB[0]\, \TFC_ADDRB[1]\, 
        \TFC_ADDRB[2]\, \TFC_ADDRB[3]\, \TFC_ADDRB[4]\, 
        \TFC_ADDRB[5]\, \TFC_ADDRB[6]\, \TFC_ADDRB[7]\, 
        TFC_RAM_BLKB_EN, TFC_RWB, \ELKS_ADDRB[0]\, 
        \ELKS_ADDRB[1]\, \ELKS_ADDRB[2]\, \ELKS_ADDRB[3]\, 
        \ELKS_ADDRB[4]\, \ELKS_ADDRB[5]\, \ELKS_ADDRB[6]\, 
        \ELKS_ADDRB[7]\, ELKS_RAM_BLKB_EN, ELKS_RWB, DEV_RST_B_c, 
        DCB_SALT_SEL_c, EXTCLK_40MHZ_c, EXT_INT_REF_SEL_c, 
        ALL_PLL_LOCK_c, P_MASTER_POR_B_c, P_USB_MASTER_EN_c, 
        CLK_40M_GL, CCC_160M_FXD, CCC_160M_ADJ, P_ELK0_SYNC_DET_c, 
        P_TFC_SYNC_DET_c, \OP_MODE_c[1]\, \OP_MODE_c[2]\, 
        \OP_MODE_c[5]\, \OP_MODE_c[6]\, USBCLK60MHZ_c, 
        ELK0_OUT_R_i_0, ELK0_OUT_F_i_0, MASTER_DCB_POR_B_i_0_i, 
        P_USB_MASTER_EN_c_0, P_USB_MASTER_EN_c_22, 
        \ELKS_ADDRB_0[6]\, \ELKS_ADDRB_0[4]\, \ELKS_ADDRB_0[2]\, 
        P_USB_MASTER_EN_c_22_0, \U_ELK1_CH/ELK_IN_F_net_1\, 
        \U_ELK1_CH/ELK_IN_R_net_1\, \U_ELK1_CH/ELK_OUT_F_i_0\, 
        \U_ELK1_CH/ELK_OUT_R_i_0\, 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[0]_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[1]_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[2]_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[3]_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[11]_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[12]_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[13]_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[14]_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[0]\, 
        \U_ELK1_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[1]\, 
        \U_ELK1_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[2]\, 
        \U_ELK1_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[3]\, 
        \U_ELK1_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[4]\, 
        \U_ELK1_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[5]\, 
        \U_ELK1_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[6]\, 
        \U_ELK1_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[7]\, 
        \U_ELK1_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/Q[0]_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/Q[1]_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/Q[2]_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/Q[3]_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/Q[4]_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/Q[5]_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/Q[6]_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/Q[7]_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/Q[8]_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/Q[9]_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/Q[10]_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/Q[11]_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/Q[12]_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/Q[13]_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[13]_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/Q[14]_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[14]_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]_net_1\, 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]_net_1\, 
        \U_ELK1_CH/U_DDR_ELK1/ELK_IN_DDR_R\, 
        \U_ELK1_CH/U_DDR_ELK1/ELK_IN_DDR_F\, \GND\, 
        \U_ELK3_CH/ELK_IN_F_net_1\, \U_ELK3_CH/ELK_IN_R_net_1\, 
        \U_ELK3_CH/ELK_OUT_F_i_0\, \U_ELK3_CH/ELK_OUT_R_i_0\, 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[0]_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[1]_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[2]_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[3]_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[11]_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[12]_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[13]_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[14]_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[0]\, 
        \U_ELK3_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[1]\, 
        \U_ELK3_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[2]\, 
        \U_ELK3_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[3]\, 
        \U_ELK3_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[4]\, 
        \U_ELK3_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[5]\, 
        \U_ELK3_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[6]\, 
        \U_ELK3_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[7]\, 
        \U_ELK3_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/Q[0]_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/Q[1]_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/Q[2]_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/Q[3]_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/Q[4]_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/Q[5]_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/Q[6]_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/Q[7]_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/Q[8]_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/Q[9]_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/Q[10]_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/Q[11]_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/Q[12]_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/Q[13]_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[13]_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/Q[14]_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[14]_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]_net_1\, 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]_net_1\, 
        \U_ELK3_CH/U_DDR_ELK1/ELK_IN_DDR_R\, 
        \U_ELK3_CH/U_DDR_ELK1/ELK_IN_DDR_F\, 
        \U50_PATTERNS/RD_USB_ADBUS[6]\, 
        \U50_PATTERNS/RD_USB_ADBUS[7]\, 
        \U50_PATTERNS/ELINK_DOUTA_6[1]\, 
        \U50_PATTERNS/ELINK_DOUTA_16[1]\, 
        \U50_PATTERNS/ELINK_DOUTA_5[6]\, 
        \U50_PATTERNS/ELINK_DOUTA_16[7]\, 
        \U50_PATTERNS/ELINK_DOUTA_5[3]\, 
        \U50_PATTERNS/ELINK_DOUTA_0[3]\, 
        \U50_PATTERNS/ELINK_DOUTA_16[0]\, 
        \U50_PATTERNS/ELINK_DOUTA_5[5]\, 
        \U50_PATTERNS/ELINK_DOUTA_0[5]\, 
        \U50_PATTERNS/ELINK_DOUTA_6[3]\, 
        \U50_PATTERNS/ELINK_DOUTA_5[1]\, 
        \U50_PATTERNS/ELINK_DOUTA_0[1]\, 
        \U50_PATTERNS/ELINK_DOUTA_3[0]\, 
        \U50_PATTERNS/ELINK_DOUTA_11[7]\, 
        \U50_PATTERNS/ELINK_DOUTA_16[3]\, 
        \U50_PATTERNS/ELINK_DOUTA_6[6]\, 
        \U50_PATTERNS/ELINK_DOUTA_6[5]\, 
        \U50_PATTERNS/ELINK_DOUTA_16[5]\, \U50_PATTERNS/TrienAux\, 
        \U50_PATTERNS/ELINK_DOUTA_13[1]\, 
        \U50_PATTERNS/ELINK_DOUTA_8[1]\, 
        \U50_PATTERNS/ELINK_DOUTA_10[1]\, 
        \U50_PATTERNS/ELINK_DOUTA_2[1]\, 
        \U50_PATTERNS/ELINK_DOUTA_1[1]\, 
        \U50_PATTERNS/ELINK_DOUTA_0[6]\, 
        \U50_PATTERNS/ELINK_DOUTA_2[6]\, 
        \U50_PATTERNS/ELINK_DOUTA_11[6]\, 
        \U50_PATTERNS/ELINK_DOUTA_10[6]\, 
        \U50_PATTERNS/ELINK_DOUTA_17[6]\, 
        \U50_PATTERNS/ELINK_DOUTA_16[6]\, 
        \U50_PATTERNS/ELINK_DOUTA_3[7]\, 
        \U50_PATTERNS/ELINK_DOUTA_1[7]\, 
        \U50_PATTERNS/ELINK_DOUTA_0[7]\, 
        \U50_PATTERNS/ELINK_DOUTA_17[7]\, 
        \U50_PATTERNS/ELINK_DOUTA_6[7]\, 
        \U50_PATTERNS/ELINK_DOUTA_5[7]\, 
        \U50_PATTERNS/ELINK_DOUTA_6[4]\, 
        \U50_PATTERNS/ELINK_DOUTA_2[4]\, 
        \U50_PATTERNS/ELINK_DOUTA_0[4]\, 
        \U50_PATTERNS/ELINK_DOUTA_8[4]\, 
        \U50_PATTERNS/ELINK_DOUTA_11[4]\, 
        \U50_PATTERNS/ELINK_DOUTA_13[4]\, 
        \U50_PATTERNS/ELINK_DOUTA_16[4]\, 
        \U50_PATTERNS/ELINK_DOUTA_13[3]\, 
        \U50_PATTERNS/ELINK_DOUTA_10[3]\, 
        \U50_PATTERNS/ELINK_DOUTA_8[3]\, 
        \U50_PATTERNS/ELINK_DOUTA_2[3]\, 
        \U50_PATTERNS/ELINK_DOUTA_1[3]\, 
        \U50_PATTERNS/ELINK_DOUTA_1[0]\, 
        \U50_PATTERNS/ELINK_DOUTA_17[0]\, 
        \U50_PATTERNS/ELINK_DOUTA_13[0]\, 
        \U50_PATTERNS/ELINK_DOUTA_10[0]\, 
        \U50_PATTERNS/ELINK_DOUTA_8[0]\, 
        \U50_PATTERNS/ELINK_DOUTA_6[0]\, 
        \U50_PATTERNS/ELINK_DOUTA_13[2]\, 
        \U50_PATTERNS/ELINK_DOUTA_17[2]\, 
        \U50_PATTERNS/ELINK_DOUTA_1[2]\, 
        \U50_PATTERNS/ELINK_DOUTA_2[2]\, 
        \U50_PATTERNS/ELINK_DOUTA_5[2]\, 
        \U50_PATTERNS/ELINK_DOUTA_6[2]\, 
        \U50_PATTERNS/ELINK_DOUTA_8[2]\, 
        \U50_PATTERNS/ELINK_DOUTA_13[5]\, 
        \U50_PATTERNS/ELINK_DOUTA_10[5]\, 
        \U50_PATTERNS/ELINK_DOUTA_8[5]\, 
        \U50_PATTERNS/ELINK_DOUTA_2[5]\, 
        \U50_PATTERNS/ELINK_DOUTA_1[5]\, 
        \U50_PATTERNS/RD_USB_ADBUS[4]\, \U50_PATTERNS/USB_RXF_B\, 
        \U50_PATTERNS/RD_USB_ADBUS[2]\, 
        \U50_PATTERNS/RD_USB_ADBUS[3]\, \U50_PATTERNS/USB_TXE_B\, 
        \U50_PATTERNS/RD_USB_ADBUS[5]\, 
        \U50_PATTERNS/RD_USB_ADBUS[1]\, 
        \U50_PATTERNS/RD_USB_ADBUS[0]\, 
        \U50_PATTERNS/ELINK_RWA[19]\, 
        \U50_PATTERNS/ELINK_RWA[18]\, 
        \U50_PATTERNS/ELINK_RWA[16]\, \U50_PATTERNS/ELINK_RWA[9]\, 
        \U50_PATTERNS/ELINK_RWA[15]\, 
        \U50_PATTERNS/ELINK_RWA[14]\, 
        \U50_PATTERNS/ELINK_RWA[12]\, 
        \U50_PATTERNS/ELINK_RWA[10]\, \U50_PATTERNS/ELINK_RWA[8]\, 
        \U50_PATTERNS/ELINK_RWA[7]\, \U50_PATTERNS/ELINK_RWA[5]\, 
        \U50_PATTERNS/ELINK_RWA[4]\, \U50_PATTERNS/ELINK_RWA[1]\, 
        \U50_PATTERNS/ELINK_RWA[11]\, \U50_PATTERNS/ELINK_RWA[3]\, 
        \U50_PATTERNS/ELINK_RWA[17]\, 
        \U50_PATTERNS/ELINK_BLKA[17]\, 
        \U50_PATTERNS/ELINK_RWA[13]\, \U50_PATTERNS/ELINK_RWA[6]\, 
        \U50_PATTERNS/ELINK_RWA[2]\, 
        \U50_PATTERNS/ELINK_DOUTA_18[0]\, 
        \U50_PATTERNS/ELINK_DOUTA_9[0]\, 
        \U50_PATTERNS/ELINK_DOUTA_15[0]\, 
        \U50_PATTERNS/ELINK_DOUTA_14[0]\, 
        \U50_PATTERNS/ELINK_DOUTA_12[0]\, 
        \U50_PATTERNS/ELINK_DOUTA_11[0]\, 
        \U50_PATTERNS/ELINK_DOUTA_19[3]\, 
        \U50_PATTERNS/ELINK_DOUTA_14[3]\, 
        \U50_PATTERNS/ELINK_DOUTA_12[3]\, 
        \U50_PATTERNS/ELINK_DOUTA_11[3]\, 
        \U50_PATTERNS/ELINK_DOUTA_9[3]\, 
        \U50_PATTERNS/ELINK_DOUTA_7[3]\, 
        \U50_PATTERNS/ELINK_DOUTA_4[3]\, 
        \U50_PATTERNS/ELINK_DOUTA_3[3]\, 
        \U50_PATTERNS/TFC_DOUTA[3]\, 
        \U50_PATTERNS/ELINK_DOUTA_19[1]\, 
        \U50_PATTERNS/ELINK_DOUTA_4[1]\, 
        \U50_PATTERNS/ELINK_DOUTA_3[1]\, 
        \U50_PATTERNS/TFC_DOUTA[1]\, 
        \U50_PATTERNS/ELINK_DOUTA_19[0]\, 
        \U50_PATTERNS/ELINK_DOUTA_7[0]\, 
        \U50_PATTERNS/ELINK_DOUTA_5[0]\, 
        \U50_PATTERNS/ELINK_DOUTA_4[0]\, 
        \U50_PATTERNS/ELINK_DOUTA_2[0]\, 
        \U50_PATTERNS/ELINK_DOUTA_0[0]\, 
        \U50_PATTERNS/TFC_DOUTA[0]\, 
        \U50_PATTERNS/ELINK_DOUTA_18[2]\, 
        \U50_PATTERNS/ELINK_DOUTA_16[2]\, 
        \U50_PATTERNS/ELINK_DOUTA_15[2]\, 
        \U50_PATTERNS/ELINK_DOUTA_17[4]\, 
        \U50_PATTERNS/ELINK_DOUTA_15[4]\, 
        \U50_PATTERNS/ELINK_DOUTA_10[4]\, 
        \U50_PATTERNS/ELINK_DOUTA_9[4]\, 
        \U50_PATTERNS/ELINK_DOUTA_7[4]\, 
        \U50_PATTERNS/ELINK_DOUTA_5[4]\, 
        \U50_PATTERNS/ELINK_DOUTA_4[4]\, 
        \U50_PATTERNS/ELINK_DOUTA_3[4]\, 
        \U50_PATTERNS/ELINK_DOUTA_1[4]\, 
        \U50_PATTERNS/TFC_DOUTA[4]\, \U50_PATTERNS/ELINK_RWA[0]\, 
        \U50_PATTERNS/ELINK_DOUTA_18[7]\, 
        \U50_PATTERNS/ELINK_DOUTA_15[7]\, 
        \U50_PATTERNS/ELINK_DOUTA_14[7]\, 
        \U50_PATTERNS/ELINK_DOUTA_13[7]\, 
        \U50_PATTERNS/ELINK_DOUTA_12[7]\, 
        \U50_PATTERNS/ELINK_DOUTA_10[7]\, 
        \U50_PATTERNS/ELINK_DOUTA_9[7]\, 
        \U50_PATTERNS/ELINK_DOUTA_8[7]\, 
        \U50_PATTERNS/ELINK_DOUTA_7[7]\, 
        \U50_PATTERNS/ELINK_DOUTA_4[7]\, 
        \U50_PATTERNS/ELINK_DOUTA_2[7]\, 
        \U50_PATTERNS/TFC_DOUTA[7]\, 
        \U50_PATTERNS/ELINK_DOUTA_18[3]\, 
        \U50_PATTERNS/ELINK_DOUTA_17[3]\, 
        \U50_PATTERNS/ELINK_DOUTA_15[3]\, 
        \U50_PATTERNS/ELINK_DOUTA_18[1]\, 
        \U50_PATTERNS/ELINK_DOUTA_17[1]\, 
        \U50_PATTERNS/ELINK_DOUTA_15[1]\, 
        \U50_PATTERNS/TFC_DOUTA[6]\, 
        \U50_PATTERNS/ELINK_DOUTA_1[6]\, 
        \U50_PATTERNS/ELINK_DOUTA_3[6]\, 
        \U50_PATTERNS/ELINK_DOUTA_4[6]\, 
        \U50_PATTERNS/ELINK_DOUTA_7[6]\, 
        \U50_PATTERNS/ELINK_DOUTA_8[6]\, 
        \U50_PATTERNS/ELINK_DOUTA_9[6]\, 
        \U50_PATTERNS/ELINK_DOUTA_12[6]\, 
        \U50_PATTERNS/ELINK_DOUTA_13[6]\, 
        \U50_PATTERNS/ELINK_DOUTA_14[6]\, 
        \U50_PATTERNS/ELINK_DOUTA_15[6]\, 
        \U50_PATTERNS/ELINK_DOUTA_18[6]\, 
        \U50_PATTERNS/ELINK_DOUTA_19[6]\, 
        \U50_PATTERNS/ELINK_DOUTA_7[1]\, 
        \U50_PATTERNS/ELINK_DOUTA_9[1]\, 
        \U50_PATTERNS/ELINK_DOUTA_11[1]\, 
        \U50_PATTERNS/ELINK_DOUTA_12[1]\, 
        \U50_PATTERNS/ELINK_DOUTA_14[1]\, 
        \U50_PATTERNS/TFC_DOUTA[5]\, 
        \U50_PATTERNS/ELINK_DOUTA_3[5]\, 
        \U50_PATTERNS/ELINK_DOUTA_4[5]\, 
        \U50_PATTERNS/ELINK_DOUTA_7[5]\, 
        \U50_PATTERNS/ELINK_DOUTA_9[5]\, 
        \U50_PATTERNS/ELINK_DOUTA_11[5]\, 
        \U50_PATTERNS/ELINK_DOUTA_12[5]\, 
        \U50_PATTERNS/ELINK_DOUTA_14[5]\, 
        \U50_PATTERNS/ELINK_DOUTA_15[5]\, 
        \U50_PATTERNS/ELINK_DOUTA_17[5]\, 
        \U50_PATTERNS/ELINK_DOUTA_18[5]\, 
        \U50_PATTERNS/ELINK_DOUTA_19[5]\, 
        \U50_PATTERNS/ELINK_BLKA[13]\, 
        \U50_PATTERNS/ELINK_BLKA[19]\, 
        \U50_PATTERNS/ELINK_BLKA[16]\, 
        \U50_PATTERNS/ELINK_BLKA[11]\, 
        \U50_PATTERNS/ELINK_BLKA[9]\, 
        \U50_PATTERNS/ELINK_BLKA[12]\, 
        \U50_PATTERNS/ELINK_BLKA[10]\, 
        \U50_PATTERNS/ELINK_BLKA[8]\, 
        \U50_PATTERNS/ELINK_BLKA[7]\, 
        \U50_PATTERNS/ELINK_BLKA[5]\, 
        \U50_PATTERNS/ELINK_BLKA[4]\, 
        \U50_PATTERNS/ELINK_BLKA[3]\, 
        \U50_PATTERNS/ELINK_BLKA[1]\, 
        \U50_PATTERNS/ELINK_BLKA[18]\, 
        \U50_PATTERNS/ELINK_BLKA[14]\, 
        \U50_PATTERNS/ELINK_BLKA[15]\, 
        \U50_PATTERNS/ELINK_BLKA[6]\, 
        \U50_PATTERNS/ELINK_BLKA[0]\, 
        \U50_PATTERNS/ELINK_BLKA[2]\, 
        \U50_PATTERNS/ELINK_DOUTA_19[7]\, 
        \U50_PATTERNS/ELINK_DOUTA_12[4]\, 
        \U50_PATTERNS/ELINK_DOUTA_14[4]\, 
        \U50_PATTERNS/ELINK_DOUTA_18[4]\, 
        \U50_PATTERNS/ELINK_DOUTA_19[4]\, 
        \U50_PATTERNS/TFC_DOUTA[2]\, 
        \U50_PATTERNS/ELINK_DOUTA_0[2]\, 
        \U50_PATTERNS/ELINK_DOUTA_3[2]\, 
        \U50_PATTERNS/ELINK_DOUTA_4[2]\, 
        \U50_PATTERNS/ELINK_DOUTA_7[2]\, 
        \U50_PATTERNS/ELINK_DOUTA_9[2]\, 
        \U50_PATTERNS/ELINK_DOUTA_10[2]\, 
        \U50_PATTERNS/ELINK_DOUTA_11[2]\, 
        \U50_PATTERNS/ELINK_DOUTA_12[2]\, 
        \U50_PATTERNS/ELINK_DOUTA_14[2]\, 
        \U50_PATTERNS/ELINK_DOUTA_19[2]\, \U50_PATTERNS/TFC_BLKA\, 
        \U50_PATTERNS/TFC_RWA\, \U50_PATTERNS/ELINK_DINA_8[0]\, 
        \U50_PATTERNS/ELINK_DINA_8[1]\, 
        \U50_PATTERNS/ELINK_DINA_8[2]\, 
        \U50_PATTERNS/ELINK_DINA_8[3]\, 
        \U50_PATTERNS/ELINK_DINA_8[4]\, 
        \U50_PATTERNS/ELINK_DINA_8[5]\, 
        \U50_PATTERNS/ELINK_DINA_8[6]\, 
        \U50_PATTERNS/ELINK_DINA_8[7]\, 
        \U50_PATTERNS/ELINK_DINA_7[0]\, 
        \U50_PATTERNS/ELINK_DINA_7[1]\, 
        \U50_PATTERNS/ELINK_DINA_7[2]\, 
        \U50_PATTERNS/ELINK_DINA_7[3]\, 
        \U50_PATTERNS/ELINK_DINA_7[4]\, 
        \U50_PATTERNS/ELINK_DINA_7[5]\, 
        \U50_PATTERNS/ELINK_DINA_7[6]\, 
        \U50_PATTERNS/ELINK_DINA_7[7]\, 
        \U50_PATTERNS/ELINK_DINA_6[0]\, 
        \U50_PATTERNS/ELINK_DINA_6[1]\, 
        \U50_PATTERNS/ELINK_DINA_6[2]\, 
        \U50_PATTERNS/ELINK_DINA_6[3]\, 
        \U50_PATTERNS/ELINK_DINA_6[4]\, 
        \U50_PATTERNS/ELINK_DINA_6[5]\, 
        \U50_PATTERNS/ELINK_DINA_6[6]\, 
        \U50_PATTERNS/ELINK_DINA_6[7]\, 
        \U50_PATTERNS/ELINK_DINA_5[0]\, 
        \U50_PATTERNS/ELINK_DINA_5[1]\, 
        \U50_PATTERNS/ELINK_DINA_5[2]\, 
        \U50_PATTERNS/ELINK_DINA_5[3]\, 
        \U50_PATTERNS/ELINK_DINA_5[4]\, 
        \U50_PATTERNS/ELINK_DINA_5[5]\, 
        \U50_PATTERNS/ELINK_DINA_5[6]\, 
        \U50_PATTERNS/ELINK_DINA_5[7]\, 
        \U50_PATTERNS/ELINK_DINA_4[0]\, 
        \U50_PATTERNS/ELINK_DINA_4[1]\, 
        \U50_PATTERNS/ELINK_DINA_4[2]\, 
        \U50_PATTERNS/ELINK_DINA_4[3]\, 
        \U50_PATTERNS/ELINK_DINA_4[4]\, 
        \U50_PATTERNS/ELINK_DINA_4[5]\, 
        \U50_PATTERNS/ELINK_DINA_4[6]\, 
        \U50_PATTERNS/ELINK_DINA_4[7]\, 
        \U50_PATTERNS/ELINK_DINA_3[0]\, 
        \U50_PATTERNS/ELINK_DINA_3[1]\, 
        \U50_PATTERNS/ELINK_DINA_3[2]\, 
        \U50_PATTERNS/ELINK_DINA_3[3]\, 
        \U50_PATTERNS/ELINK_DINA_3[4]\, 
        \U50_PATTERNS/ELINK_DINA_3[5]\, 
        \U50_PATTERNS/ELINK_DINA_3[6]\, 
        \U50_PATTERNS/ELINK_DINA_3[7]\, 
        \U50_PATTERNS/ELINK_DINA_2[0]\, 
        \U50_PATTERNS/ELINK_DINA_2[1]\, 
        \U50_PATTERNS/ELINK_DINA_2[2]\, 
        \U50_PATTERNS/ELINK_DINA_2[3]\, 
        \U50_PATTERNS/ELINK_DINA_2[4]\, 
        \U50_PATTERNS/ELINK_DINA_2[5]\, 
        \U50_PATTERNS/ELINK_DINA_2[6]\, 
        \U50_PATTERNS/ELINK_DINA_2[7]\, 
        \U50_PATTERNS/ELINK_DINA_1[0]\, 
        \U50_PATTERNS/ELINK_DINA_1[1]\, 
        \U50_PATTERNS/ELINK_DINA_1[2]\, 
        \U50_PATTERNS/ELINK_DINA_1[3]\, 
        \U50_PATTERNS/ELINK_DINA_1[4]\, 
        \U50_PATTERNS/ELINK_DINA_1[5]\, 
        \U50_PATTERNS/ELINK_DINA_1[6]\, 
        \U50_PATTERNS/ELINK_DINA_1[7]\, 
        \U50_PATTERNS/ELINK_DINA_0[0]\, 
        \U50_PATTERNS/ELINK_DINA_0[1]\, 
        \U50_PATTERNS/ELINK_DINA_0[2]\, 
        \U50_PATTERNS/ELINK_DINA_0[3]\, 
        \U50_PATTERNS/ELINK_DINA_0[4]\, 
        \U50_PATTERNS/ELINK_DINA_0[5]\, 
        \U50_PATTERNS/ELINK_DINA_0[6]\, 
        \U50_PATTERNS/ELINK_DINA_0[7]\, 
        \U50_PATTERNS/WR_USB_ADBUS[0]\, 
        \U50_PATTERNS/WR_USB_ADBUS[1]\, 
        \U50_PATTERNS/WR_USB_ADBUS[2]\, 
        \U50_PATTERNS/WR_USB_ADBUS[3]\, 
        \U50_PATTERNS/WR_USB_ADBUS[4]\, 
        \U50_PATTERNS/WR_USB_ADBUS[5]\, 
        \U50_PATTERNS/WR_USB_ADBUS[6]\, 
        \U50_PATTERNS/WR_USB_ADBUS[7]\, 
        \U50_PATTERNS/ELINK_ADDRA_1[0]\, 
        \U50_PATTERNS/ELINK_ADDRA_1[1]\, 
        \U50_PATTERNS/ELINK_ADDRA_1[2]\, 
        \U50_PATTERNS/ELINK_ADDRA_1[3]\, 
        \U50_PATTERNS/ELINK_ADDRA_1[4]\, 
        \U50_PATTERNS/ELINK_ADDRA_1[5]\, 
        \U50_PATTERNS/ELINK_ADDRA_1[6]\, 
        \U50_PATTERNS/ELINK_ADDRA_1[7]\, 
        \U50_PATTERNS/ELINK_ADDRA_0[0]\, 
        \U50_PATTERNS/ELINK_ADDRA_0[1]\, 
        \U50_PATTERNS/ELINK_ADDRA_0[2]\, 
        \U50_PATTERNS/ELINK_ADDRA_0[3]\, 
        \U50_PATTERNS/ELINK_ADDRA_0[4]\, 
        \U50_PATTERNS/ELINK_ADDRA_0[5]\, 
        \U50_PATTERNS/ELINK_ADDRA_0[6]\, 
        \U50_PATTERNS/ELINK_ADDRA_0[7]\, 
        \U50_PATTERNS/TFC_DINA[0]\, \U50_PATTERNS/TFC_DINA[1]\, 
        \U50_PATTERNS/TFC_DINA[2]\, \U50_PATTERNS/TFC_DINA[3]\, 
        \U50_PATTERNS/TFC_DINA[4]\, \U50_PATTERNS/TFC_DINA[5]\, 
        \U50_PATTERNS/TFC_DINA[6]\, \U50_PATTERNS/TFC_DINA[7]\, 
        \U50_PATTERNS/ELINK_DINA_19[0]\, 
        \U50_PATTERNS/ELINK_DINA_19[1]\, 
        \U50_PATTERNS/ELINK_DINA_19[2]\, 
        \U50_PATTERNS/ELINK_DINA_19[3]\, 
        \U50_PATTERNS/ELINK_DINA_19[4]\, 
        \U50_PATTERNS/ELINK_DINA_19[5]\, 
        \U50_PATTERNS/ELINK_DINA_19[6]\, 
        \U50_PATTERNS/ELINK_DINA_19[7]\, 
        \U50_PATTERNS/ELINK_DINA_18[0]\, 
        \U50_PATTERNS/ELINK_DINA_18[1]\, 
        \U50_PATTERNS/ELINK_DINA_18[2]\, 
        \U50_PATTERNS/ELINK_DINA_18[3]\, 
        \U50_PATTERNS/ELINK_DINA_18[4]\, 
        \U50_PATTERNS/ELINK_DINA_18[5]\, 
        \U50_PATTERNS/ELINK_DINA_18[6]\, 
        \U50_PATTERNS/ELINK_DINA_18[7]\, 
        \U50_PATTERNS/ELINK_DINA_17[0]\, 
        \U50_PATTERNS/ELINK_DINA_17[1]\, 
        \U50_PATTERNS/ELINK_DINA_17[2]\, 
        \U50_PATTERNS/ELINK_DINA_17[3]\, 
        \U50_PATTERNS/ELINK_DINA_17[4]\, 
        \U50_PATTERNS/ELINK_DINA_17[5]\, 
        \U50_PATTERNS/ELINK_DINA_17[6]\, 
        \U50_PATTERNS/ELINK_DINA_17[7]\, 
        \U50_PATTERNS/ELINK_DINA_16[0]\, 
        \U50_PATTERNS/ELINK_DINA_16[1]\, 
        \U50_PATTERNS/ELINK_DINA_16[2]\, 
        \U50_PATTERNS/ELINK_DINA_16[3]\, 
        \U50_PATTERNS/ELINK_DINA_16[4]\, 
        \U50_PATTERNS/ELINK_DINA_16[5]\, 
        \U50_PATTERNS/ELINK_DINA_16[6]\, 
        \U50_PATTERNS/ELINK_DINA_16[7]\, 
        \U50_PATTERNS/ELINK_DINA_15[0]\, 
        \U50_PATTERNS/ELINK_DINA_15[1]\, 
        \U50_PATTERNS/ELINK_DINA_15[2]\, 
        \U50_PATTERNS/ELINK_DINA_15[3]\, 
        \U50_PATTERNS/ELINK_DINA_15[4]\, 
        \U50_PATTERNS/ELINK_DINA_15[5]\, 
        \U50_PATTERNS/ELINK_DINA_15[6]\, 
        \U50_PATTERNS/ELINK_DINA_15[7]\, 
        \U50_PATTERNS/ELINK_DINA_14[0]\, 
        \U50_PATTERNS/ELINK_DINA_14[1]\, 
        \U50_PATTERNS/ELINK_DINA_14[2]\, 
        \U50_PATTERNS/ELINK_DINA_14[3]\, 
        \U50_PATTERNS/ELINK_DINA_14[4]\, 
        \U50_PATTERNS/ELINK_DINA_14[5]\, 
        \U50_PATTERNS/ELINK_DINA_14[6]\, 
        \U50_PATTERNS/ELINK_DINA_14[7]\, 
        \U50_PATTERNS/ELINK_DINA_13[0]\, 
        \U50_PATTERNS/ELINK_DINA_13[1]\, 
        \U50_PATTERNS/ELINK_DINA_13[2]\, 
        \U50_PATTERNS/ELINK_DINA_13[3]\, 
        \U50_PATTERNS/ELINK_DINA_13[4]\, 
        \U50_PATTERNS/ELINK_DINA_13[5]\, 
        \U50_PATTERNS/ELINK_DINA_13[6]\, 
        \U50_PATTERNS/ELINK_DINA_13[7]\, 
        \U50_PATTERNS/ELINK_DINA_12[0]\, 
        \U50_PATTERNS/ELINK_DINA_12[1]\, 
        \U50_PATTERNS/ELINK_DINA_12[2]\, 
        \U50_PATTERNS/ELINK_DINA_12[3]\, 
        \U50_PATTERNS/ELINK_DINA_12[4]\, 
        \U50_PATTERNS/ELINK_DINA_12[5]\, 
        \U50_PATTERNS/ELINK_DINA_12[6]\, 
        \U50_PATTERNS/ELINK_DINA_12[7]\, 
        \U50_PATTERNS/ELINK_DINA_11[0]\, 
        \U50_PATTERNS/ELINK_DINA_11[1]\, 
        \U50_PATTERNS/ELINK_DINA_11[2]\, 
        \U50_PATTERNS/ELINK_DINA_11[3]\, 
        \U50_PATTERNS/ELINK_DINA_11[4]\, 
        \U50_PATTERNS/ELINK_DINA_11[5]\, 
        \U50_PATTERNS/ELINK_DINA_11[6]\, 
        \U50_PATTERNS/ELINK_DINA_11[7]\, 
        \U50_PATTERNS/ELINK_DINA_10[0]\, 
        \U50_PATTERNS/ELINK_DINA_10[1]\, 
        \U50_PATTERNS/ELINK_DINA_10[2]\, 
        \U50_PATTERNS/ELINK_DINA_10[3]\, 
        \U50_PATTERNS/ELINK_DINA_10[4]\, 
        \U50_PATTERNS/ELINK_DINA_10[5]\, 
        \U50_PATTERNS/ELINK_DINA_10[6]\, 
        \U50_PATTERNS/ELINK_DINA_10[7]\, 
        \U50_PATTERNS/ELINK_DINA_9[0]\, 
        \U50_PATTERNS/ELINK_DINA_9[1]\, 
        \U50_PATTERNS/ELINK_DINA_9[2]\, 
        \U50_PATTERNS/ELINK_DINA_9[3]\, 
        \U50_PATTERNS/ELINK_DINA_9[4]\, 
        \U50_PATTERNS/ELINK_DINA_9[5]\, 
        \U50_PATTERNS/ELINK_DINA_9[6]\, 
        \U50_PATTERNS/ELINK_DINA_9[7]\, 
        \U50_PATTERNS/ELINK_ADDRA_16[0]\, 
        \U50_PATTERNS/ELINK_ADDRA_16[1]\, 
        \U50_PATTERNS/ELINK_ADDRA_16[2]\, 
        \U50_PATTERNS/ELINK_ADDRA_16[3]\, 
        \U50_PATTERNS/ELINK_ADDRA_16[4]\, 
        \U50_PATTERNS/ELINK_ADDRA_16[5]\, 
        \U50_PATTERNS/ELINK_ADDRA_16[6]\, 
        \U50_PATTERNS/ELINK_ADDRA_16[7]\, 
        \U50_PATTERNS/ELINK_ADDRA_15[0]\, 
        \U50_PATTERNS/ELINK_ADDRA_15[1]\, 
        \U50_PATTERNS/ELINK_ADDRA_15[2]\, 
        \U50_PATTERNS/ELINK_ADDRA_15[3]\, 
        \U50_PATTERNS/ELINK_ADDRA_15[4]\, 
        \U50_PATTERNS/ELINK_ADDRA_15[5]\, 
        \U50_PATTERNS/ELINK_ADDRA_15[6]\, 
        \U50_PATTERNS/ELINK_ADDRA_15[7]\, 
        \U50_PATTERNS/ELINK_ADDRA_14[0]\, 
        \U50_PATTERNS/ELINK_ADDRA_14[1]\, 
        \U50_PATTERNS/ELINK_ADDRA_14[2]\, 
        \U50_PATTERNS/ELINK_ADDRA_14[3]\, 
        \U50_PATTERNS/ELINK_ADDRA_14[4]\, 
        \U50_PATTERNS/ELINK_ADDRA_14[5]\, 
        \U50_PATTERNS/ELINK_ADDRA_14[6]\, 
        \U50_PATTERNS/ELINK_ADDRA_14[7]\, 
        \U50_PATTERNS/ELINK_ADDRA_13[0]\, 
        \U50_PATTERNS/ELINK_ADDRA_13[1]\, 
        \U50_PATTERNS/ELINK_ADDRA_13[2]\, 
        \U50_PATTERNS/ELINK_ADDRA_13[3]\, 
        \U50_PATTERNS/ELINK_ADDRA_13[4]\, 
        \U50_PATTERNS/ELINK_ADDRA_13[5]\, 
        \U50_PATTERNS/ELINK_ADDRA_13[6]\, 
        \U50_PATTERNS/ELINK_ADDRA_13[7]\, 
        \U50_PATTERNS/ELINK_ADDRA_12[0]\, 
        \U50_PATTERNS/ELINK_ADDRA_12[1]\, 
        \U50_PATTERNS/ELINK_ADDRA_12[2]\, 
        \U50_PATTERNS/ELINK_ADDRA_12[3]\, 
        \U50_PATTERNS/ELINK_ADDRA_12[4]\, 
        \U50_PATTERNS/ELINK_ADDRA_12[5]\, 
        \U50_PATTERNS/ELINK_ADDRA_12[6]\, 
        \U50_PATTERNS/ELINK_ADDRA_12[7]\, 
        \U50_PATTERNS/ELINK_ADDRA_11[0]\, 
        \U50_PATTERNS/ELINK_ADDRA_11[1]\, 
        \U50_PATTERNS/ELINK_ADDRA_11[2]\, 
        \U50_PATTERNS/ELINK_ADDRA_11[3]\, 
        \U50_PATTERNS/ELINK_ADDRA_11[4]\, 
        \U50_PATTERNS/ELINK_ADDRA_11[5]\, 
        \U50_PATTERNS/ELINK_ADDRA_11[6]\, 
        \U50_PATTERNS/ELINK_ADDRA_11[7]\, 
        \U50_PATTERNS/ELINK_ADDRA_10[0]\, 
        \U50_PATTERNS/ELINK_ADDRA_10[1]\, 
        \U50_PATTERNS/ELINK_ADDRA_10[2]\, 
        \U50_PATTERNS/ELINK_ADDRA_10[3]\, 
        \U50_PATTERNS/ELINK_ADDRA_10[4]\, 
        \U50_PATTERNS/ELINK_ADDRA_10[5]\, 
        \U50_PATTERNS/ELINK_ADDRA_10[6]\, 
        \U50_PATTERNS/ELINK_ADDRA_10[7]\, 
        \U50_PATTERNS/ELINK_ADDRA_9[0]\, 
        \U50_PATTERNS/ELINK_ADDRA_9[1]\, 
        \U50_PATTERNS/ELINK_ADDRA_9[2]\, 
        \U50_PATTERNS/ELINK_ADDRA_9[3]\, 
        \U50_PATTERNS/ELINK_ADDRA_9[4]\, 
        \U50_PATTERNS/ELINK_ADDRA_9[5]\, 
        \U50_PATTERNS/ELINK_ADDRA_9[6]\, 
        \U50_PATTERNS/ELINK_ADDRA_9[7]\, 
        \U50_PATTERNS/ELINK_ADDRA_8[0]\, 
        \U50_PATTERNS/ELINK_ADDRA_8[1]\, 
        \U50_PATTERNS/ELINK_ADDRA_8[2]\, 
        \U50_PATTERNS/ELINK_ADDRA_8[3]\, 
        \U50_PATTERNS/ELINK_ADDRA_8[4]\, 
        \U50_PATTERNS/ELINK_ADDRA_8[5]\, 
        \U50_PATTERNS/ELINK_ADDRA_8[6]\, 
        \U50_PATTERNS/ELINK_ADDRA_8[7]\, 
        \U50_PATTERNS/ELINK_ADDRA_7[0]\, 
        \U50_PATTERNS/ELINK_ADDRA_7[1]\, 
        \U50_PATTERNS/ELINK_ADDRA_7[2]\, 
        \U50_PATTERNS/ELINK_ADDRA_7[3]\, 
        \U50_PATTERNS/ELINK_ADDRA_7[4]\, 
        \U50_PATTERNS/ELINK_ADDRA_7[5]\, 
        \U50_PATTERNS/ELINK_ADDRA_7[6]\, 
        \U50_PATTERNS/ELINK_ADDRA_7[7]\, 
        \U50_PATTERNS/ELINK_ADDRA_6[0]\, 
        \U50_PATTERNS/ELINK_ADDRA_6[1]\, 
        \U50_PATTERNS/ELINK_ADDRA_6[2]\, 
        \U50_PATTERNS/ELINK_ADDRA_6[3]\, 
        \U50_PATTERNS/ELINK_ADDRA_6[4]\, 
        \U50_PATTERNS/ELINK_ADDRA_6[5]\, 
        \U50_PATTERNS/ELINK_ADDRA_6[6]\, 
        \U50_PATTERNS/ELINK_ADDRA_6[7]\, 
        \U50_PATTERNS/ELINK_ADDRA_5[0]\, 
        \U50_PATTERNS/ELINK_ADDRA_5[1]\, 
        \U50_PATTERNS/ELINK_ADDRA_5[2]\, 
        \U50_PATTERNS/ELINK_ADDRA_5[3]\, 
        \U50_PATTERNS/ELINK_ADDRA_5[4]\, 
        \U50_PATTERNS/ELINK_ADDRA_5[5]\, 
        \U50_PATTERNS/ELINK_ADDRA_5[6]\, 
        \U50_PATTERNS/ELINK_ADDRA_5[7]\, 
        \U50_PATTERNS/ELINK_ADDRA_4[0]\, 
        \U50_PATTERNS/ELINK_ADDRA_4[1]\, 
        \U50_PATTERNS/ELINK_ADDRA_4[2]\, 
        \U50_PATTERNS/ELINK_ADDRA_4[3]\, 
        \U50_PATTERNS/ELINK_ADDRA_4[4]\, 
        \U50_PATTERNS/ELINK_ADDRA_4[5]\, 
        \U50_PATTERNS/ELINK_ADDRA_4[6]\, 
        \U50_PATTERNS/ELINK_ADDRA_4[7]\, 
        \U50_PATTERNS/ELINK_ADDRA_3[0]\, 
        \U50_PATTERNS/ELINK_ADDRA_3[1]\, 
        \U50_PATTERNS/ELINK_ADDRA_3[2]\, 
        \U50_PATTERNS/ELINK_ADDRA_3[3]\, 
        \U50_PATTERNS/ELINK_ADDRA_3[4]\, 
        \U50_PATTERNS/ELINK_ADDRA_3[5]\, 
        \U50_PATTERNS/ELINK_ADDRA_3[6]\, 
        \U50_PATTERNS/ELINK_ADDRA_3[7]\, 
        \U50_PATTERNS/ELINK_ADDRA_2[0]\, 
        \U50_PATTERNS/ELINK_ADDRA_2[1]\, 
        \U50_PATTERNS/ELINK_ADDRA_2[2]\, 
        \U50_PATTERNS/ELINK_ADDRA_2[3]\, 
        \U50_PATTERNS/ELINK_ADDRA_2[4]\, 
        \U50_PATTERNS/ELINK_ADDRA_2[5]\, 
        \U50_PATTERNS/ELINK_ADDRA_2[6]\, 
        \U50_PATTERNS/ELINK_ADDRA_2[7]\, 
        \U50_PATTERNS/TFC_ADDRA[0]\, \U50_PATTERNS/TFC_ADDRA[1]\, 
        \U50_PATTERNS/TFC_ADDRA[2]\, \U50_PATTERNS/TFC_ADDRA[3]\, 
        \U50_PATTERNS/TFC_ADDRA[4]\, \U50_PATTERNS/TFC_ADDRA[5]\, 
        \U50_PATTERNS/TFC_ADDRA[6]\, \U50_PATTERNS/TFC_ADDRA[7]\, 
        \U50_PATTERNS/ELINK_ADDRA_19[0]\, 
        \U50_PATTERNS/ELINK_ADDRA_19[1]\, 
        \U50_PATTERNS/ELINK_ADDRA_19[2]\, 
        \U50_PATTERNS/ELINK_ADDRA_19[3]\, 
        \U50_PATTERNS/ELINK_ADDRA_19[4]\, 
        \U50_PATTERNS/ELINK_ADDRA_19[5]\, 
        \U50_PATTERNS/ELINK_ADDRA_19[6]\, 
        \U50_PATTERNS/ELINK_ADDRA_19[7]\, 
        \U50_PATTERNS/ELINK_ADDRA_18[0]\, 
        \U50_PATTERNS/ELINK_ADDRA_18[1]\, 
        \U50_PATTERNS/ELINK_ADDRA_18[2]\, 
        \U50_PATTERNS/ELINK_ADDRA_18[3]\, 
        \U50_PATTERNS/ELINK_ADDRA_18[4]\, 
        \U50_PATTERNS/ELINK_ADDRA_18[5]\, 
        \U50_PATTERNS/ELINK_ADDRA_18[6]\, 
        \U50_PATTERNS/ELINK_ADDRA_18[7]\, 
        \U50_PATTERNS/ELINK_ADDRA_17[0]\, 
        \U50_PATTERNS/ELINK_ADDRA_17[1]\, 
        \U50_PATTERNS/ELINK_ADDRA_17[2]\, 
        \U50_PATTERNS/ELINK_ADDRA_17[3]\, 
        \U50_PATTERNS/ELINK_ADDRA_17[4]\, 
        \U50_PATTERNS/ELINK_ADDRA_17[5]\, 
        \U50_PATTERNS/ELINK_ADDRA_17[6]\, 
        \U50_PATTERNS/ELINK_ADDRA_17[7]\, \VCC\, 
        \U_TFC_SERDAT_SOURCE/N_SERDAT[0]\, 
        \U_TFC_SERDAT_SOURCE/N_SERDAT[4]\, 
        \U_TFC_SERDAT_SOURCE/N_SERDAT[5]\, 
        \U_TFC_SERDAT_SOURCE/N_SERDAT[6]\, 
        \U_TFC_SERDAT_SOURCE/N_SERDAT[1]\, 
        \U_TFC_SERDAT_SOURCE/N_SERDAT[2]\, 
        \U_TFC_SERDAT_SOURCE/N_SERDAT[3]\, 
        \U_TFC_SERDAT_SOURCE/N_SERDAT[7]\, 
        \U_ELK18_CH/ELK_IN_F_net_1\, \U_ELK18_CH/ELK_IN_DDR_F\, 
        \U_ELK18_CH/ELK_IN_R_net_1\, \U_ELK18_CH/ELK_IN_DDR_R\, 
        \U_ELK18_CH/ELK_OUT_F\, \U_ELK18_CH/ELK_OUT_R\, 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[0]_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[1]_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[2]_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[3]_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[11]_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[12]_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[13]_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[14]_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[0]\, 
        \U_ELK18_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[1]\, 
        \U_ELK18_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[2]\, 
        \U_ELK18_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[3]\, 
        \U_ELK18_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[4]\, 
        \U_ELK18_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[5]\, 
        \U_ELK18_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[6]\, 
        \U_ELK18_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[7]\, 
        \U_ELK18_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/Q[0]_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/Q[1]_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/Q[2]_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/Q[3]_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/Q[4]_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/Q[5]_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/Q[6]_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/Q[7]_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/Q[8]_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/Q[9]_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/Q[10]_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/Q[11]_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/Q[12]_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/Q[13]_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[13]_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/Q[14]_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[14]_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]_net_1\, 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]_net_1\, 
        \U_ELK11_CH/ELK_IN_F_net_1\, \U_ELK11_CH/ELK_IN_DDR_F\, 
        \U_ELK11_CH/ELK_IN_R_net_1\, \U_ELK11_CH/ELK_IN_DDR_R\, 
        \U_ELK11_CH/ELK_OUT_F\, \U_ELK11_CH/ELK_OUT_R\, 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[0]_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[1]_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[2]_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[3]_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[11]_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[12]_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[13]_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[14]_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[0]\, 
        \U_ELK11_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[1]\, 
        \U_ELK11_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[2]\, 
        \U_ELK11_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[3]\, 
        \U_ELK11_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[4]\, 
        \U_ELK11_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[5]\, 
        \U_ELK11_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[6]\, 
        \U_ELK11_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[7]\, 
        \U_ELK11_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/Q[0]_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/Q[1]_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/Q[2]_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/Q[3]_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/Q[4]_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/Q[5]_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/Q[6]_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/Q[7]_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/Q[8]_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/Q[9]_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/Q[10]_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/Q[11]_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/Q[12]_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/Q[13]_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[13]_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/Q[14]_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[14]_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]_net_1\, 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]_net_1\, 
        \U_TFC_CMD_TX/N_SER_CMD_WORD_R[0]\, 
        \U_TFC_CMD_TX/START_RISE_net_1\, 
        \U_TFC_CMD_TX/N_SER_CMD_WORD_F[0]\, 
        \U_TFC_CMD_TX/N_SER_CMD_WORD_R[3]\, 
        \U_TFC_CMD_TX/SER_CMD_WORD_R[2]_net_1\, 
        \U_TFC_CMD_TX/N_SER_CMD_WORD_R[2]\, 
        \U_TFC_CMD_TX/SER_CMD_WORD_R[1]_net_1\, 
        \U_TFC_CMD_TX/N_SER_CMD_WORD_R[1]\, 
        \U_TFC_CMD_TX/SER_CMD_WORD_R[0]_net_1\, 
        \U_TFC_CMD_TX/N_SER_CMD_WORD_F[3]\, 
        \U_TFC_CMD_TX/SER_CMD_WORD_F[2]_net_1\, 
        \U_TFC_CMD_TX/N_SER_CMD_WORD_F[2]\, 
        \U_TFC_CMD_TX/SER_CMD_WORD_F[1]_net_1\, 
        \U_TFC_CMD_TX/N_SER_CMD_WORD_F[1]\, 
        \U_TFC_CMD_TX/SER_CMD_WORD_F[0]_net_1\, 
        \U_TFC_CMD_TX/N_START_RISE\, 
        \U_TFC_CMD_TX/CLK40M_GEN_DEL0_net_1\, 
        \U_TFC_CMD_TX/SER_OUT_FI_net_1\, 
        \U_TFC_CMD_TX/SER_OUT_RI_net_1\, 
        \U_TFC_CMD_TX/SER_CMD_WORD_F[3]_net_1\, 
        \U_TFC_CMD_TX/SER_CMD_WORD_R[3]_net_1\, 
        \U_ELK12_CH/ELK_IN_F_net_1\, \U_ELK12_CH/ELK_IN_DDR_F\, 
        \U_ELK12_CH/ELK_IN_R_net_1\, \U_ELK12_CH/ELK_IN_DDR_R\, 
        \U_ELK12_CH/ELK_OUT_F\, \U_ELK12_CH/ELK_OUT_R\, 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[0]_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[1]_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[2]_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[3]_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[11]_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[12]_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[13]_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[14]_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[0]\, 
        \U_ELK12_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[1]\, 
        \U_ELK12_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[2]\, 
        \U_ELK12_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[3]\, 
        \U_ELK12_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[4]\, 
        \U_ELK12_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[5]\, 
        \U_ELK12_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[6]\, 
        \U_ELK12_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[7]\, 
        \U_ELK12_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/Q[0]_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/Q[1]_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/Q[2]_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/Q[3]_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/Q[4]_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/Q[5]_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/Q[6]_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/Q[7]_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/Q[8]_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/Q[9]_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/Q[10]_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/Q[11]_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/Q[12]_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/Q[13]_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[13]_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/Q[14]_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[14]_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]_net_1\, 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]_net_1\, 
        \U_ELK13_CH/ELK_IN_F_net_1\, \U_ELK13_CH/ELK_IN_DDR_F\, 
        \U_ELK13_CH/ELK_IN_R_net_1\, \U_ELK13_CH/ELK_IN_DDR_R\, 
        \U_ELK13_CH/ELK_OUT_F\, \U_ELK13_CH/ELK_OUT_R\, 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[0]_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[1]_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[2]_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[3]_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[11]_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[12]_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[13]_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[14]_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[0]\, 
        \U_ELK13_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[1]\, 
        \U_ELK13_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[2]\, 
        \U_ELK13_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[3]\, 
        \U_ELK13_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[4]\, 
        \U_ELK13_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[5]\, 
        \U_ELK13_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[6]\, 
        \U_ELK13_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[7]\, 
        \U_ELK13_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/Q[0]_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/Q[1]_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/Q[2]_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/Q[3]_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/Q[4]_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/Q[5]_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/Q[6]_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/Q[7]_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/Q[8]_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/Q[9]_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/Q[10]_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/Q[11]_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/Q[12]_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/Q[13]_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[13]_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/Q[14]_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[14]_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]_net_1\, 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]_net_1\, 
        \U_EXEC_MASTER/MPOR_DCB_B_net_1\, 
        \U_ELK7_CH/ELK_IN_F_net_1\, \U_ELK7_CH/ELK_IN_DDR_F\, 
        \U_ELK7_CH/ELK_IN_R_net_1\, \U_ELK7_CH/ELK_IN_DDR_R\, 
        \U_ELK7_CH/ELK_OUT_F\, \U_ELK7_CH/ELK_OUT_R\, 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[0]_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[1]_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[2]_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[3]_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[11]_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[12]_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[13]_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[14]_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[0]\, 
        \U_ELK7_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[1]\, 
        \U_ELK7_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[2]\, 
        \U_ELK7_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[3]\, 
        \U_ELK7_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[4]\, 
        \U_ELK7_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[5]\, 
        \U_ELK7_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[6]\, 
        \U_ELK7_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[7]\, 
        \U_ELK7_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/Q[0]_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/Q[1]_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/Q[2]_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/Q[3]_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/Q[4]_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/Q[5]_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/Q[6]_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/Q[7]_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/Q[8]_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/Q[9]_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/Q[10]_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/Q[11]_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/Q[12]_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/Q[13]_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[13]_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/Q[14]_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[14]_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]_net_1\, 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]_net_1\, 
        \U_ELK14_CH/ELK_IN_F_net_1\, \U_ELK14_CH/ELK_IN_DDR_F\, 
        \U_ELK14_CH/ELK_IN_R_net_1\, \U_ELK14_CH/ELK_IN_DDR_R\, 
        \U_ELK14_CH/ELK_OUT_F\, \U_ELK14_CH/ELK_OUT_R\, 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[0]_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[1]_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[2]_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[3]_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[11]_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[12]_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[13]_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[14]_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[0]\, 
        \U_ELK14_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[1]\, 
        \U_ELK14_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[2]\, 
        \U_ELK14_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[3]\, 
        \U_ELK14_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[4]\, 
        \U_ELK14_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[5]\, 
        \U_ELK14_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[6]\, 
        \U_ELK14_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[7]\, 
        \U_ELK14_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/Q[0]_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/Q[1]_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/Q[2]_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/Q[3]_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/Q[4]_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/Q[5]_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/Q[6]_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/Q[7]_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/Q[8]_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/Q[9]_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/Q[10]_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/Q[11]_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/Q[12]_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/Q[13]_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[13]_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/Q[14]_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[14]_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]_net_1\, 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]_net_1\, 
        \U_ELK2_CH/ELK_IN_F_net_1\, \U_ELK2_CH/ELK_IN_DDR_F\, 
        \U_ELK2_CH/ELK_IN_R_net_1\, \U_ELK2_CH/ELK_IN_DDR_R\, 
        \U_ELK2_CH/ELK_OUT_F\, \U_ELK2_CH/ELK_OUT_R\, 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[0]_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[1]_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[2]_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[3]_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[11]_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[12]_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[13]_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[14]_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[0]\, 
        \U_ELK2_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[1]\, 
        \U_ELK2_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[2]\, 
        \U_ELK2_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[3]\, 
        \U_ELK2_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[4]\, 
        \U_ELK2_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[5]\, 
        \U_ELK2_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[6]\, 
        \U_ELK2_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[7]\, 
        \U_ELK2_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/Q[0]_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/Q[1]_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/Q[2]_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/Q[3]_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/Q[4]_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/Q[5]_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/Q[6]_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/Q[7]_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/Q[8]_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/Q[9]_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/Q[10]_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/Q[11]_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/Q[12]_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/Q[13]_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[13]_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/Q[14]_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[14]_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]_net_1\, 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]_net_1\, 
        \U_ELK4_CH/ELK_IN_F_net_1\, \U_ELK4_CH/ELK_IN_R_net_1\, 
        \U_ELK4_CH/ELK_OUT_F_i_0\, \U_ELK4_CH/ELK_OUT_R_i_0\, 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[0]_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[1]_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[2]_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[3]_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[11]_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[12]_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[13]_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[14]_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[0]\, 
        \U_ELK4_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[1]\, 
        \U_ELK4_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[2]\, 
        \U_ELK4_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[3]\, 
        \U_ELK4_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[4]\, 
        \U_ELK4_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[5]\, 
        \U_ELK4_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[6]\, 
        \U_ELK4_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[7]\, 
        \U_ELK4_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/Q[0]_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/Q[1]_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/Q[2]_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/Q[3]_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/Q[4]_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/Q[5]_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/Q[6]_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/Q[7]_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/Q[8]_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/Q[9]_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/Q[10]_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/Q[11]_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/Q[12]_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/Q[13]_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[13]_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/Q[14]_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[14]_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]_net_1\, 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]_net_1\, 
        \U_ELK4_CH/U_DDR_ELK1/ELK_IN_DDR_R\, 
        \U_ELK4_CH/U_DDR_ELK1/ELK_IN_DDR_F\, 
        \U_ELK6_CH/ELK_IN_F_net_1\, \U_ELK6_CH/ELK_IN_DDR_F\, 
        \U_ELK6_CH/ELK_IN_R_net_1\, \U_ELK6_CH/ELK_IN_DDR_R\, 
        \U_ELK6_CH/ELK_OUT_F\, \U_ELK6_CH/ELK_OUT_R\, 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[0]_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[1]_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[2]_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[3]_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[11]_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[12]_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[13]_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[14]_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[0]\, 
        \U_ELK6_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[1]\, 
        \U_ELK6_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[2]\, 
        \U_ELK6_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[3]\, 
        \U_ELK6_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[4]\, 
        \U_ELK6_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[5]\, 
        \U_ELK6_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[6]\, 
        \U_ELK6_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[7]\, 
        \U_ELK6_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/Q[0]_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/Q[1]_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/Q[2]_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/Q[3]_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/Q[4]_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/Q[5]_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/Q[6]_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/Q[7]_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/Q[8]_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/Q[9]_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/Q[10]_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/Q[11]_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/Q[12]_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/Q[13]_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[13]_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/Q[14]_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[14]_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]_net_1\, 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]_net_1\, 
        \U_MASTER_DES/AUX_MODE\, \U_MASTER_DES/AUX_SDIN\, 
        \U_MASTER_DES/AUX_SUPDATE\, \U_MASTER_DES/AUX_SSHIFT\, 
        \U_MASTER_DES/CCC_RX_CLK_LOCK\, 
        \U_ELK16_CH/ELK_IN_F_net_1\, \U_ELK16_CH/ELK_IN_DDR_F\, 
        \U_ELK16_CH/ELK_IN_R_net_1\, \U_ELK16_CH/ELK_IN_DDR_R\, 
        \U_ELK16_CH/ELK_OUT_F\, \U_ELK16_CH/ELK_OUT_R\, 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[0]_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[1]_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[2]_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[3]_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[11]_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[12]_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[13]_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[14]_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[0]\, 
        \U_ELK16_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[1]\, 
        \U_ELK16_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[2]\, 
        \U_ELK16_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[3]\, 
        \U_ELK16_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[4]\, 
        \U_ELK16_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[5]\, 
        \U_ELK16_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[6]\, 
        \U_ELK16_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[7]\, 
        \U_ELK16_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/Q[0]_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/Q[1]_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/Q[2]_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/Q[3]_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/Q[4]_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/Q[5]_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/Q[6]_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/Q[7]_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/Q[8]_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/Q[9]_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/Q[10]_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/Q[11]_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/Q[12]_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/Q[13]_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[13]_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/Q[14]_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[14]_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]_net_1\, 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]_net_1\, 
        \U_DDR_ELK0/ELK0_IN_DDR_R\, \U_DDR_ELK0/ELK0_IN_DDR_F\, 
        \U_ELK19_CH/ELK_IN_F_net_1\, \U_ELK19_CH/ELK_IN_DDR_F\, 
        \U_ELK19_CH/ELK_IN_R_net_1\, \U_ELK19_CH/ELK_IN_DDR_R\, 
        \U_ELK19_CH/ELK_OUT_F\, \U_ELK19_CH/ELK_OUT_R\, 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[0]_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[1]_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[2]_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[3]_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[11]_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[12]_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[13]_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[14]_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[0]\, 
        \U_ELK19_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[1]\, 
        \U_ELK19_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[2]\, 
        \U_ELK19_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[3]\, 
        \U_ELK19_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[4]\, 
        \U_ELK19_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[5]\, 
        \U_ELK19_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[6]\, 
        \U_ELK19_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[7]\, 
        \U_ELK19_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/Q[0]_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/Q[1]_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/Q[2]_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/Q[3]_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/Q[4]_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/Q[5]_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/Q[6]_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/Q[7]_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/Q[8]_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/Q[9]_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/Q[10]_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/Q[11]_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/Q[12]_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/Q[13]_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[13]_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/Q[14]_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[14]_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]_net_1\, 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]_net_1\, 
        \U_ELK9_CH/ELK_IN_F_net_1\, \U_ELK9_CH/ELK_IN_DDR_F\, 
        \U_ELK9_CH/ELK_IN_R_net_1\, \U_ELK9_CH/ELK_IN_DDR_R\, 
        \U_ELK9_CH/ELK_OUT_F\, \U_ELK9_CH/ELK_OUT_R\, 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[0]_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[1]_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[2]_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[3]_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[11]_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[12]_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[13]_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[14]_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[0]\, 
        \U_ELK9_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[1]\, 
        \U_ELK9_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[2]\, 
        \U_ELK9_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[3]\, 
        \U_ELK9_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[4]\, 
        \U_ELK9_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[5]\, 
        \U_ELK9_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[6]\, 
        \U_ELK9_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[7]\, 
        \U_ELK9_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/Q[0]_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/Q[1]_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/Q[2]_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/Q[3]_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/Q[4]_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/Q[5]_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/Q[6]_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/Q[7]_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/Q[8]_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/Q[9]_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/Q[10]_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/Q[11]_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/Q[12]_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/Q[13]_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[13]_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/Q[14]_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[14]_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]_net_1\, 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]_net_1\, 
        \U_ELK8_CH/ELK_IN_F_net_1\, \U_ELK8_CH/ELK_IN_DDR_F\, 
        \U_ELK8_CH/ELK_IN_R_net_1\, \U_ELK8_CH/ELK_IN_DDR_R\, 
        \U_ELK8_CH/ELK_OUT_F\, \U_ELK8_CH/ELK_OUT_R\, 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[0]_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[1]_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[2]_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[3]_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[11]_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[12]_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[13]_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[14]_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[0]\, 
        \U_ELK8_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[1]\, 
        \U_ELK8_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[2]\, 
        \U_ELK8_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[3]\, 
        \U_ELK8_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[4]\, 
        \U_ELK8_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[5]\, 
        \U_ELK8_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[6]\, 
        \U_ELK8_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[7]\, 
        \U_ELK8_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/Q[0]_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/Q[1]_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/Q[2]_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/Q[3]_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/Q[4]_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/Q[5]_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/Q[6]_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/Q[7]_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/Q[8]_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/Q[9]_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/Q[10]_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/Q[11]_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/Q[12]_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/Q[13]_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[13]_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/Q[14]_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[14]_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]_net_1\, 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]_net_1\, 
        \U_ELK17_CH/ELK_IN_F_net_1\, \U_ELK17_CH/ELK_IN_DDR_F\, 
        \U_ELK17_CH/ELK_IN_R_net_1\, \U_ELK17_CH/ELK_IN_DDR_R\, 
        \U_ELK17_CH/ELK_OUT_F\, \U_ELK17_CH/ELK_OUT_R\, 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[0]_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[1]_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[2]_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[3]_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[11]_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[12]_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[13]_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[14]_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[0]\, 
        \U_ELK17_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[1]\, 
        \U_ELK17_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[2]\, 
        \U_ELK17_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[3]\, 
        \U_ELK17_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[4]\, 
        \U_ELK17_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[5]\, 
        \U_ELK17_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[6]\, 
        \U_ELK17_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[7]\, 
        \U_ELK17_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/Q[0]_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/Q[1]_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/Q[2]_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/Q[3]_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/Q[4]_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/Q[5]_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/Q[6]_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/Q[7]_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/Q[8]_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/Q[9]_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/Q[10]_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/Q[11]_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/Q[12]_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/Q[13]_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[13]_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/Q[14]_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[14]_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]_net_1\, 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]_net_1\, 
        \U_ELK15_CH/ELK_IN_F_net_1\, \U_ELK15_CH/ELK_IN_DDR_F\, 
        \U_ELK15_CH/ELK_IN_R_net_1\, \U_ELK15_CH/ELK_IN_DDR_R\, 
        \U_ELK15_CH/ELK_OUT_F\, \U_ELK15_CH/ELK_OUT_R\, 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[0]_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[1]_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[2]_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[3]_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[11]_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[12]_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[13]_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[14]_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[0]\, 
        \U_ELK15_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[1]\, 
        \U_ELK15_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[2]\, 
        \U_ELK15_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[3]\, 
        \U_ELK15_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[4]\, 
        \U_ELK15_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[5]\, 
        \U_ELK15_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[6]\, 
        \U_ELK15_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[7]\, 
        \U_ELK15_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/Q[0]_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/Q[1]_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/Q[2]_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/Q[3]_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/Q[4]_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/Q[5]_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/Q[6]_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/Q[7]_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/Q[8]_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/Q[9]_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/Q[10]_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/Q[11]_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/Q[12]_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/Q[13]_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[13]_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/Q[14]_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[14]_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]_net_1\, 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]_net_1\, 
        \U_ELK5_CH/ELK_IN_F_net_1\, \U_ELK5_CH/ELK_IN_DDR_F\, 
        \U_ELK5_CH/ELK_IN_R_net_1\, \U_ELK5_CH/ELK_IN_DDR_R\, 
        \U_ELK5_CH/ELK_OUT_F\, \U_ELK5_CH/ELK_OUT_R\, 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[0]_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[1]_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[2]_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[3]_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[11]_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[12]_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[13]_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[14]_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[0]\, 
        \U_ELK5_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[1]\, 
        \U_ELK5_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[2]\, 
        \U_ELK5_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[3]\, 
        \U_ELK5_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[4]\, 
        \U_ELK5_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[5]\, 
        \U_ELK5_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[6]\, 
        \U_ELK5_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[7]\, 
        \U_ELK5_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/Q[0]_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/Q[1]_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/Q[2]_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/Q[3]_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/Q[4]_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/Q[5]_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/Q[6]_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/Q[7]_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/Q[8]_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/Q[9]_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/Q[10]_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/Q[11]_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/Q[12]_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/Q[13]_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[13]_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/Q[14]_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[14]_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]_net_1\, 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]_net_1\, 
        \U_ELK10_CH/ELK_IN_F_net_1\, \U_ELK10_CH/ELK_IN_DDR_F\, 
        \U_ELK10_CH/ELK_IN_R_net_1\, \U_ELK10_CH/ELK_IN_DDR_R\, 
        \U_ELK10_CH/ELK_OUT_F\, \U_ELK10_CH/ELK_OUT_R\, 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[0]_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[1]_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[2]_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[3]_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[11]_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[12]_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[13]_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[14]_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[0]\, 
        \U_ELK10_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[1]\, 
        \U_ELK10_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[2]\, 
        \U_ELK10_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[3]\, 
        \U_ELK10_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[4]\, 
        \U_ELK10_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[5]\, 
        \U_ELK10_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[6]\, 
        \U_ELK10_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[7]\, 
        \U_ELK10_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/Q[0]_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/Q[1]_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/Q[2]_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/Q[3]_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/Q[4]_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/Q[5]_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/Q[6]_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/Q[7]_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/Q[8]_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/Q[9]_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/Q[10]_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/Q[11]_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/Q[12]_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/Q[13]_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[13]_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/Q[14]_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[14]_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]_net_1\, 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]_net_1\, 
        \USBCLK60MHZ_pad/U0/NET1\, 
        \U60_TS_RD_BUF/\\\\TRIBUFF_F_24U[0]\\\\/U0/NET1\, 
        \U60_TS_RD_BUF/\\\\TRIBUFF_F_24U[0]\\\\/U0/NET2\, 
        \U_ELK13_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2_N2P\, 
        \U_ELK13_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, 
        \U_ELK13_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET2\, 
        \U_ELK13_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET3\, 
        \U_ELK13_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\, 
        \DEV_RST_B_pad/U0/NET1\, 
        \U_ELK16_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2_N2P\, 
        \U_ELK16_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, 
        \U_ELK16_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET2\, 
        \U_ELK16_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET3\, 
        \U_ELK16_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\, 
        \U_ELK19_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2_N2P\, 
        \U_ELK19_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, 
        \U_ELK19_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET2\, 
        \U_ELK19_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET3\, 
        \U_ELK19_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\, 
        \U_DDR_TFC/BIBUF_LVDS_0/U0/U2_N2P\, 
        \U_DDR_TFC/BIBUF_LVDS_0/U0/NET1\, 
        \U_DDR_TFC/BIBUF_LVDS_0/U0/NET2\, 
        \U_DDR_TFC/BIBUF_LVDS_0/U0/NET3\, 
        \U_DDR_TFC/BIBUF_LVDS_0/U0/NET4\, 
        \U_ELK6_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2_N2P\, 
        \U_ELK6_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, 
        \U_ELK6_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET2\, 
        \U_ELK6_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET3\, 
        \U_ELK6_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\, 
        \U0A_40M_REFCLK/\\\\BIBUF_LVDS[0]\\\\/U0/U2_N2P\, 
        \U0A_40M_REFCLK/\\\\BIBUF_LVDS[0]\\\\/U0/NET1\, 
        \U0A_40M_REFCLK/\\\\BIBUF_LVDS[0]\\\\/U0/NET2\, 
        \U0A_40M_REFCLK/\\\\BIBUF_LVDS[0]\\\\/U0/NET3\, 
        \U0A_40M_REFCLK/\\\\BIBUF_LVDS[0]\\\\/U0/NET4\, 
        \U_ELK7_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2_N2P\, 
        \U_ELK7_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, 
        \U_ELK7_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET2\, 
        \U_ELK7_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET3\, 
        \U_ELK7_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\, 
        \P_USB_RXF_B_pad/U0/NET1\, 
        \U_ELK15_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2_N2P\, 
        \U_ELK15_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, 
        \U_ELK15_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET2\, 
        \U_ELK15_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET3\, 
        \U_ELK15_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\, 
        \P_OP_MODE5_AAE_pad/U0/NET1\, 
        \P_OP_MODE5_AAE_pad/U0/NET2\, \ALL_PLL_LOCK_pad/U0/NET1\, 
        \ALL_PLL_LOCK_pad/U0/NET2\, \P_ELK0_SYNC_DET_pad/U0/NET1\, 
        \P_ELK0_SYNC_DET_pad/U0/NET2\, 
        \U_ELK4_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2_N2P\, 
        \U_ELK4_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, 
        \U_ELK4_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET2\, 
        \U_ELK4_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET3\, 
        \U_ELK4_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\, 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[0]\\\\/U0/NET1\, 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[0]\\\\/U0/NET2\, 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[0]\\\\/U0/NET3\, 
        \P_OP_MODE6_EE_pad/U0/NET1\, \P_OP_MODE6_EE_pad/U0/NET2\, 
        \P_OP_MODE2_TE_pad/U0/NET1\, \P_OP_MODE2_TE_pad/U0/NET2\, 
        \U_DDR_ELK0/BIBUF_LVDS_0/U0/U2_N2P\, 
        \U_DDR_ELK0/BIBUF_LVDS_0/U0/NET1\, 
        \U_DDR_ELK0/BIBUF_LVDS_0/U0/NET2\, 
        \U_DDR_ELK0/BIBUF_LVDS_0/U0/NET3\, 
        \U_DDR_ELK0/BIBUF_LVDS_0/U0/NET4\, 
        \U_ELK10_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2_N2P\, 
        \U_ELK10_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, 
        \U_ELK10_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET2\, 
        \U_ELK10_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET3\, 
        \U_ELK10_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\, 
        \P_TFC_SYNC_DET_pad/U0/NET1\, 
        \P_TFC_SYNC_DET_pad/U0/NET2\, 
        \U_ELK12_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2_N2P\, 
        \U_ELK12_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, 
        \U_ELK12_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET2\, 
        \U_ELK12_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET3\, 
        \U_ELK12_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\, 
        \P_MASTER_POR_B_pad/U0/NET1\, 
        \P_MASTER_POR_B_pad/U0/NET2\, 
        \U63_TS_SIWU_BUF/\\\\TRIBUFF_F_24U[0]\\\\/U0/NET1\, 
        \U63_TS_SIWU_BUF/\\\\TRIBUFF_F_24U[0]\\\\/U0/NET2\, 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[6]\\\\/U0/NET1\, 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[6]\\\\/U0/NET2\, 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[6]\\\\/U0/NET3\, 
        \U_ELK3_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2_N2P\, 
        \U_ELK3_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, 
        \U_ELK3_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET2\, 
        \U_ELK3_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET3\, 
        \U_ELK3_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\, 
        \P_OP_MODE1_SPE_pad/U0/NET1\, 
        \P_OP_MODE1_SPE_pad/U0/NET2\, 
        \U0B_TX40M_REFCLK/\\\\OUTBUF_LVDS[0]\\\\/U0/NET1\, 
        \U0B_TX40M_REFCLK/\\\\OUTBUF_LVDS[0]\\\\/U0/NET2\, 
        \U_ELK5_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2_N2P\, 
        \U_ELK5_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, 
        \U_ELK5_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET2\, 
        \U_ELK5_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET3\, 
        \U_ELK5_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\, 
        \P_USB_MASTER_EN_pad/U0/NET1\, 
        \P_USB_MASTER_EN_pad/U0/NET2\, \P_USB_TXE_B_pad/U0/NET1\, 
        \U_ELK17_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2_N2P\, 
        \U_ELK17_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, 
        \U_ELK17_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET2\, 
        \U_ELK17_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET3\, 
        \U_ELK17_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\, 
        \P_CLK_40M_GL_pad/U0/NET1\, \P_CLK_40M_GL_pad/U0/NET2\, 
        \U_ELK1_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2_N2P\, 
        \U_ELK1_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, 
        \U_ELK1_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET2\, 
        \U_ELK1_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET3\, 
        \U_ELK1_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\, 
        \U_ELK14_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2_N2P\, 
        \U_ELK14_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, 
        \U_ELK14_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET2\, 
        \U_ELK14_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET3\, 
        \U_ELK14_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\, 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[3]\\\\/U0/NET1\, 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[3]\\\\/U0/NET2\, 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[3]\\\\/U0/NET3\, 
        \U62_TS_OE_BUF/\\\\TRIBUFF_F_24U[0]\\\\/U0/NET1\, 
        \U62_TS_OE_BUF/\\\\TRIBUFF_F_24U[0]\\\\/U0/NET2\, 
        \U_ELK8_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2_N2P\, 
        \U_ELK8_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, 
        \U_ELK8_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET2\, 
        \U_ELK8_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET3\, 
        \U_ELK8_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\, 
        \U_ELK11_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2_N2P\, 
        \U_ELK11_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, 
        \U_ELK11_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET2\, 
        \U_ELK11_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET3\, 
        \U_ELK11_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\, 
        \P_CCC_160M_FXD_pad/U0/NET1\, 
        \P_CCC_160M_FXD_pad/U0/NET2\, 
        \U_REFCLKBUF/\\\\BIBUF_LVDS[0]\\\\/U0/U2_N2P\, 
        \U_REFCLKBUF/\\\\BIBUF_LVDS[0]\\\\/U0/NET1\, 
        \U_REFCLKBUF/\\\\BIBUF_LVDS[0]\\\\/U0/NET2\, 
        \U_REFCLKBUF/\\\\BIBUF_LVDS[0]\\\\/U0/NET3\, 
        \U_REFCLKBUF/\\\\BIBUF_LVDS[0]\\\\/U0/NET4\, 
        \U_ELK2_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2_N2P\, 
        \U_ELK2_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, 
        \U_ELK2_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET2\, 
        \U_ELK2_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET3\, 
        \U_ELK2_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\, 
        \U_ELK9_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2_N2P\, 
        \U_ELK9_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, 
        \U_ELK9_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET2\, 
        \U_ELK9_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET3\, 
        \U_ELK9_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\, 
        \P_CCC_160M_ADJ_pad/U0/NET1\, 
        \P_CCC_160M_ADJ_pad/U0/NET2\, 
        \U61_TS_WR_BUF/\\\\TRIBUFF_F_24U[0]\\\\/U0/NET1\, 
        \U61_TS_WR_BUF/\\\\TRIBUFF_F_24U[0]\\\\/U0/NET2\, 
        \U_ELK18_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2_N2P\, 
        \U_ELK18_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, 
        \U_ELK18_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET2\, 
        \U_ELK18_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET3\, 
        \U_ELK18_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\, 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[4]\\\\/U0/NET1\, 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[4]\\\\/U0/NET2\, 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[4]\\\\/U0/NET3\, 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[7]\\\\/U0/NET1\, 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[7]\\\\/U0/NET2\, 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[7]\\\\/U0/NET3\, 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[2]\\\\/U0/NET1\, 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[2]\\\\/U0/NET2\, 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[2]\\\\/U0/NET3\, 
        \DCB_SALT_SEL_pad/U0/NET1\, 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[1]\\\\/U0/NET1\, 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[1]\\\\/U0/NET2\, 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[1]\\\\/U0/NET3\, 
        \U0_200M_BUF/\\\\INBUF_LVDS[0]\\\\/U0/U2_N2P\, 
        \U0_200M_BUF/\\\\INBUF_LVDS[0]\\\\/U0/NET1\, 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[5]\\\\/U0/NET1\, 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[5]\\\\/U0/NET2\, 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[5]\\\\/U0/NET3\, 
        \EXTCLK_40MHZ_pad/U0/NET1\, \EXTCLK_40MHZ_pad/U0/NET2\, 
        \EXT_INT_REF_SEL_pad/U0/NET1\, ALIGN_ACTIVE, 
        \BIT_OS_SEL[0]\, \BIT_OS_SEL[1]\, \BIT_OS_SEL[2]\, 
        \BIT_OS_SEL_0[0]\, \BIT_OS_SEL_0[1]\, \BIT_OS_SEL_0[2]\, 
        \BIT_OS_SEL_1[0]\, \BIT_OS_SEL_1[1]\, \BIT_OS_SEL_1[2]\, 
        \BIT_OS_SEL_2[0]\, \BIT_OS_SEL_2[1]\, \BIT_OS_SEL_2[2]\, 
        \BIT_OS_SEL_3[0]\, \BIT_OS_SEL_3[1]\, \BIT_OS_SEL_3[2]\, 
        \BIT_OS_SEL_4[0]\, \BIT_OS_SEL_4[1]\, \BIT_OS_SEL_4[2]\, 
        \BIT_OS_SEL_5[0]\, \BIT_OS_SEL_5[1]\, \BIT_OS_SEL_5[2]\, 
        \BIT_OS_SEL_6[1]\, \BIT_OS_SEL_6[2]\, \BIT_OS_SEL_7[2]\, 
        \ELK0_IN_F\, \ELK0_IN_R\, \ELK0_TX_DAT[0]\, 
        \ELK0_TX_DAT[1]\, \ELK0_TX_DAT[2]\, \ELK0_TX_DAT[3]\, 
        \ELK0_TX_DAT[4]\, \ELK0_TX_DAT[5]\, \ELK0_TX_DAT[6]\, 
        \ELK0_TX_DAT[7]\, \ELKS_STOP_ADDR[0]\, 
        \ELKS_STOP_ADDR[1]\, \ELKS_STOP_ADDR[2]\, 
        \ELKS_STOP_ADDR[3]\, \ELKS_STOP_ADDR[4]\, 
        \ELKS_STOP_ADDR[5]\, \ELKS_STOP_ADDR[6]\, 
        \ELKS_STOP_ADDR[7]\, \ELKS_STRT_ADDR[0]\, 
        \ELKS_STRT_ADDR[1]\, \ELKS_STRT_ADDR[2]\, 
        \ELKS_STRT_ADDR[3]\, \ELKS_STRT_ADDR[4]\, 
        \ELKS_STRT_ADDR[5]\, \ELKS_STRT_ADDR[6]\, 
        \ELKS_STRT_ADDR[7]\, HIEFFPLA_NET_0_115805, 
        HIEFFPLA_NET_0_115806, HIEFFPLA_NET_0_115807, 
        HIEFFPLA_NET_0_115808, HIEFFPLA_NET_0_115809, 
        HIEFFPLA_NET_0_115810, HIEFFPLA_NET_0_115811, 
        HIEFFPLA_NET_0_115812, HIEFFPLA_NET_0_115813, 
        HIEFFPLA_NET_0_115814, HIEFFPLA_NET_0_115815, 
        HIEFFPLA_NET_0_115816, HIEFFPLA_NET_0_115817, 
        HIEFFPLA_NET_0_115818, HIEFFPLA_NET_0_115819, 
        HIEFFPLA_NET_0_115820, HIEFFPLA_NET_0_115821, 
        HIEFFPLA_NET_0_115822, HIEFFPLA_NET_0_115823, 
        HIEFFPLA_NET_0_115824, HIEFFPLA_NET_0_115825, 
        HIEFFPLA_NET_0_115826, HIEFFPLA_NET_0_115827, 
        HIEFFPLA_NET_0_115828, HIEFFPLA_NET_0_115829, 
        HIEFFPLA_NET_0_115830, HIEFFPLA_NET_0_115831, 
        HIEFFPLA_NET_0_115832, HIEFFPLA_NET_0_115833, 
        HIEFFPLA_NET_0_115834, HIEFFPLA_NET_0_115835, 
        HIEFFPLA_NET_0_115836, HIEFFPLA_NET_0_115837, 
        HIEFFPLA_NET_0_115838, HIEFFPLA_NET_0_115839, 
        HIEFFPLA_NET_0_115840, HIEFFPLA_NET_0_115841, 
        HIEFFPLA_NET_0_115842, HIEFFPLA_NET_0_115843, 
        HIEFFPLA_NET_0_115844, HIEFFPLA_NET_0_115845, 
        HIEFFPLA_NET_0_115846, HIEFFPLA_NET_0_115847, 
        HIEFFPLA_NET_0_115848, HIEFFPLA_NET_0_115866, 
        HIEFFPLA_NET_0_115867, HIEFFPLA_NET_0_115868, 
        HIEFFPLA_NET_0_115869, HIEFFPLA_NET_0_115870, 
        HIEFFPLA_NET_0_115871, HIEFFPLA_NET_0_115872, 
        HIEFFPLA_NET_0_115873, HIEFFPLA_NET_0_115874, 
        HIEFFPLA_NET_0_115875, HIEFFPLA_NET_0_115876, 
        HIEFFPLA_NET_0_115877, HIEFFPLA_NET_0_115878, 
        HIEFFPLA_NET_0_115879, HIEFFPLA_NET_0_115880, 
        HIEFFPLA_NET_0_115881, HIEFFPLA_NET_0_115882, 
        HIEFFPLA_NET_0_115883, HIEFFPLA_NET_0_115884, 
        HIEFFPLA_NET_0_115885, HIEFFPLA_NET_0_115886, 
        HIEFFPLA_NET_0_115887, HIEFFPLA_NET_0_115888, 
        HIEFFPLA_NET_0_115889, HIEFFPLA_NET_0_115890, 
        HIEFFPLA_NET_0_115891, HIEFFPLA_NET_0_115892, 
        HIEFFPLA_NET_0_115893, HIEFFPLA_NET_0_115894, 
        HIEFFPLA_NET_0_115895, HIEFFPLA_NET_0_115896, 
        HIEFFPLA_NET_0_115897, HIEFFPLA_NET_0_115898, 
        HIEFFPLA_NET_0_115899, HIEFFPLA_NET_0_115900, 
        HIEFFPLA_NET_0_115901, HIEFFPLA_NET_0_115902, 
        HIEFFPLA_NET_0_115903, HIEFFPLA_NET_0_115904, 
        HIEFFPLA_NET_0_115905, HIEFFPLA_NET_0_115906, 
        HIEFFPLA_NET_0_115907, HIEFFPLA_NET_0_115908, 
        HIEFFPLA_NET_0_115909, HIEFFPLA_NET_0_115910, 
        HIEFFPLA_NET_0_115911, HIEFFPLA_NET_0_115912, 
        HIEFFPLA_NET_0_115913, HIEFFPLA_NET_0_115914, 
        HIEFFPLA_NET_0_115915, HIEFFPLA_NET_0_115916, 
        HIEFFPLA_NET_0_115917, HIEFFPLA_NET_0_115918, 
        HIEFFPLA_NET_0_115919, HIEFFPLA_NET_0_115920, 
        HIEFFPLA_NET_0_115921, HIEFFPLA_NET_0_115922, 
        HIEFFPLA_NET_0_115923, HIEFFPLA_NET_0_115924, 
        HIEFFPLA_NET_0_115925, HIEFFPLA_NET_0_115926, 
        HIEFFPLA_NET_0_115927, HIEFFPLA_NET_0_115928, 
        HIEFFPLA_NET_0_115929, HIEFFPLA_NET_0_115930, 
        HIEFFPLA_NET_0_115931, HIEFFPLA_NET_0_115932, 
        HIEFFPLA_NET_0_115933, HIEFFPLA_NET_0_115934, 
        HIEFFPLA_NET_0_115935, HIEFFPLA_NET_0_115936, 
        HIEFFPLA_NET_0_115937, HIEFFPLA_NET_0_115938, 
        HIEFFPLA_NET_0_115939, HIEFFPLA_NET_0_115940, 
        HIEFFPLA_NET_0_115941, HIEFFPLA_NET_0_115942, 
        HIEFFPLA_NET_0_115943, HIEFFPLA_NET_0_115944, 
        HIEFFPLA_NET_0_115945, HIEFFPLA_NET_0_115946, 
        HIEFFPLA_NET_0_115947, HIEFFPLA_NET_0_115948, 
        HIEFFPLA_NET_0_115949, HIEFFPLA_NET_0_115950, 
        HIEFFPLA_NET_0_115951, HIEFFPLA_NET_0_115952, 
        HIEFFPLA_NET_0_115953, HIEFFPLA_NET_0_115954, 
        HIEFFPLA_NET_0_115955, HIEFFPLA_NET_0_115956, 
        HIEFFPLA_NET_0_115957, HIEFFPLA_NET_0_115958, 
        HIEFFPLA_NET_0_115959, HIEFFPLA_NET_0_115960, 
        HIEFFPLA_NET_0_115961, HIEFFPLA_NET_0_115962, 
        HIEFFPLA_NET_0_115963, HIEFFPLA_NET_0_115964, 
        HIEFFPLA_NET_0_115965, HIEFFPLA_NET_0_115966, 
        HIEFFPLA_NET_0_115967, HIEFFPLA_NET_0_115968, 
        HIEFFPLA_NET_0_115969, HIEFFPLA_NET_0_115970, 
        HIEFFPLA_NET_0_115971, HIEFFPLA_NET_0_115972, 
        HIEFFPLA_NET_0_115973, HIEFFPLA_NET_0_115974, 
        HIEFFPLA_NET_0_115975, HIEFFPLA_NET_0_115976, 
        HIEFFPLA_NET_0_115977, HIEFFPLA_NET_0_115978, 
        HIEFFPLA_NET_0_115979, HIEFFPLA_NET_0_115980, 
        HIEFFPLA_NET_0_115981, HIEFFPLA_NET_0_115982, 
        HIEFFPLA_NET_0_115983, HIEFFPLA_NET_0_115984, 
        HIEFFPLA_NET_0_115985, HIEFFPLA_NET_0_115986, 
        HIEFFPLA_NET_0_115987, HIEFFPLA_NET_0_115988, 
        HIEFFPLA_NET_0_115989, HIEFFPLA_NET_0_115990, 
        HIEFFPLA_NET_0_115991, HIEFFPLA_NET_0_115992, 
        HIEFFPLA_NET_0_115993, HIEFFPLA_NET_0_115994, 
        HIEFFPLA_NET_0_115995, HIEFFPLA_NET_0_115996, 
        HIEFFPLA_NET_0_115997, HIEFFPLA_NET_0_115998, 
        HIEFFPLA_NET_0_115999, HIEFFPLA_NET_0_116000, 
        HIEFFPLA_NET_0_116001, HIEFFPLA_NET_0_116002, 
        HIEFFPLA_NET_0_116003, HIEFFPLA_NET_0_116004, 
        HIEFFPLA_NET_0_116005, HIEFFPLA_NET_0_116006, 
        HIEFFPLA_NET_0_116007, HIEFFPLA_NET_0_116008, 
        HIEFFPLA_NET_0_116009, HIEFFPLA_NET_0_116010, 
        HIEFFPLA_NET_0_116011, HIEFFPLA_NET_0_116012, 
        HIEFFPLA_NET_0_116013, HIEFFPLA_NET_0_116014, 
        HIEFFPLA_NET_0_116015, HIEFFPLA_NET_0_116016, 
        HIEFFPLA_NET_0_116017, HIEFFPLA_NET_0_116018, 
        HIEFFPLA_NET_0_116019, HIEFFPLA_NET_0_116020, 
        HIEFFPLA_NET_0_116021, HIEFFPLA_NET_0_116022, 
        HIEFFPLA_NET_0_116023, HIEFFPLA_NET_0_116024, 
        HIEFFPLA_NET_0_116025, HIEFFPLA_NET_0_116026, 
        HIEFFPLA_NET_0_116027, HIEFFPLA_NET_0_116028, 
        HIEFFPLA_NET_0_116029, HIEFFPLA_NET_0_116030, 
        HIEFFPLA_NET_0_116031, HIEFFPLA_NET_0_116032, 
        HIEFFPLA_NET_0_116033, HIEFFPLA_NET_0_116034, 
        HIEFFPLA_NET_0_116035, HIEFFPLA_NET_0_116036, 
        HIEFFPLA_NET_0_116037, HIEFFPLA_NET_0_116038, 
        HIEFFPLA_NET_0_116039, HIEFFPLA_NET_0_116040, 
        HIEFFPLA_NET_0_116041, HIEFFPLA_NET_0_116042, 
        HIEFFPLA_NET_0_116043, HIEFFPLA_NET_0_116044, 
        HIEFFPLA_NET_0_116045, HIEFFPLA_NET_0_116046, 
        HIEFFPLA_NET_0_116047, HIEFFPLA_NET_0_116048, 
        HIEFFPLA_NET_0_116049, HIEFFPLA_NET_0_116050, 
        HIEFFPLA_NET_0_116051, HIEFFPLA_NET_0_116052, 
        HIEFFPLA_NET_0_116053, HIEFFPLA_NET_0_116054, 
        HIEFFPLA_NET_0_116055, HIEFFPLA_NET_0_116056, 
        HIEFFPLA_NET_0_116057, HIEFFPLA_NET_0_116058, 
        HIEFFPLA_NET_0_116059, HIEFFPLA_NET_0_116060, 
        HIEFFPLA_NET_0_116061, HIEFFPLA_NET_0_116062, 
        HIEFFPLA_NET_0_116063, HIEFFPLA_NET_0_116064, 
        HIEFFPLA_NET_0_116065, HIEFFPLA_NET_0_116066, 
        HIEFFPLA_NET_0_116067, HIEFFPLA_NET_0_116068, 
        HIEFFPLA_NET_0_116069, HIEFFPLA_NET_0_116070, 
        HIEFFPLA_NET_0_116071, HIEFFPLA_NET_0_116072, 
        HIEFFPLA_NET_0_116073, HIEFFPLA_NET_0_116074, 
        HIEFFPLA_NET_0_116075, HIEFFPLA_NET_0_116076, 
        HIEFFPLA_NET_0_116077, HIEFFPLA_NET_0_116078, 
        HIEFFPLA_NET_0_116079, HIEFFPLA_NET_0_116080, 
        HIEFFPLA_NET_0_116081, HIEFFPLA_NET_0_116082, 
        HIEFFPLA_NET_0_116083, HIEFFPLA_NET_0_116084, 
        HIEFFPLA_NET_0_116085, HIEFFPLA_NET_0_116086, 
        HIEFFPLA_NET_0_116087, HIEFFPLA_NET_0_116088, 
        HIEFFPLA_NET_0_116089, HIEFFPLA_NET_0_116090, 
        HIEFFPLA_NET_0_116091, HIEFFPLA_NET_0_116092, 
        HIEFFPLA_NET_0_116093, HIEFFPLA_NET_0_116094, 
        HIEFFPLA_NET_0_116095, HIEFFPLA_NET_0_116096, 
        HIEFFPLA_NET_0_116097, HIEFFPLA_NET_0_116098, 
        HIEFFPLA_NET_0_116099, HIEFFPLA_NET_0_116100, 
        HIEFFPLA_NET_0_116101, HIEFFPLA_NET_0_116102, 
        HIEFFPLA_NET_0_116103, HIEFFPLA_NET_0_116104, 
        HIEFFPLA_NET_0_116105, HIEFFPLA_NET_0_116106, 
        HIEFFPLA_NET_0_116107, HIEFFPLA_NET_0_116108, 
        HIEFFPLA_NET_0_116109, HIEFFPLA_NET_0_116110, 
        HIEFFPLA_NET_0_116111, HIEFFPLA_NET_0_116112, 
        HIEFFPLA_NET_0_116113, HIEFFPLA_NET_0_116114, 
        HIEFFPLA_NET_0_116115, HIEFFPLA_NET_0_116116, 
        HIEFFPLA_NET_0_116117, HIEFFPLA_NET_0_116118, 
        HIEFFPLA_NET_0_116119, HIEFFPLA_NET_0_116120, 
        HIEFFPLA_NET_0_116121, HIEFFPLA_NET_0_116122, 
        HIEFFPLA_NET_0_116123, HIEFFPLA_NET_0_116124, 
        HIEFFPLA_NET_0_116125, HIEFFPLA_NET_0_116126, 
        HIEFFPLA_NET_0_116127, HIEFFPLA_NET_0_116128, 
        HIEFFPLA_NET_0_116129, HIEFFPLA_NET_0_116130, 
        HIEFFPLA_NET_0_116131, HIEFFPLA_NET_0_116132, 
        HIEFFPLA_NET_0_116133, HIEFFPLA_NET_0_116134, 
        HIEFFPLA_NET_0_116135, HIEFFPLA_NET_0_116136, 
        HIEFFPLA_NET_0_116137, HIEFFPLA_NET_0_116138, 
        HIEFFPLA_NET_0_116139, HIEFFPLA_NET_0_116140, 
        HIEFFPLA_NET_0_116141, HIEFFPLA_NET_0_116142, 
        HIEFFPLA_NET_0_116143, HIEFFPLA_NET_0_116144, 
        HIEFFPLA_NET_0_116145, HIEFFPLA_NET_0_116146, 
        HIEFFPLA_NET_0_116147, HIEFFPLA_NET_0_116148, 
        HIEFFPLA_NET_0_116149, HIEFFPLA_NET_0_116150, 
        HIEFFPLA_NET_0_116151, HIEFFPLA_NET_0_116152, 
        HIEFFPLA_NET_0_116153, HIEFFPLA_NET_0_116154, 
        HIEFFPLA_NET_0_116155, HIEFFPLA_NET_0_116156, 
        HIEFFPLA_NET_0_116157, HIEFFPLA_NET_0_116158, 
        HIEFFPLA_NET_0_116159, HIEFFPLA_NET_0_116160, 
        HIEFFPLA_NET_0_116161, HIEFFPLA_NET_0_116162, 
        HIEFFPLA_NET_0_116163, HIEFFPLA_NET_0_116164, 
        HIEFFPLA_NET_0_116165, HIEFFPLA_NET_0_116166, 
        HIEFFPLA_NET_0_116167, HIEFFPLA_NET_0_116168, 
        HIEFFPLA_NET_0_116169, HIEFFPLA_NET_0_116170, 
        HIEFFPLA_NET_0_116171, HIEFFPLA_NET_0_116172, 
        HIEFFPLA_NET_0_116173, HIEFFPLA_NET_0_116174, 
        HIEFFPLA_NET_0_116175, HIEFFPLA_NET_0_116176, 
        HIEFFPLA_NET_0_116177, HIEFFPLA_NET_0_116178, 
        HIEFFPLA_NET_0_116179, HIEFFPLA_NET_0_116180, 
        HIEFFPLA_NET_0_116181, HIEFFPLA_NET_0_116182, 
        HIEFFPLA_NET_0_116183, HIEFFPLA_NET_0_116184, 
        HIEFFPLA_NET_0_116185, HIEFFPLA_NET_0_116186, 
        HIEFFPLA_NET_0_116187, HIEFFPLA_NET_0_116188, 
        HIEFFPLA_NET_0_116189, HIEFFPLA_NET_0_116190, 
        HIEFFPLA_NET_0_116191, HIEFFPLA_NET_0_116192, 
        HIEFFPLA_NET_0_116193, HIEFFPLA_NET_0_116194, 
        HIEFFPLA_NET_0_116195, HIEFFPLA_NET_0_116196, 
        HIEFFPLA_NET_0_116197, HIEFFPLA_NET_0_116198, 
        HIEFFPLA_NET_0_116199, HIEFFPLA_NET_0_116200, 
        HIEFFPLA_NET_0_116201, HIEFFPLA_NET_0_116202, 
        HIEFFPLA_NET_0_116203, HIEFFPLA_NET_0_116204, 
        HIEFFPLA_NET_0_116205, HIEFFPLA_NET_0_116206, 
        HIEFFPLA_NET_0_116207, HIEFFPLA_NET_0_116208, 
        HIEFFPLA_NET_0_116209, HIEFFPLA_NET_0_116210, 
        HIEFFPLA_NET_0_116211, HIEFFPLA_NET_0_116212, 
        HIEFFPLA_NET_0_116213, HIEFFPLA_NET_0_116214, 
        HIEFFPLA_NET_0_116215, HIEFFPLA_NET_0_116216, 
        HIEFFPLA_NET_0_116217, HIEFFPLA_NET_0_116218, 
        HIEFFPLA_NET_0_116219, HIEFFPLA_NET_0_116220, 
        HIEFFPLA_NET_0_116221, HIEFFPLA_NET_0_116222, 
        HIEFFPLA_NET_0_116223, HIEFFPLA_NET_0_116224, 
        HIEFFPLA_NET_0_116225, HIEFFPLA_NET_0_116226, 
        HIEFFPLA_NET_0_116227, HIEFFPLA_NET_0_116228, 
        HIEFFPLA_NET_0_116229, HIEFFPLA_NET_0_116230, 
        HIEFFPLA_NET_0_116231, HIEFFPLA_NET_0_116232, 
        HIEFFPLA_NET_0_116233, HIEFFPLA_NET_0_116234, 
        HIEFFPLA_NET_0_116235, HIEFFPLA_NET_0_116236, 
        HIEFFPLA_NET_0_116237, HIEFFPLA_NET_0_116238, 
        HIEFFPLA_NET_0_116239, HIEFFPLA_NET_0_116240, 
        HIEFFPLA_NET_0_116241, HIEFFPLA_NET_0_116242, 
        HIEFFPLA_NET_0_116243, HIEFFPLA_NET_0_116244, 
        HIEFFPLA_NET_0_116245, HIEFFPLA_NET_0_116246, 
        HIEFFPLA_NET_0_116247, HIEFFPLA_NET_0_116248, 
        HIEFFPLA_NET_0_116249, HIEFFPLA_NET_0_116250, 
        HIEFFPLA_NET_0_116251, HIEFFPLA_NET_0_116252, 
        HIEFFPLA_NET_0_116253, HIEFFPLA_NET_0_116254, 
        HIEFFPLA_NET_0_116255, HIEFFPLA_NET_0_116256, 
        HIEFFPLA_NET_0_116257, HIEFFPLA_NET_0_116258, 
        HIEFFPLA_NET_0_116259, HIEFFPLA_NET_0_116260, 
        HIEFFPLA_NET_0_116261, HIEFFPLA_NET_0_116262, 
        HIEFFPLA_NET_0_116263, HIEFFPLA_NET_0_116264, 
        HIEFFPLA_NET_0_116265, HIEFFPLA_NET_0_116266, 
        HIEFFPLA_NET_0_116267, HIEFFPLA_NET_0_116268, 
        HIEFFPLA_NET_0_116269, HIEFFPLA_NET_0_116270, 
        HIEFFPLA_NET_0_116271, HIEFFPLA_NET_0_116272, 
        HIEFFPLA_NET_0_116273, HIEFFPLA_NET_0_116274, 
        HIEFFPLA_NET_0_116275, HIEFFPLA_NET_0_116276, 
        HIEFFPLA_NET_0_116277, HIEFFPLA_NET_0_116278, 
        HIEFFPLA_NET_0_116279, HIEFFPLA_NET_0_116280, 
        HIEFFPLA_NET_0_116281, HIEFFPLA_NET_0_116282, 
        HIEFFPLA_NET_0_116283, HIEFFPLA_NET_0_116284, 
        HIEFFPLA_NET_0_116285, HIEFFPLA_NET_0_116286, 
        HIEFFPLA_NET_0_116287, HIEFFPLA_NET_0_116288, 
        HIEFFPLA_NET_0_116289, HIEFFPLA_NET_0_116290, 
        HIEFFPLA_NET_0_116291, HIEFFPLA_NET_0_116292, 
        HIEFFPLA_NET_0_116293, HIEFFPLA_NET_0_116294, 
        HIEFFPLA_NET_0_116295, HIEFFPLA_NET_0_116296, 
        HIEFFPLA_NET_0_116297, HIEFFPLA_NET_0_116298, 
        HIEFFPLA_NET_0_116299, HIEFFPLA_NET_0_116300, 
        HIEFFPLA_NET_0_116301, HIEFFPLA_NET_0_116302, 
        HIEFFPLA_NET_0_116303, HIEFFPLA_NET_0_116304, 
        HIEFFPLA_NET_0_116305, HIEFFPLA_NET_0_116306, 
        HIEFFPLA_NET_0_116307, HIEFFPLA_NET_0_116308, 
        HIEFFPLA_NET_0_116309, HIEFFPLA_NET_0_116310, 
        HIEFFPLA_NET_0_116311, HIEFFPLA_NET_0_116312, 
        HIEFFPLA_NET_0_116313, HIEFFPLA_NET_0_116314, 
        HIEFFPLA_NET_0_116315, HIEFFPLA_NET_0_116316, 
        HIEFFPLA_NET_0_116317, HIEFFPLA_NET_0_116318, 
        HIEFFPLA_NET_0_116319, HIEFFPLA_NET_0_116320, 
        HIEFFPLA_NET_0_116321, HIEFFPLA_NET_0_116322, 
        HIEFFPLA_NET_0_116323, HIEFFPLA_NET_0_116324, 
        HIEFFPLA_NET_0_116325, HIEFFPLA_NET_0_116326, 
        HIEFFPLA_NET_0_116327, HIEFFPLA_NET_0_116328, 
        HIEFFPLA_NET_0_116329, HIEFFPLA_NET_0_116330, 
        HIEFFPLA_NET_0_116331, HIEFFPLA_NET_0_116332, 
        HIEFFPLA_NET_0_116333, HIEFFPLA_NET_0_116334, 
        HIEFFPLA_NET_0_116335, HIEFFPLA_NET_0_116336, 
        HIEFFPLA_NET_0_116337, HIEFFPLA_NET_0_116338, 
        HIEFFPLA_NET_0_116339, HIEFFPLA_NET_0_116340, 
        HIEFFPLA_NET_0_116341, HIEFFPLA_NET_0_116342, 
        HIEFFPLA_NET_0_116343, HIEFFPLA_NET_0_116344, 
        HIEFFPLA_NET_0_116345, HIEFFPLA_NET_0_116346, 
        HIEFFPLA_NET_0_116347, HIEFFPLA_NET_0_116348, 
        HIEFFPLA_NET_0_116349, HIEFFPLA_NET_0_116350, 
        HIEFFPLA_NET_0_116351, HIEFFPLA_NET_0_116352, 
        HIEFFPLA_NET_0_116353, HIEFFPLA_NET_0_116354, 
        HIEFFPLA_NET_0_116355, HIEFFPLA_NET_0_116356, 
        HIEFFPLA_NET_0_116357, HIEFFPLA_NET_0_116358, 
        HIEFFPLA_NET_0_116359, HIEFFPLA_NET_0_116360, 
        HIEFFPLA_NET_0_116361, HIEFFPLA_NET_0_116362, 
        HIEFFPLA_NET_0_116363, HIEFFPLA_NET_0_116364, 
        HIEFFPLA_NET_0_116365, HIEFFPLA_NET_0_116366, 
        HIEFFPLA_NET_0_116367, HIEFFPLA_NET_0_116368, 
        HIEFFPLA_NET_0_116369, HIEFFPLA_NET_0_116370, 
        HIEFFPLA_NET_0_116371, HIEFFPLA_NET_0_116372, 
        HIEFFPLA_NET_0_116373, HIEFFPLA_NET_0_116374, 
        HIEFFPLA_NET_0_116375, HIEFFPLA_NET_0_116376, 
        HIEFFPLA_NET_0_116377, HIEFFPLA_NET_0_116378, 
        HIEFFPLA_NET_0_116379, HIEFFPLA_NET_0_116380, 
        HIEFFPLA_NET_0_116381, HIEFFPLA_NET_0_116382, 
        HIEFFPLA_NET_0_116383, HIEFFPLA_NET_0_116384, 
        HIEFFPLA_NET_0_116385, HIEFFPLA_NET_0_116386, 
        HIEFFPLA_NET_0_116387, HIEFFPLA_NET_0_116388, 
        HIEFFPLA_NET_0_116389, HIEFFPLA_NET_0_116390, 
        HIEFFPLA_NET_0_116391, HIEFFPLA_NET_0_116392, 
        HIEFFPLA_NET_0_116393, HIEFFPLA_NET_0_116394, 
        HIEFFPLA_NET_0_116395, HIEFFPLA_NET_0_116396, 
        HIEFFPLA_NET_0_116397, HIEFFPLA_NET_0_116398, 
        HIEFFPLA_NET_0_116399, HIEFFPLA_NET_0_116400, 
        HIEFFPLA_NET_0_116401, HIEFFPLA_NET_0_116402, 
        HIEFFPLA_NET_0_116403, HIEFFPLA_NET_0_116404, 
        HIEFFPLA_NET_0_116405, HIEFFPLA_NET_0_116406, 
        HIEFFPLA_NET_0_116407, HIEFFPLA_NET_0_116408, 
        HIEFFPLA_NET_0_116409, HIEFFPLA_NET_0_116410, 
        HIEFFPLA_NET_0_116411, HIEFFPLA_NET_0_116412, 
        HIEFFPLA_NET_0_116413, HIEFFPLA_NET_0_116414, 
        HIEFFPLA_NET_0_116415, HIEFFPLA_NET_0_116416, 
        HIEFFPLA_NET_0_116417, HIEFFPLA_NET_0_116418, 
        HIEFFPLA_NET_0_116419, HIEFFPLA_NET_0_116420, 
        HIEFFPLA_NET_0_116421, HIEFFPLA_NET_0_116422, 
        HIEFFPLA_NET_0_116423, HIEFFPLA_NET_0_116424, 
        HIEFFPLA_NET_0_116425, HIEFFPLA_NET_0_116426, 
        HIEFFPLA_NET_0_116427, HIEFFPLA_NET_0_116428, 
        HIEFFPLA_NET_0_116429, HIEFFPLA_NET_0_116430, 
        HIEFFPLA_NET_0_116431, HIEFFPLA_NET_0_116432, 
        HIEFFPLA_NET_0_116433, HIEFFPLA_NET_0_116434, 
        HIEFFPLA_NET_0_116435, HIEFFPLA_NET_0_116436, 
        HIEFFPLA_NET_0_116437, HIEFFPLA_NET_0_116438, 
        HIEFFPLA_NET_0_116439, HIEFFPLA_NET_0_116440, 
        HIEFFPLA_NET_0_116441, HIEFFPLA_NET_0_116442, 
        HIEFFPLA_NET_0_116443, HIEFFPLA_NET_0_116444, 
        HIEFFPLA_NET_0_116445, HIEFFPLA_NET_0_116446, 
        HIEFFPLA_NET_0_116447, HIEFFPLA_NET_0_116448, 
        HIEFFPLA_NET_0_116449, HIEFFPLA_NET_0_116450, 
        HIEFFPLA_NET_0_116451, HIEFFPLA_NET_0_116452, 
        HIEFFPLA_NET_0_116453, HIEFFPLA_NET_0_116454, 
        HIEFFPLA_NET_0_116455, HIEFFPLA_NET_0_116456, 
        HIEFFPLA_NET_0_116457, HIEFFPLA_NET_0_116458, 
        HIEFFPLA_NET_0_116459, HIEFFPLA_NET_0_116460, 
        HIEFFPLA_NET_0_116461, HIEFFPLA_NET_0_116462, 
        HIEFFPLA_NET_0_116463, HIEFFPLA_NET_0_116464, 
        HIEFFPLA_NET_0_116465, HIEFFPLA_NET_0_116466, 
        HIEFFPLA_NET_0_116467, HIEFFPLA_NET_0_116468, 
        HIEFFPLA_NET_0_116469, HIEFFPLA_NET_0_116470, 
        HIEFFPLA_NET_0_116471, HIEFFPLA_NET_0_116472, 
        HIEFFPLA_NET_0_116473, HIEFFPLA_NET_0_116474, 
        HIEFFPLA_NET_0_116475, HIEFFPLA_NET_0_116476, 
        HIEFFPLA_NET_0_116477, HIEFFPLA_NET_0_116478, 
        HIEFFPLA_NET_0_116479, HIEFFPLA_NET_0_116480, 
        HIEFFPLA_NET_0_116481, HIEFFPLA_NET_0_116482, 
        HIEFFPLA_NET_0_116483, HIEFFPLA_NET_0_116484, 
        HIEFFPLA_NET_0_116485, HIEFFPLA_NET_0_116486, 
        HIEFFPLA_NET_0_116487, HIEFFPLA_NET_0_116488, 
        HIEFFPLA_NET_0_116489, HIEFFPLA_NET_0_116490, 
        HIEFFPLA_NET_0_116491, HIEFFPLA_NET_0_116492, 
        HIEFFPLA_NET_0_116493, HIEFFPLA_NET_0_116494, 
        HIEFFPLA_NET_0_116495, HIEFFPLA_NET_0_116496, 
        HIEFFPLA_NET_0_116497, HIEFFPLA_NET_0_116498, 
        HIEFFPLA_NET_0_116499, HIEFFPLA_NET_0_116500, 
        HIEFFPLA_NET_0_116501, HIEFFPLA_NET_0_116502, 
        HIEFFPLA_NET_0_116503, HIEFFPLA_NET_0_116504, 
        HIEFFPLA_NET_0_116505, HIEFFPLA_NET_0_116506, 
        HIEFFPLA_NET_0_116507, HIEFFPLA_NET_0_116508, 
        HIEFFPLA_NET_0_116509, HIEFFPLA_NET_0_116510, 
        HIEFFPLA_NET_0_116511, HIEFFPLA_NET_0_116512, 
        HIEFFPLA_NET_0_116513, HIEFFPLA_NET_0_116514, 
        HIEFFPLA_NET_0_116515, HIEFFPLA_NET_0_116516, 
        HIEFFPLA_NET_0_116517, HIEFFPLA_NET_0_116518, 
        HIEFFPLA_NET_0_116519, HIEFFPLA_NET_0_116520, 
        HIEFFPLA_NET_0_116521, HIEFFPLA_NET_0_116522, 
        HIEFFPLA_NET_0_116523, HIEFFPLA_NET_0_116524, 
        HIEFFPLA_NET_0_116525, HIEFFPLA_NET_0_116526, 
        HIEFFPLA_NET_0_116527, HIEFFPLA_NET_0_116528, 
        HIEFFPLA_NET_0_116529, HIEFFPLA_NET_0_116530, 
        HIEFFPLA_NET_0_116531, HIEFFPLA_NET_0_116532, 
        HIEFFPLA_NET_0_116533, HIEFFPLA_NET_0_116534, 
        HIEFFPLA_NET_0_116535, HIEFFPLA_NET_0_116536, 
        HIEFFPLA_NET_0_116537, HIEFFPLA_NET_0_116538, 
        HIEFFPLA_NET_0_116539, HIEFFPLA_NET_0_116540, 
        HIEFFPLA_NET_0_116541, HIEFFPLA_NET_0_116542, 
        HIEFFPLA_NET_0_116543, HIEFFPLA_NET_0_116544, 
        HIEFFPLA_NET_0_116545, HIEFFPLA_NET_0_116546, 
        HIEFFPLA_NET_0_116547, HIEFFPLA_NET_0_116548, 
        HIEFFPLA_NET_0_116549, HIEFFPLA_NET_0_116550, 
        HIEFFPLA_NET_0_116551, HIEFFPLA_NET_0_116552, 
        HIEFFPLA_NET_0_116553, HIEFFPLA_NET_0_116554, 
        HIEFFPLA_NET_0_116555, HIEFFPLA_NET_0_116556, 
        HIEFFPLA_NET_0_116557, HIEFFPLA_NET_0_116558, 
        HIEFFPLA_NET_0_116559, HIEFFPLA_NET_0_116560, 
        HIEFFPLA_NET_0_116561, HIEFFPLA_NET_0_116562, 
        HIEFFPLA_NET_0_116563, HIEFFPLA_NET_0_116564, 
        HIEFFPLA_NET_0_116565, HIEFFPLA_NET_0_116566, 
        HIEFFPLA_NET_0_116567, HIEFFPLA_NET_0_116568, 
        HIEFFPLA_NET_0_116569, HIEFFPLA_NET_0_116570, 
        HIEFFPLA_NET_0_116571, HIEFFPLA_NET_0_116572, 
        HIEFFPLA_NET_0_116573, HIEFFPLA_NET_0_116574, 
        HIEFFPLA_NET_0_116575, HIEFFPLA_NET_0_116576, 
        HIEFFPLA_NET_0_116577, HIEFFPLA_NET_0_116578, 
        HIEFFPLA_NET_0_116579, HIEFFPLA_NET_0_116580, 
        HIEFFPLA_NET_0_116581, HIEFFPLA_NET_0_116582, 
        HIEFFPLA_NET_0_116583, HIEFFPLA_NET_0_116584, 
        HIEFFPLA_NET_0_116585, HIEFFPLA_NET_0_116586, 
        HIEFFPLA_NET_0_116587, HIEFFPLA_NET_0_116588, 
        HIEFFPLA_NET_0_116589, HIEFFPLA_NET_0_116590, 
        HIEFFPLA_NET_0_116591, HIEFFPLA_NET_0_116592, 
        HIEFFPLA_NET_0_116593, HIEFFPLA_NET_0_116594, 
        HIEFFPLA_NET_0_116595, HIEFFPLA_NET_0_116596, 
        HIEFFPLA_NET_0_116597, HIEFFPLA_NET_0_116598, 
        HIEFFPLA_NET_0_116599, HIEFFPLA_NET_0_116600, 
        HIEFFPLA_NET_0_116601, HIEFFPLA_NET_0_116602, 
        HIEFFPLA_NET_0_116603, HIEFFPLA_NET_0_116604, 
        HIEFFPLA_NET_0_116605, HIEFFPLA_NET_0_116606, 
        HIEFFPLA_NET_0_116607, HIEFFPLA_NET_0_116608, 
        HIEFFPLA_NET_0_116609, HIEFFPLA_NET_0_116610, 
        HIEFFPLA_NET_0_116611, HIEFFPLA_NET_0_116612, 
        HIEFFPLA_NET_0_116613, HIEFFPLA_NET_0_116614, 
        HIEFFPLA_NET_0_116615, HIEFFPLA_NET_0_116616, 
        HIEFFPLA_NET_0_116617, HIEFFPLA_NET_0_116618, 
        HIEFFPLA_NET_0_116619, HIEFFPLA_NET_0_116620, 
        HIEFFPLA_NET_0_116621, HIEFFPLA_NET_0_116622, 
        HIEFFPLA_NET_0_116623, HIEFFPLA_NET_0_116624, 
        HIEFFPLA_NET_0_116625, HIEFFPLA_NET_0_116626, 
        HIEFFPLA_NET_0_116627, HIEFFPLA_NET_0_116628, 
        HIEFFPLA_NET_0_116629, HIEFFPLA_NET_0_116630, 
        HIEFFPLA_NET_0_116631, HIEFFPLA_NET_0_116632, 
        HIEFFPLA_NET_0_116633, HIEFFPLA_NET_0_116634, 
        HIEFFPLA_NET_0_116635, HIEFFPLA_NET_0_116636, 
        HIEFFPLA_NET_0_116637, HIEFFPLA_NET_0_116638, 
        HIEFFPLA_NET_0_116639, HIEFFPLA_NET_0_116640, 
        HIEFFPLA_NET_0_116641, HIEFFPLA_NET_0_116642, 
        HIEFFPLA_NET_0_116643, HIEFFPLA_NET_0_116644, 
        HIEFFPLA_NET_0_116645, HIEFFPLA_NET_0_116646, 
        HIEFFPLA_NET_0_116647, HIEFFPLA_NET_0_116648, 
        HIEFFPLA_NET_0_116649, HIEFFPLA_NET_0_116650, 
        HIEFFPLA_NET_0_116651, HIEFFPLA_NET_0_116652, 
        HIEFFPLA_NET_0_116653, HIEFFPLA_NET_0_116654, 
        HIEFFPLA_NET_0_116655, HIEFFPLA_NET_0_116656, 
        HIEFFPLA_NET_0_116657, HIEFFPLA_NET_0_116658, 
        HIEFFPLA_NET_0_116659, HIEFFPLA_NET_0_116660, 
        HIEFFPLA_NET_0_116661, HIEFFPLA_NET_0_116662, 
        HIEFFPLA_NET_0_116663, HIEFFPLA_NET_0_116664, 
        HIEFFPLA_NET_0_116665, HIEFFPLA_NET_0_116666, 
        HIEFFPLA_NET_0_116667, HIEFFPLA_NET_0_116668, 
        HIEFFPLA_NET_0_116669, HIEFFPLA_NET_0_116670, 
        HIEFFPLA_NET_0_116671, HIEFFPLA_NET_0_116672, 
        HIEFFPLA_NET_0_116673, HIEFFPLA_NET_0_116674, 
        HIEFFPLA_NET_0_116675, HIEFFPLA_NET_0_116676, 
        HIEFFPLA_NET_0_116677, HIEFFPLA_NET_0_116678, 
        HIEFFPLA_NET_0_116679, HIEFFPLA_NET_0_116680, 
        HIEFFPLA_NET_0_116681, HIEFFPLA_NET_0_116682, 
        HIEFFPLA_NET_0_116683, HIEFFPLA_NET_0_116684, 
        HIEFFPLA_NET_0_116685, HIEFFPLA_NET_0_116686, 
        HIEFFPLA_NET_0_116687, HIEFFPLA_NET_0_116688, 
        HIEFFPLA_NET_0_116689, HIEFFPLA_NET_0_116690, 
        HIEFFPLA_NET_0_116691, HIEFFPLA_NET_0_116692, 
        HIEFFPLA_NET_0_116693, HIEFFPLA_NET_0_116694, 
        HIEFFPLA_NET_0_116695, HIEFFPLA_NET_0_116696, 
        HIEFFPLA_NET_0_116697, HIEFFPLA_NET_0_116698, 
        HIEFFPLA_NET_0_116699, HIEFFPLA_NET_0_116700, 
        HIEFFPLA_NET_0_116701, HIEFFPLA_NET_0_116702, 
        HIEFFPLA_NET_0_116703, HIEFFPLA_NET_0_116704, 
        HIEFFPLA_NET_0_116705, HIEFFPLA_NET_0_116706, 
        HIEFFPLA_NET_0_116707, HIEFFPLA_NET_0_116708, 
        HIEFFPLA_NET_0_116709, HIEFFPLA_NET_0_116710, 
        HIEFFPLA_NET_0_116711, HIEFFPLA_NET_0_116712, 
        HIEFFPLA_NET_0_116713, HIEFFPLA_NET_0_116714, 
        HIEFFPLA_NET_0_116715, HIEFFPLA_NET_0_116716, 
        HIEFFPLA_NET_0_116717, HIEFFPLA_NET_0_116718, 
        HIEFFPLA_NET_0_116719, HIEFFPLA_NET_0_116720, 
        HIEFFPLA_NET_0_116721, HIEFFPLA_NET_0_116722, 
        HIEFFPLA_NET_0_116723, HIEFFPLA_NET_0_116724, 
        HIEFFPLA_NET_0_116725, HIEFFPLA_NET_0_116726, 
        HIEFFPLA_NET_0_116727, HIEFFPLA_NET_0_116728, 
        HIEFFPLA_NET_0_116729, HIEFFPLA_NET_0_116730, 
        HIEFFPLA_NET_0_116731, HIEFFPLA_NET_0_116732, 
        HIEFFPLA_NET_0_116733, HIEFFPLA_NET_0_116734, 
        HIEFFPLA_NET_0_116735, HIEFFPLA_NET_0_116736, 
        HIEFFPLA_NET_0_116737, HIEFFPLA_NET_0_116738, 
        HIEFFPLA_NET_0_116739, HIEFFPLA_NET_0_116740, 
        HIEFFPLA_NET_0_116741, HIEFFPLA_NET_0_116742, 
        HIEFFPLA_NET_0_116743, HIEFFPLA_NET_0_116744, 
        HIEFFPLA_NET_0_116745, HIEFFPLA_NET_0_116746, 
        HIEFFPLA_NET_0_116747, HIEFFPLA_NET_0_116748, 
        HIEFFPLA_NET_0_116749, HIEFFPLA_NET_0_116750, 
        HIEFFPLA_NET_0_116751, HIEFFPLA_NET_0_116752, 
        HIEFFPLA_NET_0_116753, HIEFFPLA_NET_0_116754, 
        HIEFFPLA_NET_0_116755, HIEFFPLA_NET_0_116756, 
        HIEFFPLA_NET_0_116757, HIEFFPLA_NET_0_116758, 
        HIEFFPLA_NET_0_116759, HIEFFPLA_NET_0_116760, 
        HIEFFPLA_NET_0_116761, HIEFFPLA_NET_0_116762, 
        HIEFFPLA_NET_0_116763, HIEFFPLA_NET_0_116764, 
        HIEFFPLA_NET_0_116765, HIEFFPLA_NET_0_116766, 
        HIEFFPLA_NET_0_116767, HIEFFPLA_NET_0_116768, 
        HIEFFPLA_NET_0_116769, HIEFFPLA_NET_0_116770, 
        HIEFFPLA_NET_0_116771, HIEFFPLA_NET_0_116772, 
        HIEFFPLA_NET_0_116773, HIEFFPLA_NET_0_116774, 
        HIEFFPLA_NET_0_116775, HIEFFPLA_NET_0_116776, 
        HIEFFPLA_NET_0_116777, HIEFFPLA_NET_0_116778, 
        HIEFFPLA_NET_0_116779, HIEFFPLA_NET_0_116780, 
        HIEFFPLA_NET_0_116781, HIEFFPLA_NET_0_116782, 
        HIEFFPLA_NET_0_116783, HIEFFPLA_NET_0_116784, 
        HIEFFPLA_NET_0_116785, HIEFFPLA_NET_0_116786, 
        HIEFFPLA_NET_0_116787, HIEFFPLA_NET_0_116788, 
        HIEFFPLA_NET_0_116789, HIEFFPLA_NET_0_116790, 
        HIEFFPLA_NET_0_116791, HIEFFPLA_NET_0_116792, 
        HIEFFPLA_NET_0_116793, HIEFFPLA_NET_0_116794, 
        HIEFFPLA_NET_0_116795, HIEFFPLA_NET_0_116796, 
        HIEFFPLA_NET_0_116797, HIEFFPLA_NET_0_116798, 
        HIEFFPLA_NET_0_116799, HIEFFPLA_NET_0_116800, 
        HIEFFPLA_NET_0_116801, HIEFFPLA_NET_0_116802, 
        HIEFFPLA_NET_0_116803, HIEFFPLA_NET_0_116804, 
        HIEFFPLA_NET_0_116805, HIEFFPLA_NET_0_116806, 
        HIEFFPLA_NET_0_116807, HIEFFPLA_NET_0_116808, 
        HIEFFPLA_NET_0_116809, HIEFFPLA_NET_0_116810, 
        HIEFFPLA_NET_0_116811, HIEFFPLA_NET_0_116812, 
        HIEFFPLA_NET_0_116813, HIEFFPLA_NET_0_116814, 
        HIEFFPLA_NET_0_116815, HIEFFPLA_NET_0_116816, 
        HIEFFPLA_NET_0_116817, HIEFFPLA_NET_0_116818, 
        HIEFFPLA_NET_0_116819, HIEFFPLA_NET_0_116820, 
        HIEFFPLA_NET_0_116821, HIEFFPLA_NET_0_116822, 
        HIEFFPLA_NET_0_116823, HIEFFPLA_NET_0_116824, 
        HIEFFPLA_NET_0_116825, HIEFFPLA_NET_0_116826, 
        HIEFFPLA_NET_0_116827, HIEFFPLA_NET_0_116828, 
        HIEFFPLA_NET_0_116829, HIEFFPLA_NET_0_116830, 
        HIEFFPLA_NET_0_116831, HIEFFPLA_NET_0_116832, 
        HIEFFPLA_NET_0_116833, HIEFFPLA_NET_0_116834, 
        HIEFFPLA_NET_0_116835, HIEFFPLA_NET_0_116836, 
        HIEFFPLA_NET_0_116837, HIEFFPLA_NET_0_116838, 
        HIEFFPLA_NET_0_116839, HIEFFPLA_NET_0_116840, 
        HIEFFPLA_NET_0_116841, HIEFFPLA_NET_0_116842, 
        HIEFFPLA_NET_0_116843, HIEFFPLA_NET_0_116844, 
        HIEFFPLA_NET_0_116845, HIEFFPLA_NET_0_116846, 
        HIEFFPLA_NET_0_116847, HIEFFPLA_NET_0_116848, 
        HIEFFPLA_NET_0_116849, HIEFFPLA_NET_0_116850, 
        HIEFFPLA_NET_0_116851, HIEFFPLA_NET_0_116852, 
        HIEFFPLA_NET_0_116853, HIEFFPLA_NET_0_116854, 
        HIEFFPLA_NET_0_116855, HIEFFPLA_NET_0_116856, 
        HIEFFPLA_NET_0_116857, HIEFFPLA_NET_0_116858, 
        HIEFFPLA_NET_0_116859, HIEFFPLA_NET_0_116860, 
        HIEFFPLA_NET_0_116861, HIEFFPLA_NET_0_116862, 
        HIEFFPLA_NET_0_116863, HIEFFPLA_NET_0_116864, 
        HIEFFPLA_NET_0_116865, HIEFFPLA_NET_0_116866, 
        HIEFFPLA_NET_0_116867, HIEFFPLA_NET_0_116868, 
        HIEFFPLA_NET_0_116869, HIEFFPLA_NET_0_116870, 
        HIEFFPLA_NET_0_116871, HIEFFPLA_NET_0_116872, 
        HIEFFPLA_NET_0_116873, HIEFFPLA_NET_0_116874, 
        HIEFFPLA_NET_0_116875, HIEFFPLA_NET_0_116876, 
        HIEFFPLA_NET_0_116877, HIEFFPLA_NET_0_116878, 
        HIEFFPLA_NET_0_116879, HIEFFPLA_NET_0_116880, 
        HIEFFPLA_NET_0_116881, HIEFFPLA_NET_0_116882, 
        HIEFFPLA_NET_0_116883, HIEFFPLA_NET_0_116884, 
        HIEFFPLA_NET_0_116885, HIEFFPLA_NET_0_116886, 
        HIEFFPLA_NET_0_116887, HIEFFPLA_NET_0_116888, 
        HIEFFPLA_NET_0_116889, HIEFFPLA_NET_0_116890, 
        HIEFFPLA_NET_0_116891, HIEFFPLA_NET_0_116892, 
        HIEFFPLA_NET_0_116893, HIEFFPLA_NET_0_116894, 
        HIEFFPLA_NET_0_116895, HIEFFPLA_NET_0_116896, 
        HIEFFPLA_NET_0_116897, HIEFFPLA_NET_0_116898, 
        HIEFFPLA_NET_0_116899, HIEFFPLA_NET_0_116900, 
        HIEFFPLA_NET_0_116901, HIEFFPLA_NET_0_116902, 
        HIEFFPLA_NET_0_116903, HIEFFPLA_NET_0_116904, 
        HIEFFPLA_NET_0_116905, HIEFFPLA_NET_0_116906, 
        HIEFFPLA_NET_0_116907, HIEFFPLA_NET_0_116924, 
        HIEFFPLA_NET_0_116925, HIEFFPLA_NET_0_116926, 
        HIEFFPLA_NET_0_116927, HIEFFPLA_NET_0_116928, 
        HIEFFPLA_NET_0_116929, HIEFFPLA_NET_0_116930, 
        HIEFFPLA_NET_0_116931, HIEFFPLA_NET_0_116932, 
        HIEFFPLA_NET_0_116933, HIEFFPLA_NET_0_116934, 
        HIEFFPLA_NET_0_116935, HIEFFPLA_NET_0_116936, 
        HIEFFPLA_NET_0_116937, HIEFFPLA_NET_0_116938, 
        HIEFFPLA_NET_0_116939, HIEFFPLA_NET_0_116940, 
        HIEFFPLA_NET_0_116941, HIEFFPLA_NET_0_116942, 
        HIEFFPLA_NET_0_116943, HIEFFPLA_NET_0_116944, 
        HIEFFPLA_NET_0_116945, HIEFFPLA_NET_0_116946, 
        HIEFFPLA_NET_0_116947, HIEFFPLA_NET_0_116948, 
        HIEFFPLA_NET_0_116949, HIEFFPLA_NET_0_116950, 
        HIEFFPLA_NET_0_116951, HIEFFPLA_NET_0_116952, 
        HIEFFPLA_NET_0_116953, HIEFFPLA_NET_0_116954, 
        HIEFFPLA_NET_0_116955, HIEFFPLA_NET_0_116956, 
        HIEFFPLA_NET_0_116957, HIEFFPLA_NET_0_116958, 
        HIEFFPLA_NET_0_116959, HIEFFPLA_NET_0_116960, 
        HIEFFPLA_NET_0_116961, HIEFFPLA_NET_0_116962, 
        HIEFFPLA_NET_0_116963, HIEFFPLA_NET_0_116964, 
        HIEFFPLA_NET_0_116965, HIEFFPLA_NET_0_116966, 
        HIEFFPLA_NET_0_116967, HIEFFPLA_NET_0_116968, 
        HIEFFPLA_NET_0_116969, HIEFFPLA_NET_0_116970, 
        HIEFFPLA_NET_0_116971, HIEFFPLA_NET_0_116972, 
        HIEFFPLA_NET_0_116973, HIEFFPLA_NET_0_116974, 
        HIEFFPLA_NET_0_116975, HIEFFPLA_NET_0_116976, 
        HIEFFPLA_NET_0_116977, HIEFFPLA_NET_0_116978, 
        HIEFFPLA_NET_0_116979, HIEFFPLA_NET_0_116980, 
        HIEFFPLA_NET_0_116981, HIEFFPLA_NET_0_116982, 
        HIEFFPLA_NET_0_116983, HIEFFPLA_NET_0_116984, 
        HIEFFPLA_NET_0_116985, HIEFFPLA_NET_0_116986, 
        HIEFFPLA_NET_0_116987, HIEFFPLA_NET_0_116988, 
        HIEFFPLA_NET_0_116989, HIEFFPLA_NET_0_116990, 
        HIEFFPLA_NET_0_116991, HIEFFPLA_NET_0_116992, 
        HIEFFPLA_NET_0_116993, HIEFFPLA_NET_0_116994, 
        HIEFFPLA_NET_0_116995, HIEFFPLA_NET_0_116996, 
        HIEFFPLA_NET_0_116997, HIEFFPLA_NET_0_116998, 
        HIEFFPLA_NET_0_116999, HIEFFPLA_NET_0_117000, 
        HIEFFPLA_NET_0_117001, HIEFFPLA_NET_0_117002, 
        HIEFFPLA_NET_0_117003, HIEFFPLA_NET_0_117004, 
        HIEFFPLA_NET_0_117005, HIEFFPLA_NET_0_117006, 
        HIEFFPLA_NET_0_117007, HIEFFPLA_NET_0_117008, 
        HIEFFPLA_NET_0_117009, HIEFFPLA_NET_0_117010, 
        HIEFFPLA_NET_0_117011, HIEFFPLA_NET_0_117012, 
        HIEFFPLA_NET_0_117013, HIEFFPLA_NET_0_117014, 
        HIEFFPLA_NET_0_117015, HIEFFPLA_NET_0_117016, 
        HIEFFPLA_NET_0_117017, HIEFFPLA_NET_0_117018, 
        HIEFFPLA_NET_0_117019, HIEFFPLA_NET_0_117020, 
        HIEFFPLA_NET_0_117021, HIEFFPLA_NET_0_117022, 
        HIEFFPLA_NET_0_117023, HIEFFPLA_NET_0_117024, 
        HIEFFPLA_NET_0_117025, HIEFFPLA_NET_0_117026, 
        HIEFFPLA_NET_0_117027, HIEFFPLA_NET_0_117028, 
        HIEFFPLA_NET_0_117029, HIEFFPLA_NET_0_117030, 
        HIEFFPLA_NET_0_117031, HIEFFPLA_NET_0_117032, 
        HIEFFPLA_NET_0_117033, HIEFFPLA_NET_0_117034, 
        HIEFFPLA_NET_0_117035, HIEFFPLA_NET_0_117036, 
        HIEFFPLA_NET_0_117037, HIEFFPLA_NET_0_117038, 
        HIEFFPLA_NET_0_117039, HIEFFPLA_NET_0_117040, 
        HIEFFPLA_NET_0_117041, HIEFFPLA_NET_0_117042, 
        HIEFFPLA_NET_0_117043, HIEFFPLA_NET_0_117044, 
        HIEFFPLA_NET_0_117045, HIEFFPLA_NET_0_117046, 
        HIEFFPLA_NET_0_117047, HIEFFPLA_NET_0_117048, 
        HIEFFPLA_NET_0_117049, HIEFFPLA_NET_0_117050, 
        HIEFFPLA_NET_0_117051, HIEFFPLA_NET_0_117052, 
        HIEFFPLA_NET_0_117053, HIEFFPLA_NET_0_117054, 
        HIEFFPLA_NET_0_117055, HIEFFPLA_NET_0_117056, 
        HIEFFPLA_NET_0_117057, HIEFFPLA_NET_0_117058, 
        HIEFFPLA_NET_0_117059, HIEFFPLA_NET_0_117060, 
        HIEFFPLA_NET_0_117061, HIEFFPLA_NET_0_117062, 
        HIEFFPLA_NET_0_117063, HIEFFPLA_NET_0_117064, 
        HIEFFPLA_NET_0_117065, HIEFFPLA_NET_0_117066, 
        HIEFFPLA_NET_0_117067, HIEFFPLA_NET_0_117068, 
        HIEFFPLA_NET_0_117069, HIEFFPLA_NET_0_117070, 
        HIEFFPLA_NET_0_117071, HIEFFPLA_NET_0_117072, 
        HIEFFPLA_NET_0_117073, HIEFFPLA_NET_0_117074, 
        HIEFFPLA_NET_0_117075, HIEFFPLA_NET_0_117076, 
        HIEFFPLA_NET_0_117077, HIEFFPLA_NET_0_117078, 
        HIEFFPLA_NET_0_117079, HIEFFPLA_NET_0_117080, 
        HIEFFPLA_NET_0_117081, HIEFFPLA_NET_0_117082, 
        HIEFFPLA_NET_0_117083, HIEFFPLA_NET_0_117084, 
        HIEFFPLA_NET_0_117085, HIEFFPLA_NET_0_117086, 
        HIEFFPLA_NET_0_117087, HIEFFPLA_NET_0_117088, 
        HIEFFPLA_NET_0_117089, HIEFFPLA_NET_0_117090, 
        HIEFFPLA_NET_0_117091, HIEFFPLA_NET_0_117092, 
        HIEFFPLA_NET_0_117093, HIEFFPLA_NET_0_117094, 
        HIEFFPLA_NET_0_117095, HIEFFPLA_NET_0_117096, 
        HIEFFPLA_NET_0_117097, HIEFFPLA_NET_0_117098, 
        HIEFFPLA_NET_0_117099, HIEFFPLA_NET_0_117100, 
        HIEFFPLA_NET_0_117101, HIEFFPLA_NET_0_117102, 
        HIEFFPLA_NET_0_117103, HIEFFPLA_NET_0_117104, 
        HIEFFPLA_NET_0_117105, HIEFFPLA_NET_0_117106, 
        HIEFFPLA_NET_0_117107, HIEFFPLA_NET_0_117108, 
        HIEFFPLA_NET_0_117109, HIEFFPLA_NET_0_117110, 
        HIEFFPLA_NET_0_117111, HIEFFPLA_NET_0_117112, 
        HIEFFPLA_NET_0_117113, HIEFFPLA_NET_0_117114, 
        HIEFFPLA_NET_0_117115, HIEFFPLA_NET_0_117116, 
        HIEFFPLA_NET_0_117117, HIEFFPLA_NET_0_117118, 
        HIEFFPLA_NET_0_117119, HIEFFPLA_NET_0_117120, 
        HIEFFPLA_NET_0_117121, HIEFFPLA_NET_0_117122, 
        HIEFFPLA_NET_0_117123, HIEFFPLA_NET_0_117124, 
        HIEFFPLA_NET_0_117125, HIEFFPLA_NET_0_117126, 
        HIEFFPLA_NET_0_117127, HIEFFPLA_NET_0_117128, 
        HIEFFPLA_NET_0_117129, HIEFFPLA_NET_0_117130, 
        HIEFFPLA_NET_0_117131, HIEFFPLA_NET_0_117132, 
        HIEFFPLA_NET_0_117133, HIEFFPLA_NET_0_117134, 
        HIEFFPLA_NET_0_117135, HIEFFPLA_NET_0_117136, 
        HIEFFPLA_NET_0_117137, HIEFFPLA_NET_0_117138, 
        HIEFFPLA_NET_0_117139, HIEFFPLA_NET_0_117140, 
        HIEFFPLA_NET_0_117141, HIEFFPLA_NET_0_117142, 
        HIEFFPLA_NET_0_117143, HIEFFPLA_NET_0_117144, 
        HIEFFPLA_NET_0_117145, HIEFFPLA_NET_0_117146, 
        HIEFFPLA_NET_0_117147, HIEFFPLA_NET_0_117148, 
        HIEFFPLA_NET_0_117149, HIEFFPLA_NET_0_117150, 
        HIEFFPLA_NET_0_117151, HIEFFPLA_NET_0_117152, 
        HIEFFPLA_NET_0_117153, HIEFFPLA_NET_0_117154, 
        HIEFFPLA_NET_0_117155, HIEFFPLA_NET_0_117156, 
        HIEFFPLA_NET_0_117157, HIEFFPLA_NET_0_117158, 
        HIEFFPLA_NET_0_117159, HIEFFPLA_NET_0_117160, 
        HIEFFPLA_NET_0_117161, HIEFFPLA_NET_0_117162, 
        HIEFFPLA_NET_0_117163, HIEFFPLA_NET_0_117164, 
        HIEFFPLA_NET_0_117165, HIEFFPLA_NET_0_117166, 
        HIEFFPLA_NET_0_117167, HIEFFPLA_NET_0_117168, 
        HIEFFPLA_NET_0_117169, HIEFFPLA_NET_0_117170, 
        HIEFFPLA_NET_0_117171, HIEFFPLA_NET_0_117172, 
        HIEFFPLA_NET_0_117173, HIEFFPLA_NET_0_117174, 
        HIEFFPLA_NET_0_117175, HIEFFPLA_NET_0_117176, 
        HIEFFPLA_NET_0_117177, HIEFFPLA_NET_0_117178, 
        HIEFFPLA_NET_0_117179, HIEFFPLA_NET_0_117180, 
        HIEFFPLA_NET_0_117181, HIEFFPLA_NET_0_117182, 
        HIEFFPLA_NET_0_117183, HIEFFPLA_NET_0_117184, 
        HIEFFPLA_NET_0_117185, HIEFFPLA_NET_0_117186, 
        HIEFFPLA_NET_0_117187, HIEFFPLA_NET_0_117188, 
        HIEFFPLA_NET_0_117189, HIEFFPLA_NET_0_117190, 
        HIEFFPLA_NET_0_117191, HIEFFPLA_NET_0_117192, 
        HIEFFPLA_NET_0_117193, HIEFFPLA_NET_0_117194, 
        HIEFFPLA_NET_0_117195, HIEFFPLA_NET_0_117196, 
        HIEFFPLA_NET_0_117197, HIEFFPLA_NET_0_117198, 
        HIEFFPLA_NET_0_117199, HIEFFPLA_NET_0_117200, 
        HIEFFPLA_NET_0_117201, HIEFFPLA_NET_0_117202, 
        HIEFFPLA_NET_0_117203, HIEFFPLA_NET_0_117204, 
        HIEFFPLA_NET_0_117205, HIEFFPLA_NET_0_117206, 
        HIEFFPLA_NET_0_117207, HIEFFPLA_NET_0_117208, 
        HIEFFPLA_NET_0_117209, HIEFFPLA_NET_0_117210, 
        HIEFFPLA_NET_0_117211, HIEFFPLA_NET_0_117212, 
        HIEFFPLA_NET_0_117213, HIEFFPLA_NET_0_117214, 
        HIEFFPLA_NET_0_117215, HIEFFPLA_NET_0_117216, 
        HIEFFPLA_NET_0_117217, HIEFFPLA_NET_0_117218, 
        HIEFFPLA_NET_0_117219, HIEFFPLA_NET_0_117220, 
        HIEFFPLA_NET_0_117221, HIEFFPLA_NET_0_117222, 
        HIEFFPLA_NET_0_117223, HIEFFPLA_NET_0_117224, 
        HIEFFPLA_NET_0_117225, HIEFFPLA_NET_0_117226, 
        HIEFFPLA_NET_0_117227, HIEFFPLA_NET_0_117228, 
        HIEFFPLA_NET_0_117229, HIEFFPLA_NET_0_117230, 
        HIEFFPLA_NET_0_117231, HIEFFPLA_NET_0_117232, 
        HIEFFPLA_NET_0_117233, HIEFFPLA_NET_0_117234, 
        HIEFFPLA_NET_0_117235, HIEFFPLA_NET_0_117236, 
        HIEFFPLA_NET_0_117237, HIEFFPLA_NET_0_117238, 
        HIEFFPLA_NET_0_117239, HIEFFPLA_NET_0_117240, 
        HIEFFPLA_NET_0_117241, HIEFFPLA_NET_0_117242, 
        HIEFFPLA_NET_0_117243, HIEFFPLA_NET_0_117244, 
        HIEFFPLA_NET_0_117245, HIEFFPLA_NET_0_117246, 
        HIEFFPLA_NET_0_117247, HIEFFPLA_NET_0_117248, 
        HIEFFPLA_NET_0_117249, HIEFFPLA_NET_0_117250, 
        HIEFFPLA_NET_0_117251, HIEFFPLA_NET_0_117252, 
        HIEFFPLA_NET_0_117253, HIEFFPLA_NET_0_117254, 
        HIEFFPLA_NET_0_117255, HIEFFPLA_NET_0_117256, 
        HIEFFPLA_NET_0_117257, HIEFFPLA_NET_0_117258, 
        HIEFFPLA_NET_0_117259, HIEFFPLA_NET_0_117260, 
        HIEFFPLA_NET_0_117261, HIEFFPLA_NET_0_117262, 
        HIEFFPLA_NET_0_117263, HIEFFPLA_NET_0_117264, 
        HIEFFPLA_NET_0_117265, HIEFFPLA_NET_0_117266, 
        HIEFFPLA_NET_0_117267, HIEFFPLA_NET_0_117268, 
        HIEFFPLA_NET_0_117269, HIEFFPLA_NET_0_117270, 
        HIEFFPLA_NET_0_117271, HIEFFPLA_NET_0_117272, 
        HIEFFPLA_NET_0_117273, HIEFFPLA_NET_0_117274, 
        HIEFFPLA_NET_0_117275, HIEFFPLA_NET_0_117276, 
        HIEFFPLA_NET_0_117277, HIEFFPLA_NET_0_117278, 
        HIEFFPLA_NET_0_117279, HIEFFPLA_NET_0_117280, 
        HIEFFPLA_NET_0_117281, HIEFFPLA_NET_0_117282, 
        HIEFFPLA_NET_0_117283, HIEFFPLA_NET_0_117284, 
        HIEFFPLA_NET_0_117285, HIEFFPLA_NET_0_117286, 
        HIEFFPLA_NET_0_117287, HIEFFPLA_NET_0_117288, 
        HIEFFPLA_NET_0_117289, HIEFFPLA_NET_0_117290, 
        HIEFFPLA_NET_0_117291, HIEFFPLA_NET_0_117292, 
        HIEFFPLA_NET_0_117293, HIEFFPLA_NET_0_117294, 
        HIEFFPLA_NET_0_117295, HIEFFPLA_NET_0_117296, 
        HIEFFPLA_NET_0_117297, HIEFFPLA_NET_0_117298, 
        HIEFFPLA_NET_0_117299, HIEFFPLA_NET_0_117300, 
        HIEFFPLA_NET_0_117301, HIEFFPLA_NET_0_117302, 
        HIEFFPLA_NET_0_117303, HIEFFPLA_NET_0_117304, 
        HIEFFPLA_NET_0_117305, HIEFFPLA_NET_0_117306, 
        HIEFFPLA_NET_0_117307, HIEFFPLA_NET_0_117308, 
        HIEFFPLA_NET_0_117309, HIEFFPLA_NET_0_117310, 
        HIEFFPLA_NET_0_117311, HIEFFPLA_NET_0_117312, 
        HIEFFPLA_NET_0_117313, HIEFFPLA_NET_0_117314, 
        HIEFFPLA_NET_0_117315, HIEFFPLA_NET_0_117316, 
        HIEFFPLA_NET_0_117317, HIEFFPLA_NET_0_117318, 
        HIEFFPLA_NET_0_117319, HIEFFPLA_NET_0_117320, 
        HIEFFPLA_NET_0_117321, HIEFFPLA_NET_0_117322, 
        HIEFFPLA_NET_0_117323, HIEFFPLA_NET_0_117324, 
        HIEFFPLA_NET_0_117325, HIEFFPLA_NET_0_117326, 
        HIEFFPLA_NET_0_117327, HIEFFPLA_NET_0_117328, 
        HIEFFPLA_NET_0_117329, HIEFFPLA_NET_0_117330, 
        HIEFFPLA_NET_0_117331, HIEFFPLA_NET_0_117332, 
        HIEFFPLA_NET_0_117333, HIEFFPLA_NET_0_117334, 
        HIEFFPLA_NET_0_117335, HIEFFPLA_NET_0_117336, 
        HIEFFPLA_NET_0_117337, HIEFFPLA_NET_0_117338, 
        HIEFFPLA_NET_0_117339, HIEFFPLA_NET_0_117340, 
        HIEFFPLA_NET_0_117341, HIEFFPLA_NET_0_117342, 
        HIEFFPLA_NET_0_117343, HIEFFPLA_NET_0_117344, 
        HIEFFPLA_NET_0_117345, HIEFFPLA_NET_0_117346, 
        HIEFFPLA_NET_0_117347, HIEFFPLA_NET_0_117348, 
        HIEFFPLA_NET_0_117349, HIEFFPLA_NET_0_117350, 
        HIEFFPLA_NET_0_117351, HIEFFPLA_NET_0_117352, 
        HIEFFPLA_NET_0_117353, HIEFFPLA_NET_0_117354, 
        HIEFFPLA_NET_0_117355, HIEFFPLA_NET_0_117356, 
        HIEFFPLA_NET_0_117357, HIEFFPLA_NET_0_117358, 
        HIEFFPLA_NET_0_117359, HIEFFPLA_NET_0_117360, 
        HIEFFPLA_NET_0_117361, HIEFFPLA_NET_0_117362, 
        HIEFFPLA_NET_0_117363, HIEFFPLA_NET_0_117364, 
        HIEFFPLA_NET_0_117365, HIEFFPLA_NET_0_117366, 
        HIEFFPLA_NET_0_117367, HIEFFPLA_NET_0_117368, 
        HIEFFPLA_NET_0_117369, HIEFFPLA_NET_0_117370, 
        HIEFFPLA_NET_0_117371, HIEFFPLA_NET_0_117372, 
        HIEFFPLA_NET_0_117373, HIEFFPLA_NET_0_117374, 
        HIEFFPLA_NET_0_117375, HIEFFPLA_NET_0_117376, 
        HIEFFPLA_NET_0_117377, HIEFFPLA_NET_0_117378, 
        HIEFFPLA_NET_0_117379, HIEFFPLA_NET_0_117380, 
        HIEFFPLA_NET_0_117381, HIEFFPLA_NET_0_117382, 
        HIEFFPLA_NET_0_117383, HIEFFPLA_NET_0_117384, 
        HIEFFPLA_NET_0_117385, HIEFFPLA_NET_0_117386, 
        HIEFFPLA_NET_0_117387, HIEFFPLA_NET_0_117388, 
        HIEFFPLA_NET_0_117389, HIEFFPLA_NET_0_117390, 
        HIEFFPLA_NET_0_117391, HIEFFPLA_NET_0_117392, 
        HIEFFPLA_NET_0_117393, HIEFFPLA_NET_0_117394, 
        HIEFFPLA_NET_0_117395, HIEFFPLA_NET_0_117396, 
        HIEFFPLA_NET_0_117397, HIEFFPLA_NET_0_117398, 
        HIEFFPLA_NET_0_117399, HIEFFPLA_NET_0_117400, 
        HIEFFPLA_NET_0_117401, HIEFFPLA_NET_0_117402, 
        HIEFFPLA_NET_0_117403, HIEFFPLA_NET_0_117404, 
        HIEFFPLA_NET_0_117405, HIEFFPLA_NET_0_117406, 
        HIEFFPLA_NET_0_117407, HIEFFPLA_NET_0_117408, 
        HIEFFPLA_NET_0_117409, HIEFFPLA_NET_0_117410, 
        HIEFFPLA_NET_0_117411, HIEFFPLA_NET_0_117412, 
        HIEFFPLA_NET_0_117413, HIEFFPLA_NET_0_117414, 
        HIEFFPLA_NET_0_117415, HIEFFPLA_NET_0_117416, 
        HIEFFPLA_NET_0_117417, HIEFFPLA_NET_0_117418, 
        HIEFFPLA_NET_0_117419, HIEFFPLA_NET_0_117420, 
        HIEFFPLA_NET_0_117421, HIEFFPLA_NET_0_117422, 
        HIEFFPLA_NET_0_117423, HIEFFPLA_NET_0_117424, 
        HIEFFPLA_NET_0_117425, HIEFFPLA_NET_0_117426, 
        HIEFFPLA_NET_0_117427, HIEFFPLA_NET_0_117428, 
        HIEFFPLA_NET_0_117429, HIEFFPLA_NET_0_117430, 
        HIEFFPLA_NET_0_117431, HIEFFPLA_NET_0_117432, 
        HIEFFPLA_NET_0_117433, HIEFFPLA_NET_0_117434, 
        HIEFFPLA_NET_0_117435, HIEFFPLA_NET_0_117436, 
        HIEFFPLA_NET_0_117437, HIEFFPLA_NET_0_117438, 
        HIEFFPLA_NET_0_117439, HIEFFPLA_NET_0_117440, 
        HIEFFPLA_NET_0_117441, HIEFFPLA_NET_0_117442, 
        HIEFFPLA_NET_0_117443, HIEFFPLA_NET_0_117444, 
        HIEFFPLA_NET_0_117445, HIEFFPLA_NET_0_117446, 
        HIEFFPLA_NET_0_117447, HIEFFPLA_NET_0_117448, 
        HIEFFPLA_NET_0_117449, HIEFFPLA_NET_0_117450, 
        HIEFFPLA_NET_0_117451, HIEFFPLA_NET_0_117452, 
        HIEFFPLA_NET_0_117453, HIEFFPLA_NET_0_117454, 
        HIEFFPLA_NET_0_117455, HIEFFPLA_NET_0_117456, 
        HIEFFPLA_NET_0_117457, HIEFFPLA_NET_0_117458, 
        HIEFFPLA_NET_0_117459, HIEFFPLA_NET_0_117460, 
        HIEFFPLA_NET_0_117461, HIEFFPLA_NET_0_117462, 
        HIEFFPLA_NET_0_117463, HIEFFPLA_NET_0_117464, 
        HIEFFPLA_NET_0_117465, HIEFFPLA_NET_0_117466, 
        HIEFFPLA_NET_0_117467, HIEFFPLA_NET_0_117468, 
        HIEFFPLA_NET_0_117469, HIEFFPLA_NET_0_117470, 
        HIEFFPLA_NET_0_117471, HIEFFPLA_NET_0_117472, 
        HIEFFPLA_NET_0_117473, HIEFFPLA_NET_0_117474, 
        HIEFFPLA_NET_0_117475, HIEFFPLA_NET_0_117476, 
        HIEFFPLA_NET_0_117477, HIEFFPLA_NET_0_117478, 
        HIEFFPLA_NET_0_117479, HIEFFPLA_NET_0_117480, 
        HIEFFPLA_NET_0_117481, HIEFFPLA_NET_0_117482, 
        HIEFFPLA_NET_0_117483, HIEFFPLA_NET_0_117484, 
        HIEFFPLA_NET_0_117485, HIEFFPLA_NET_0_117486, 
        HIEFFPLA_NET_0_117487, HIEFFPLA_NET_0_117488, 
        HIEFFPLA_NET_0_117489, HIEFFPLA_NET_0_117490, 
        HIEFFPLA_NET_0_117491, HIEFFPLA_NET_0_117492, 
        HIEFFPLA_NET_0_117493, HIEFFPLA_NET_0_117494, 
        HIEFFPLA_NET_0_117495, HIEFFPLA_NET_0_117496, 
        HIEFFPLA_NET_0_117497, HIEFFPLA_NET_0_117498, 
        HIEFFPLA_NET_0_117499, HIEFFPLA_NET_0_117500, 
        HIEFFPLA_NET_0_117501, HIEFFPLA_NET_0_117502, 
        HIEFFPLA_NET_0_117503, HIEFFPLA_NET_0_117504, 
        HIEFFPLA_NET_0_117505, HIEFFPLA_NET_0_117506, 
        HIEFFPLA_NET_0_117507, HIEFFPLA_NET_0_117508, 
        HIEFFPLA_NET_0_117509, HIEFFPLA_NET_0_117510, 
        HIEFFPLA_NET_0_117511, HIEFFPLA_NET_0_117512, 
        HIEFFPLA_NET_0_117513, HIEFFPLA_NET_0_117514, 
        HIEFFPLA_NET_0_117515, HIEFFPLA_NET_0_117516, 
        HIEFFPLA_NET_0_117517, HIEFFPLA_NET_0_117518, 
        HIEFFPLA_NET_0_117519, HIEFFPLA_NET_0_117520, 
        HIEFFPLA_NET_0_117521, HIEFFPLA_NET_0_117522, 
        HIEFFPLA_NET_0_117523, HIEFFPLA_NET_0_117524, 
        HIEFFPLA_NET_0_117525, HIEFFPLA_NET_0_117526, 
        HIEFFPLA_NET_0_117527, HIEFFPLA_NET_0_117528, 
        HIEFFPLA_NET_0_117529, HIEFFPLA_NET_0_117530, 
        HIEFFPLA_NET_0_117531, HIEFFPLA_NET_0_117532, 
        HIEFFPLA_NET_0_117533, HIEFFPLA_NET_0_117534, 
        HIEFFPLA_NET_0_117535, HIEFFPLA_NET_0_117536, 
        HIEFFPLA_NET_0_117537, HIEFFPLA_NET_0_117538, 
        HIEFFPLA_NET_0_117539, HIEFFPLA_NET_0_117540, 
        HIEFFPLA_NET_0_117541, HIEFFPLA_NET_0_117542, 
        HIEFFPLA_NET_0_117543, HIEFFPLA_NET_0_117544, 
        HIEFFPLA_NET_0_117545, HIEFFPLA_NET_0_117546, 
        HIEFFPLA_NET_0_117547, HIEFFPLA_NET_0_117548, 
        HIEFFPLA_NET_0_117549, HIEFFPLA_NET_0_117550, 
        HIEFFPLA_NET_0_117551, HIEFFPLA_NET_0_117552, 
        HIEFFPLA_NET_0_117553, HIEFFPLA_NET_0_117554, 
        HIEFFPLA_NET_0_117555, HIEFFPLA_NET_0_117556, 
        HIEFFPLA_NET_0_117557, HIEFFPLA_NET_0_117558, 
        HIEFFPLA_NET_0_117559, HIEFFPLA_NET_0_117560, 
        HIEFFPLA_NET_0_117561, HIEFFPLA_NET_0_117562, 
        HIEFFPLA_NET_0_117563, HIEFFPLA_NET_0_117564, 
        HIEFFPLA_NET_0_117565, HIEFFPLA_NET_0_117566, 
        HIEFFPLA_NET_0_117567, HIEFFPLA_NET_0_117568, 
        HIEFFPLA_NET_0_117569, HIEFFPLA_NET_0_117570, 
        HIEFFPLA_NET_0_117571, HIEFFPLA_NET_0_117572, 
        HIEFFPLA_NET_0_117573, HIEFFPLA_NET_0_117574, 
        HIEFFPLA_NET_0_117575, HIEFFPLA_NET_0_117576, 
        HIEFFPLA_NET_0_117577, HIEFFPLA_NET_0_117578, 
        HIEFFPLA_NET_0_117579, HIEFFPLA_NET_0_117580, 
        HIEFFPLA_NET_0_117581, HIEFFPLA_NET_0_117582, 
        HIEFFPLA_NET_0_117583, HIEFFPLA_NET_0_117584, 
        HIEFFPLA_NET_0_117585, HIEFFPLA_NET_0_117586, 
        HIEFFPLA_NET_0_117587, HIEFFPLA_NET_0_117588, 
        HIEFFPLA_NET_0_117589, HIEFFPLA_NET_0_117590, 
        HIEFFPLA_NET_0_117591, HIEFFPLA_NET_0_117592, 
        HIEFFPLA_NET_0_117593, HIEFFPLA_NET_0_117594, 
        HIEFFPLA_NET_0_117595, HIEFFPLA_NET_0_117596, 
        HIEFFPLA_NET_0_117597, HIEFFPLA_NET_0_117598, 
        HIEFFPLA_NET_0_117599, HIEFFPLA_NET_0_117600, 
        HIEFFPLA_NET_0_117601, HIEFFPLA_NET_0_117602, 
        HIEFFPLA_NET_0_117603, HIEFFPLA_NET_0_117604, 
        HIEFFPLA_NET_0_117605, HIEFFPLA_NET_0_117606, 
        HIEFFPLA_NET_0_117607, HIEFFPLA_NET_0_117609, 
        HIEFFPLA_NET_0_117610, HIEFFPLA_NET_0_117611, 
        HIEFFPLA_NET_0_117612, HIEFFPLA_NET_0_117613, 
        HIEFFPLA_NET_0_117614, HIEFFPLA_NET_0_117615, 
        HIEFFPLA_NET_0_117616, HIEFFPLA_NET_0_117617, 
        HIEFFPLA_NET_0_117618, HIEFFPLA_NET_0_117619, 
        HIEFFPLA_NET_0_117620, HIEFFPLA_NET_0_117621, 
        HIEFFPLA_NET_0_117622, HIEFFPLA_NET_0_117623, 
        HIEFFPLA_NET_0_117624, HIEFFPLA_NET_0_117625, 
        HIEFFPLA_NET_0_117626, HIEFFPLA_NET_0_117627, 
        HIEFFPLA_NET_0_117628, HIEFFPLA_NET_0_117629, 
        HIEFFPLA_NET_0_117630, HIEFFPLA_NET_0_117631, 
        HIEFFPLA_NET_0_117632, HIEFFPLA_NET_0_117633, 
        HIEFFPLA_NET_0_117634, HIEFFPLA_NET_0_117635, 
        HIEFFPLA_NET_0_117636, HIEFFPLA_NET_0_117637, 
        HIEFFPLA_NET_0_117638, HIEFFPLA_NET_0_117639, 
        HIEFFPLA_NET_0_117640, HIEFFPLA_NET_0_117641, 
        HIEFFPLA_NET_0_117642, HIEFFPLA_NET_0_117643, 
        HIEFFPLA_NET_0_117644, HIEFFPLA_NET_0_117645, 
        HIEFFPLA_NET_0_117646, HIEFFPLA_NET_0_117647, 
        HIEFFPLA_NET_0_117648, HIEFFPLA_NET_0_117649, 
        HIEFFPLA_NET_0_117650, HIEFFPLA_NET_0_117651, 
        HIEFFPLA_NET_0_117652, HIEFFPLA_NET_0_117653, 
        HIEFFPLA_NET_0_117654, HIEFFPLA_NET_0_117655, 
        HIEFFPLA_NET_0_117656, HIEFFPLA_NET_0_117657, 
        HIEFFPLA_NET_0_117658, HIEFFPLA_NET_0_117659, 
        HIEFFPLA_NET_0_117660, HIEFFPLA_NET_0_117661, 
        HIEFFPLA_NET_0_117662, HIEFFPLA_NET_0_117663, 
        HIEFFPLA_NET_0_117664, HIEFFPLA_NET_0_117665, 
        HIEFFPLA_NET_0_117666, HIEFFPLA_NET_0_117667, 
        HIEFFPLA_NET_0_117668, HIEFFPLA_NET_0_117669, 
        HIEFFPLA_NET_0_117670, HIEFFPLA_NET_0_117671, 
        HIEFFPLA_NET_0_117672, HIEFFPLA_NET_0_117673, 
        HIEFFPLA_NET_0_117674, HIEFFPLA_NET_0_117675, 
        HIEFFPLA_NET_0_117676, HIEFFPLA_NET_0_117677, 
        HIEFFPLA_NET_0_117678, HIEFFPLA_NET_0_117679, 
        HIEFFPLA_NET_0_117680, HIEFFPLA_NET_0_117681, 
        HIEFFPLA_NET_0_117682, HIEFFPLA_NET_0_117683, 
        HIEFFPLA_NET_0_117684, HIEFFPLA_NET_0_117685, 
        HIEFFPLA_NET_0_117686, HIEFFPLA_NET_0_117687, 
        HIEFFPLA_NET_0_117688, HIEFFPLA_NET_0_117689, 
        HIEFFPLA_NET_0_117690, HIEFFPLA_NET_0_117691, 
        HIEFFPLA_NET_0_117692, HIEFFPLA_NET_0_117693, 
        HIEFFPLA_NET_0_117694, HIEFFPLA_NET_0_117695, 
        HIEFFPLA_NET_0_117696, HIEFFPLA_NET_0_117697, 
        HIEFFPLA_NET_0_117698, HIEFFPLA_NET_0_117699, 
        HIEFFPLA_NET_0_117700, HIEFFPLA_NET_0_117701, 
        HIEFFPLA_NET_0_117702, HIEFFPLA_NET_0_117703, 
        HIEFFPLA_NET_0_117704, HIEFFPLA_NET_0_117705, 
        HIEFFPLA_NET_0_117706, HIEFFPLA_NET_0_117707, 
        HIEFFPLA_NET_0_117708, HIEFFPLA_NET_0_117709, 
        HIEFFPLA_NET_0_117710, HIEFFPLA_NET_0_117711, 
        HIEFFPLA_NET_0_117712, HIEFFPLA_NET_0_117713, 
        HIEFFPLA_NET_0_117714, HIEFFPLA_NET_0_117715, 
        HIEFFPLA_NET_0_117716, HIEFFPLA_NET_0_117717, 
        HIEFFPLA_NET_0_117718, HIEFFPLA_NET_0_117719, 
        HIEFFPLA_NET_0_117720, HIEFFPLA_NET_0_117721, 
        HIEFFPLA_NET_0_117722, HIEFFPLA_NET_0_117723, 
        HIEFFPLA_NET_0_117724, HIEFFPLA_NET_0_117725, 
        HIEFFPLA_NET_0_117726, HIEFFPLA_NET_0_117727, 
        HIEFFPLA_NET_0_117728, HIEFFPLA_NET_0_117729, 
        HIEFFPLA_NET_0_117730, HIEFFPLA_NET_0_117731, 
        HIEFFPLA_NET_0_117732, HIEFFPLA_NET_0_117733, 
        HIEFFPLA_NET_0_117734, HIEFFPLA_NET_0_117735, 
        HIEFFPLA_NET_0_117736, HIEFFPLA_NET_0_117737, 
        HIEFFPLA_NET_0_117738, HIEFFPLA_NET_0_117739, 
        HIEFFPLA_NET_0_117740, HIEFFPLA_NET_0_117741, 
        HIEFFPLA_NET_0_117742, HIEFFPLA_NET_0_117743, 
        HIEFFPLA_NET_0_117744, HIEFFPLA_NET_0_117745, 
        HIEFFPLA_NET_0_117746, HIEFFPLA_NET_0_117747, 
        HIEFFPLA_NET_0_117748, HIEFFPLA_NET_0_117749, 
        HIEFFPLA_NET_0_117750, HIEFFPLA_NET_0_117751, 
        HIEFFPLA_NET_0_117752, HIEFFPLA_NET_0_117753, 
        HIEFFPLA_NET_0_117754, HIEFFPLA_NET_0_117755, 
        HIEFFPLA_NET_0_117756, HIEFFPLA_NET_0_117757, 
        HIEFFPLA_NET_0_117758, HIEFFPLA_NET_0_117759, 
        HIEFFPLA_NET_0_117760, HIEFFPLA_NET_0_117761, 
        HIEFFPLA_NET_0_117762, HIEFFPLA_NET_0_117763, 
        HIEFFPLA_NET_0_117764, HIEFFPLA_NET_0_117765, 
        HIEFFPLA_NET_0_117766, HIEFFPLA_NET_0_117767, 
        HIEFFPLA_NET_0_117768, HIEFFPLA_NET_0_117769, 
        HIEFFPLA_NET_0_117770, HIEFFPLA_NET_0_117771, 
        HIEFFPLA_NET_0_117772, HIEFFPLA_NET_0_117773, 
        HIEFFPLA_NET_0_117774, HIEFFPLA_NET_0_117775, 
        HIEFFPLA_NET_0_117776, HIEFFPLA_NET_0_117777, 
        HIEFFPLA_NET_0_117778, HIEFFPLA_NET_0_117779, 
        HIEFFPLA_NET_0_117780, HIEFFPLA_NET_0_117781, 
        HIEFFPLA_NET_0_117782, HIEFFPLA_NET_0_117783, 
        HIEFFPLA_NET_0_117784, HIEFFPLA_NET_0_117785, 
        HIEFFPLA_NET_0_117786, HIEFFPLA_NET_0_117787, 
        HIEFFPLA_NET_0_117788, HIEFFPLA_NET_0_117789, 
        HIEFFPLA_NET_0_117790, HIEFFPLA_NET_0_117791, 
        HIEFFPLA_NET_0_117792, HIEFFPLA_NET_0_117793, 
        HIEFFPLA_NET_0_117794, HIEFFPLA_NET_0_117795, 
        HIEFFPLA_NET_0_117796, HIEFFPLA_NET_0_117797, 
        HIEFFPLA_NET_0_117798, HIEFFPLA_NET_0_117799, 
        HIEFFPLA_NET_0_117800, HIEFFPLA_NET_0_117801, 
        HIEFFPLA_NET_0_117810, HIEFFPLA_NET_0_117811, 
        HIEFFPLA_NET_0_117812, HIEFFPLA_NET_0_117813, 
        HIEFFPLA_NET_0_117814, HIEFFPLA_NET_0_117815, 
        HIEFFPLA_NET_0_117816, HIEFFPLA_NET_0_117817, 
        HIEFFPLA_NET_0_117818, HIEFFPLA_NET_0_117819, 
        HIEFFPLA_NET_0_117820, HIEFFPLA_NET_0_117821, 
        HIEFFPLA_NET_0_117822, HIEFFPLA_NET_0_117823, 
        HIEFFPLA_NET_0_117824, HIEFFPLA_NET_0_117825, 
        HIEFFPLA_NET_0_117826, HIEFFPLA_NET_0_117827, 
        HIEFFPLA_NET_0_117828, HIEFFPLA_NET_0_117829, 
        HIEFFPLA_NET_0_117830, HIEFFPLA_NET_0_117831, 
        HIEFFPLA_NET_0_117832, HIEFFPLA_NET_0_117833, 
        HIEFFPLA_NET_0_117834, HIEFFPLA_NET_0_117835, 
        HIEFFPLA_NET_0_117836, HIEFFPLA_NET_0_117837, 
        HIEFFPLA_NET_0_117838, HIEFFPLA_NET_0_117839, 
        HIEFFPLA_NET_0_117840, HIEFFPLA_NET_0_117841, 
        HIEFFPLA_NET_0_117842, HIEFFPLA_NET_0_117843, 
        HIEFFPLA_NET_0_117844, HIEFFPLA_NET_0_117845, 
        HIEFFPLA_NET_0_117846, HIEFFPLA_NET_0_117855, 
        HIEFFPLA_NET_0_117856, HIEFFPLA_NET_0_117857, 
        HIEFFPLA_NET_0_117858, HIEFFPLA_NET_0_117859, 
        HIEFFPLA_NET_0_117860, HIEFFPLA_NET_0_117861, 
        HIEFFPLA_NET_0_117862, HIEFFPLA_NET_0_117863, 
        HIEFFPLA_NET_0_117864, HIEFFPLA_NET_0_117865, 
        HIEFFPLA_NET_0_117866, HIEFFPLA_NET_0_117867, 
        HIEFFPLA_NET_0_117868, HIEFFPLA_NET_0_117869, 
        HIEFFPLA_NET_0_117870, HIEFFPLA_NET_0_117871, 
        HIEFFPLA_NET_0_117872, HIEFFPLA_NET_0_117873, 
        HIEFFPLA_NET_0_117874, HIEFFPLA_NET_0_117875, 
        HIEFFPLA_NET_0_117876, HIEFFPLA_NET_0_117877, 
        HIEFFPLA_NET_0_117878, HIEFFPLA_NET_0_117879, 
        HIEFFPLA_NET_0_117880, HIEFFPLA_NET_0_117881, 
        HIEFFPLA_NET_0_117882, HIEFFPLA_NET_0_117883, 
        HIEFFPLA_NET_0_117884, HIEFFPLA_NET_0_117885, 
        HIEFFPLA_NET_0_117886, HIEFFPLA_NET_0_117887, 
        HIEFFPLA_NET_0_117888, HIEFFPLA_NET_0_117889, 
        HIEFFPLA_NET_0_117890, HIEFFPLA_NET_0_117891, 
        HIEFFPLA_NET_0_117900, HIEFFPLA_NET_0_117901, 
        HIEFFPLA_NET_0_117902, HIEFFPLA_NET_0_117903, 
        HIEFFPLA_NET_0_117904, HIEFFPLA_NET_0_117905, 
        HIEFFPLA_NET_0_117906, HIEFFPLA_NET_0_117907, 
        HIEFFPLA_NET_0_117908, HIEFFPLA_NET_0_117909, 
        HIEFFPLA_NET_0_117910, HIEFFPLA_NET_0_117911, 
        HIEFFPLA_NET_0_117912, HIEFFPLA_NET_0_117913, 
        HIEFFPLA_NET_0_117914, HIEFFPLA_NET_0_117915, 
        HIEFFPLA_NET_0_117916, HIEFFPLA_NET_0_117917, 
        HIEFFPLA_NET_0_117918, HIEFFPLA_NET_0_117919, 
        HIEFFPLA_NET_0_117920, HIEFFPLA_NET_0_117921, 
        HIEFFPLA_NET_0_117922, HIEFFPLA_NET_0_117923, 
        HIEFFPLA_NET_0_117924, HIEFFPLA_NET_0_117925, 
        HIEFFPLA_NET_0_117926, HIEFFPLA_NET_0_117927, 
        HIEFFPLA_NET_0_117928, HIEFFPLA_NET_0_117929, 
        HIEFFPLA_NET_0_117930, HIEFFPLA_NET_0_117931, 
        HIEFFPLA_NET_0_117932, HIEFFPLA_NET_0_117933, 
        HIEFFPLA_NET_0_117934, HIEFFPLA_NET_0_117935, 
        HIEFFPLA_NET_0_117936, HIEFFPLA_NET_0_117945, 
        HIEFFPLA_NET_0_117946, HIEFFPLA_NET_0_117947, 
        HIEFFPLA_NET_0_117948, HIEFFPLA_NET_0_117949, 
        HIEFFPLA_NET_0_117950, HIEFFPLA_NET_0_117951, 
        HIEFFPLA_NET_0_117952, HIEFFPLA_NET_0_117953, 
        HIEFFPLA_NET_0_117954, HIEFFPLA_NET_0_117955, 
        HIEFFPLA_NET_0_117956, HIEFFPLA_NET_0_117957, 
        HIEFFPLA_NET_0_117958, HIEFFPLA_NET_0_117959, 
        HIEFFPLA_NET_0_117960, HIEFFPLA_NET_0_117961, 
        HIEFFPLA_NET_0_117962, HIEFFPLA_NET_0_117963, 
        HIEFFPLA_NET_0_117964, HIEFFPLA_NET_0_117965, 
        HIEFFPLA_NET_0_117966, HIEFFPLA_NET_0_117967, 
        HIEFFPLA_NET_0_117968, HIEFFPLA_NET_0_117969, 
        HIEFFPLA_NET_0_117970, HIEFFPLA_NET_0_117971, 
        HIEFFPLA_NET_0_117972, HIEFFPLA_NET_0_117973, 
        HIEFFPLA_NET_0_117974, HIEFFPLA_NET_0_117975, 
        HIEFFPLA_NET_0_117976, HIEFFPLA_NET_0_117977, 
        HIEFFPLA_NET_0_117978, HIEFFPLA_NET_0_117979, 
        HIEFFPLA_NET_0_117980, HIEFFPLA_NET_0_117981, 
        HIEFFPLA_NET_0_117990, HIEFFPLA_NET_0_117991, 
        HIEFFPLA_NET_0_117992, HIEFFPLA_NET_0_117993, 
        HIEFFPLA_NET_0_117994, HIEFFPLA_NET_0_117995, 
        HIEFFPLA_NET_0_117996, HIEFFPLA_NET_0_117997, 
        HIEFFPLA_NET_0_117998, HIEFFPLA_NET_0_117999, 
        HIEFFPLA_NET_0_118000, HIEFFPLA_NET_0_118001, 
        HIEFFPLA_NET_0_118002, HIEFFPLA_NET_0_118003, 
        HIEFFPLA_NET_0_118004, HIEFFPLA_NET_0_118005, 
        HIEFFPLA_NET_0_118006, HIEFFPLA_NET_0_118007, 
        HIEFFPLA_NET_0_118008, HIEFFPLA_NET_0_118009, 
        HIEFFPLA_NET_0_118010, HIEFFPLA_NET_0_118011, 
        HIEFFPLA_NET_0_118012, HIEFFPLA_NET_0_118013, 
        HIEFFPLA_NET_0_118014, HIEFFPLA_NET_0_118015, 
        HIEFFPLA_NET_0_118016, HIEFFPLA_NET_0_118017, 
        HIEFFPLA_NET_0_118018, HIEFFPLA_NET_0_118019, 
        HIEFFPLA_NET_0_118020, HIEFFPLA_NET_0_118021, 
        HIEFFPLA_NET_0_118022, HIEFFPLA_NET_0_118023, 
        HIEFFPLA_NET_0_118024, HIEFFPLA_NET_0_118025, 
        HIEFFPLA_NET_0_118026, HIEFFPLA_NET_0_118035, 
        HIEFFPLA_NET_0_118036, HIEFFPLA_NET_0_118037, 
        HIEFFPLA_NET_0_118038, HIEFFPLA_NET_0_118039, 
        HIEFFPLA_NET_0_118040, HIEFFPLA_NET_0_118041, 
        HIEFFPLA_NET_0_118042, HIEFFPLA_NET_0_118043, 
        HIEFFPLA_NET_0_118044, HIEFFPLA_NET_0_118045, 
        HIEFFPLA_NET_0_118046, HIEFFPLA_NET_0_118047, 
        HIEFFPLA_NET_0_118048, HIEFFPLA_NET_0_118049, 
        HIEFFPLA_NET_0_118050, HIEFFPLA_NET_0_118051, 
        HIEFFPLA_NET_0_118052, HIEFFPLA_NET_0_118053, 
        HIEFFPLA_NET_0_118054, HIEFFPLA_NET_0_118055, 
        HIEFFPLA_NET_0_118056, HIEFFPLA_NET_0_118057, 
        HIEFFPLA_NET_0_118058, HIEFFPLA_NET_0_118059, 
        HIEFFPLA_NET_0_118060, HIEFFPLA_NET_0_118061, 
        HIEFFPLA_NET_0_118062, HIEFFPLA_NET_0_118063, 
        HIEFFPLA_NET_0_118064, HIEFFPLA_NET_0_118065, 
        HIEFFPLA_NET_0_118066, HIEFFPLA_NET_0_118067, 
        HIEFFPLA_NET_0_118068, HIEFFPLA_NET_0_118069, 
        HIEFFPLA_NET_0_118070, HIEFFPLA_NET_0_118071, 
        HIEFFPLA_NET_0_118080, HIEFFPLA_NET_0_118081, 
        HIEFFPLA_NET_0_118082, HIEFFPLA_NET_0_118083, 
        HIEFFPLA_NET_0_118084, HIEFFPLA_NET_0_118085, 
        HIEFFPLA_NET_0_118086, HIEFFPLA_NET_0_118087, 
        HIEFFPLA_NET_0_118088, HIEFFPLA_NET_0_118089, 
        HIEFFPLA_NET_0_118090, HIEFFPLA_NET_0_118091, 
        HIEFFPLA_NET_0_118092, HIEFFPLA_NET_0_118093, 
        HIEFFPLA_NET_0_118094, HIEFFPLA_NET_0_118095, 
        HIEFFPLA_NET_0_118096, HIEFFPLA_NET_0_118097, 
        HIEFFPLA_NET_0_118098, HIEFFPLA_NET_0_118099, 
        HIEFFPLA_NET_0_118100, HIEFFPLA_NET_0_118101, 
        HIEFFPLA_NET_0_118102, HIEFFPLA_NET_0_118103, 
        HIEFFPLA_NET_0_118104, HIEFFPLA_NET_0_118105, 
        HIEFFPLA_NET_0_118106, HIEFFPLA_NET_0_118107, 
        HIEFFPLA_NET_0_118108, HIEFFPLA_NET_0_118109, 
        HIEFFPLA_NET_0_118110, HIEFFPLA_NET_0_118111, 
        HIEFFPLA_NET_0_118112, HIEFFPLA_NET_0_118113, 
        HIEFFPLA_NET_0_118114, HIEFFPLA_NET_0_118115, 
        HIEFFPLA_NET_0_118116, HIEFFPLA_NET_0_118125, 
        HIEFFPLA_NET_0_118126, HIEFFPLA_NET_0_118127, 
        HIEFFPLA_NET_0_118128, HIEFFPLA_NET_0_118129, 
        HIEFFPLA_NET_0_118130, HIEFFPLA_NET_0_118131, 
        HIEFFPLA_NET_0_118132, HIEFFPLA_NET_0_118133, 
        HIEFFPLA_NET_0_118134, HIEFFPLA_NET_0_118135, 
        HIEFFPLA_NET_0_118136, HIEFFPLA_NET_0_118137, 
        HIEFFPLA_NET_0_118138, HIEFFPLA_NET_0_118139, 
        HIEFFPLA_NET_0_118140, HIEFFPLA_NET_0_118141, 
        HIEFFPLA_NET_0_118142, HIEFFPLA_NET_0_118143, 
        HIEFFPLA_NET_0_118144, HIEFFPLA_NET_0_118145, 
        HIEFFPLA_NET_0_118146, HIEFFPLA_NET_0_118147, 
        HIEFFPLA_NET_0_118148, HIEFFPLA_NET_0_118149, 
        HIEFFPLA_NET_0_118150, HIEFFPLA_NET_0_118151, 
        HIEFFPLA_NET_0_118152, HIEFFPLA_NET_0_118153, 
        HIEFFPLA_NET_0_118154, HIEFFPLA_NET_0_118155, 
        HIEFFPLA_NET_0_118156, HIEFFPLA_NET_0_118157, 
        HIEFFPLA_NET_0_118158, HIEFFPLA_NET_0_118159, 
        HIEFFPLA_NET_0_118160, HIEFFPLA_NET_0_118161, 
        HIEFFPLA_NET_0_118170, HIEFFPLA_NET_0_118171, 
        HIEFFPLA_NET_0_118172, HIEFFPLA_NET_0_118173, 
        HIEFFPLA_NET_0_118174, HIEFFPLA_NET_0_118175, 
        HIEFFPLA_NET_0_118176, HIEFFPLA_NET_0_118177, 
        HIEFFPLA_NET_0_118178, HIEFFPLA_NET_0_118179, 
        HIEFFPLA_NET_0_118180, HIEFFPLA_NET_0_118181, 
        HIEFFPLA_NET_0_118182, HIEFFPLA_NET_0_118183, 
        HIEFFPLA_NET_0_118184, HIEFFPLA_NET_0_118185, 
        HIEFFPLA_NET_0_118186, HIEFFPLA_NET_0_118187, 
        HIEFFPLA_NET_0_118188, HIEFFPLA_NET_0_118189, 
        HIEFFPLA_NET_0_118190, HIEFFPLA_NET_0_118191, 
        HIEFFPLA_NET_0_118192, HIEFFPLA_NET_0_118193, 
        HIEFFPLA_NET_0_118194, HIEFFPLA_NET_0_118195, 
        HIEFFPLA_NET_0_118196, HIEFFPLA_NET_0_118197, 
        HIEFFPLA_NET_0_118198, HIEFFPLA_NET_0_118199, 
        HIEFFPLA_NET_0_118200, HIEFFPLA_NET_0_118201, 
        HIEFFPLA_NET_0_118202, HIEFFPLA_NET_0_118203, 
        HIEFFPLA_NET_0_118204, HIEFFPLA_NET_0_118205, 
        HIEFFPLA_NET_0_118206, HIEFFPLA_NET_0_118215, 
        HIEFFPLA_NET_0_118216, HIEFFPLA_NET_0_118217, 
        HIEFFPLA_NET_0_118218, HIEFFPLA_NET_0_118219, 
        HIEFFPLA_NET_0_118220, HIEFFPLA_NET_0_118221, 
        HIEFFPLA_NET_0_118222, HIEFFPLA_NET_0_118223, 
        HIEFFPLA_NET_0_118224, HIEFFPLA_NET_0_118225, 
        HIEFFPLA_NET_0_118226, HIEFFPLA_NET_0_118227, 
        HIEFFPLA_NET_0_118228, HIEFFPLA_NET_0_118229, 
        HIEFFPLA_NET_0_118230, HIEFFPLA_NET_0_118231, 
        HIEFFPLA_NET_0_118232, HIEFFPLA_NET_0_118233, 
        HIEFFPLA_NET_0_118234, HIEFFPLA_NET_0_118235, 
        HIEFFPLA_NET_0_118236, HIEFFPLA_NET_0_118237, 
        HIEFFPLA_NET_0_118238, HIEFFPLA_NET_0_118239, 
        HIEFFPLA_NET_0_118240, HIEFFPLA_NET_0_118241, 
        HIEFFPLA_NET_0_118242, HIEFFPLA_NET_0_118243, 
        HIEFFPLA_NET_0_118244, HIEFFPLA_NET_0_118245, 
        HIEFFPLA_NET_0_118246, HIEFFPLA_NET_0_118247, 
        HIEFFPLA_NET_0_118248, HIEFFPLA_NET_0_118249, 
        HIEFFPLA_NET_0_118250, HIEFFPLA_NET_0_118251, 
        HIEFFPLA_NET_0_118260, HIEFFPLA_NET_0_118261, 
        HIEFFPLA_NET_0_118262, HIEFFPLA_NET_0_118263, 
        HIEFFPLA_NET_0_118264, HIEFFPLA_NET_0_118265, 
        HIEFFPLA_NET_0_118266, HIEFFPLA_NET_0_118267, 
        HIEFFPLA_NET_0_118268, HIEFFPLA_NET_0_118269, 
        HIEFFPLA_NET_0_118270, HIEFFPLA_NET_0_118271, 
        HIEFFPLA_NET_0_118272, HIEFFPLA_NET_0_118273, 
        HIEFFPLA_NET_0_118274, HIEFFPLA_NET_0_118275, 
        HIEFFPLA_NET_0_118276, HIEFFPLA_NET_0_118277, 
        HIEFFPLA_NET_0_118278, HIEFFPLA_NET_0_118279, 
        HIEFFPLA_NET_0_118280, HIEFFPLA_NET_0_118281, 
        HIEFFPLA_NET_0_118282, HIEFFPLA_NET_0_118283, 
        HIEFFPLA_NET_0_118284, HIEFFPLA_NET_0_118285, 
        HIEFFPLA_NET_0_118286, HIEFFPLA_NET_0_118287, 
        HIEFFPLA_NET_0_118288, HIEFFPLA_NET_0_118289, 
        HIEFFPLA_NET_0_118290, HIEFFPLA_NET_0_118291, 
        HIEFFPLA_NET_0_118292, HIEFFPLA_NET_0_118293, 
        HIEFFPLA_NET_0_118294, HIEFFPLA_NET_0_118295, 
        HIEFFPLA_NET_0_118296, HIEFFPLA_NET_0_118305, 
        HIEFFPLA_NET_0_118306, HIEFFPLA_NET_0_118307, 
        HIEFFPLA_NET_0_118308, HIEFFPLA_NET_0_118309, 
        HIEFFPLA_NET_0_118310, HIEFFPLA_NET_0_118311, 
        HIEFFPLA_NET_0_118312, HIEFFPLA_NET_0_118313, 
        HIEFFPLA_NET_0_118314, HIEFFPLA_NET_0_118315, 
        HIEFFPLA_NET_0_118316, HIEFFPLA_NET_0_118317, 
        HIEFFPLA_NET_0_118318, HIEFFPLA_NET_0_118319, 
        HIEFFPLA_NET_0_118320, HIEFFPLA_NET_0_118321, 
        HIEFFPLA_NET_0_118322, HIEFFPLA_NET_0_118323, 
        HIEFFPLA_NET_0_118324, HIEFFPLA_NET_0_118325, 
        HIEFFPLA_NET_0_118326, HIEFFPLA_NET_0_118327, 
        HIEFFPLA_NET_0_118328, HIEFFPLA_NET_0_118329, 
        HIEFFPLA_NET_0_118330, HIEFFPLA_NET_0_118331, 
        HIEFFPLA_NET_0_118332, HIEFFPLA_NET_0_118333, 
        HIEFFPLA_NET_0_118334, HIEFFPLA_NET_0_118335, 
        HIEFFPLA_NET_0_118336, HIEFFPLA_NET_0_118337, 
        HIEFFPLA_NET_0_118338, HIEFFPLA_NET_0_118339, 
        HIEFFPLA_NET_0_118340, HIEFFPLA_NET_0_118341, 
        HIEFFPLA_NET_0_118350, HIEFFPLA_NET_0_118351, 
        HIEFFPLA_NET_0_118352, HIEFFPLA_NET_0_118353, 
        HIEFFPLA_NET_0_118354, HIEFFPLA_NET_0_118355, 
        HIEFFPLA_NET_0_118356, HIEFFPLA_NET_0_118357, 
        HIEFFPLA_NET_0_118358, HIEFFPLA_NET_0_118359, 
        HIEFFPLA_NET_0_118360, HIEFFPLA_NET_0_118361, 
        HIEFFPLA_NET_0_118362, HIEFFPLA_NET_0_118363, 
        HIEFFPLA_NET_0_118364, HIEFFPLA_NET_0_118365, 
        HIEFFPLA_NET_0_118366, HIEFFPLA_NET_0_118367, 
        HIEFFPLA_NET_0_118368, HIEFFPLA_NET_0_118369, 
        HIEFFPLA_NET_0_118370, HIEFFPLA_NET_0_118371, 
        HIEFFPLA_NET_0_118372, HIEFFPLA_NET_0_118373, 
        HIEFFPLA_NET_0_118374, HIEFFPLA_NET_0_118375, 
        HIEFFPLA_NET_0_118376, HIEFFPLA_NET_0_118377, 
        HIEFFPLA_NET_0_118378, HIEFFPLA_NET_0_118379, 
        HIEFFPLA_NET_0_118380, HIEFFPLA_NET_0_118381, 
        HIEFFPLA_NET_0_118382, HIEFFPLA_NET_0_118383, 
        HIEFFPLA_NET_0_118384, HIEFFPLA_NET_0_118385, 
        HIEFFPLA_NET_0_118386, HIEFFPLA_NET_0_118395, 
        HIEFFPLA_NET_0_118396, HIEFFPLA_NET_0_118397, 
        HIEFFPLA_NET_0_118398, HIEFFPLA_NET_0_118399, 
        HIEFFPLA_NET_0_118400, HIEFFPLA_NET_0_118401, 
        HIEFFPLA_NET_0_118402, HIEFFPLA_NET_0_118403, 
        HIEFFPLA_NET_0_118404, HIEFFPLA_NET_0_118405, 
        HIEFFPLA_NET_0_118406, HIEFFPLA_NET_0_118407, 
        HIEFFPLA_NET_0_118408, HIEFFPLA_NET_0_118409, 
        HIEFFPLA_NET_0_118410, HIEFFPLA_NET_0_118411, 
        HIEFFPLA_NET_0_118412, HIEFFPLA_NET_0_118413, 
        HIEFFPLA_NET_0_118414, HIEFFPLA_NET_0_118415, 
        HIEFFPLA_NET_0_118416, HIEFFPLA_NET_0_118417, 
        HIEFFPLA_NET_0_118418, HIEFFPLA_NET_0_118419, 
        HIEFFPLA_NET_0_118420, HIEFFPLA_NET_0_118421, 
        HIEFFPLA_NET_0_118422, HIEFFPLA_NET_0_118423, 
        HIEFFPLA_NET_0_118424, HIEFFPLA_NET_0_118425, 
        HIEFFPLA_NET_0_118426, HIEFFPLA_NET_0_118427, 
        HIEFFPLA_NET_0_118428, HIEFFPLA_NET_0_118429, 
        HIEFFPLA_NET_0_118430, HIEFFPLA_NET_0_118431, 
        HIEFFPLA_NET_0_118440, HIEFFPLA_NET_0_118441, 
        HIEFFPLA_NET_0_118442, HIEFFPLA_NET_0_118443, 
        HIEFFPLA_NET_0_118444, HIEFFPLA_NET_0_118445, 
        HIEFFPLA_NET_0_118446, HIEFFPLA_NET_0_118447, 
        HIEFFPLA_NET_0_118448, HIEFFPLA_NET_0_118449, 
        HIEFFPLA_NET_0_118450, HIEFFPLA_NET_0_118451, 
        HIEFFPLA_NET_0_118452, HIEFFPLA_NET_0_118453, 
        HIEFFPLA_NET_0_118454, HIEFFPLA_NET_0_118455, 
        HIEFFPLA_NET_0_118456, HIEFFPLA_NET_0_118457, 
        HIEFFPLA_NET_0_118458, HIEFFPLA_NET_0_118459, 
        HIEFFPLA_NET_0_118460, HIEFFPLA_NET_0_118461, 
        HIEFFPLA_NET_0_118462, HIEFFPLA_NET_0_118463, 
        HIEFFPLA_NET_0_118464, HIEFFPLA_NET_0_118465, 
        HIEFFPLA_NET_0_118466, HIEFFPLA_NET_0_118467, 
        HIEFFPLA_NET_0_118468, HIEFFPLA_NET_0_118469, 
        HIEFFPLA_NET_0_118470, HIEFFPLA_NET_0_118471, 
        HIEFFPLA_NET_0_118472, HIEFFPLA_NET_0_118473, 
        HIEFFPLA_NET_0_118474, HIEFFPLA_NET_0_118475, 
        HIEFFPLA_NET_0_118476, HIEFFPLA_NET_0_118485, 
        HIEFFPLA_NET_0_118486, HIEFFPLA_NET_0_118487, 
        HIEFFPLA_NET_0_118488, HIEFFPLA_NET_0_118489, 
        HIEFFPLA_NET_0_118490, HIEFFPLA_NET_0_118491, 
        HIEFFPLA_NET_0_118492, HIEFFPLA_NET_0_118493, 
        HIEFFPLA_NET_0_118494, HIEFFPLA_NET_0_118495, 
        HIEFFPLA_NET_0_118496, HIEFFPLA_NET_0_118497, 
        HIEFFPLA_NET_0_118498, HIEFFPLA_NET_0_118499, 
        HIEFFPLA_NET_0_118500, HIEFFPLA_NET_0_118501, 
        HIEFFPLA_NET_0_118502, HIEFFPLA_NET_0_118503, 
        HIEFFPLA_NET_0_118504, HIEFFPLA_NET_0_118505, 
        HIEFFPLA_NET_0_118506, HIEFFPLA_NET_0_118507, 
        HIEFFPLA_NET_0_118508, HIEFFPLA_NET_0_118509, 
        HIEFFPLA_NET_0_118510, HIEFFPLA_NET_0_118511, 
        HIEFFPLA_NET_0_118512, HIEFFPLA_NET_0_118513, 
        HIEFFPLA_NET_0_118514, HIEFFPLA_NET_0_118515, 
        HIEFFPLA_NET_0_118516, HIEFFPLA_NET_0_118517, 
        HIEFFPLA_NET_0_118518, HIEFFPLA_NET_0_118519, 
        HIEFFPLA_NET_0_118520, HIEFFPLA_NET_0_118521, 
        HIEFFPLA_NET_0_118530, HIEFFPLA_NET_0_118531, 
        HIEFFPLA_NET_0_118532, HIEFFPLA_NET_0_118533, 
        HIEFFPLA_NET_0_118534, HIEFFPLA_NET_0_118535, 
        HIEFFPLA_NET_0_118536, HIEFFPLA_NET_0_118537, 
        HIEFFPLA_NET_0_118538, HIEFFPLA_NET_0_118539, 
        HIEFFPLA_NET_0_118540, HIEFFPLA_NET_0_118541, 
        HIEFFPLA_NET_0_118542, HIEFFPLA_NET_0_118543, 
        HIEFFPLA_NET_0_118544, HIEFFPLA_NET_0_118545, 
        HIEFFPLA_NET_0_118546, HIEFFPLA_NET_0_118547, 
        HIEFFPLA_NET_0_118548, HIEFFPLA_NET_0_118549, 
        HIEFFPLA_NET_0_118550, HIEFFPLA_NET_0_118551, 
        HIEFFPLA_NET_0_118552, HIEFFPLA_NET_0_118553, 
        HIEFFPLA_NET_0_118554, HIEFFPLA_NET_0_118555, 
        HIEFFPLA_NET_0_118556, HIEFFPLA_NET_0_118557, 
        HIEFFPLA_NET_0_118558, HIEFFPLA_NET_0_118559, 
        HIEFFPLA_NET_0_118560, HIEFFPLA_NET_0_118561, 
        HIEFFPLA_NET_0_118562, HIEFFPLA_NET_0_118563, 
        HIEFFPLA_NET_0_118564, HIEFFPLA_NET_0_118565, 
        HIEFFPLA_NET_0_118566, HIEFFPLA_NET_0_118575, 
        HIEFFPLA_NET_0_118576, HIEFFPLA_NET_0_118577, 
        HIEFFPLA_NET_0_118578, HIEFFPLA_NET_0_118579, 
        HIEFFPLA_NET_0_118580, HIEFFPLA_NET_0_118581, 
        HIEFFPLA_NET_0_118582, HIEFFPLA_NET_0_118583, 
        HIEFFPLA_NET_0_118584, HIEFFPLA_NET_0_118585, 
        HIEFFPLA_NET_0_118586, HIEFFPLA_NET_0_118587, 
        HIEFFPLA_NET_0_118588, HIEFFPLA_NET_0_118589, 
        HIEFFPLA_NET_0_118590, HIEFFPLA_NET_0_118591, 
        HIEFFPLA_NET_0_118592, HIEFFPLA_NET_0_118593, 
        HIEFFPLA_NET_0_118594, HIEFFPLA_NET_0_118595, 
        HIEFFPLA_NET_0_118596, HIEFFPLA_NET_0_118597, 
        HIEFFPLA_NET_0_118598, HIEFFPLA_NET_0_118599, 
        HIEFFPLA_NET_0_118600, HIEFFPLA_NET_0_118601, 
        HIEFFPLA_NET_0_118602, HIEFFPLA_NET_0_118603, 
        HIEFFPLA_NET_0_118604, HIEFFPLA_NET_0_118605, 
        HIEFFPLA_NET_0_118606, HIEFFPLA_NET_0_118607, 
        HIEFFPLA_NET_0_118608, HIEFFPLA_NET_0_118609, 
        HIEFFPLA_NET_0_118610, HIEFFPLA_NET_0_118611, 
        HIEFFPLA_NET_0_118620, HIEFFPLA_NET_0_118621, 
        HIEFFPLA_NET_0_118622, HIEFFPLA_NET_0_118623, 
        HIEFFPLA_NET_0_118624, HIEFFPLA_NET_0_118625, 
        HIEFFPLA_NET_0_118626, HIEFFPLA_NET_0_118627, 
        HIEFFPLA_NET_0_118628, HIEFFPLA_NET_0_118629, 
        HIEFFPLA_NET_0_118630, HIEFFPLA_NET_0_118631, 
        HIEFFPLA_NET_0_118632, HIEFFPLA_NET_0_118633, 
        HIEFFPLA_NET_0_118634, HIEFFPLA_NET_0_118635, 
        HIEFFPLA_NET_0_118636, HIEFFPLA_NET_0_118637, 
        HIEFFPLA_NET_0_118638, HIEFFPLA_NET_0_118639, 
        HIEFFPLA_NET_0_118640, HIEFFPLA_NET_0_118641, 
        HIEFFPLA_NET_0_118642, HIEFFPLA_NET_0_118643, 
        HIEFFPLA_NET_0_118644, HIEFFPLA_NET_0_118645, 
        HIEFFPLA_NET_0_118646, HIEFFPLA_NET_0_118647, 
        HIEFFPLA_NET_0_118648, HIEFFPLA_NET_0_118649, 
        HIEFFPLA_NET_0_118650, HIEFFPLA_NET_0_118651, 
        HIEFFPLA_NET_0_118652, HIEFFPLA_NET_0_118653, 
        HIEFFPLA_NET_0_118654, HIEFFPLA_NET_0_118655, 
        HIEFFPLA_NET_0_118656, HIEFFPLA_NET_0_118657, 
        HIEFFPLA_NET_0_118658, HIEFFPLA_NET_0_118659, 
        HIEFFPLA_NET_0_118660, HIEFFPLA_NET_0_118661, 
        HIEFFPLA_NET_0_118662, HIEFFPLA_NET_0_118663, 
        HIEFFPLA_NET_0_118664, HIEFFPLA_NET_0_118665, 
        HIEFFPLA_NET_0_118666, HIEFFPLA_NET_0_118667, 
        HIEFFPLA_NET_0_118668, HIEFFPLA_NET_0_118669, 
        HIEFFPLA_NET_0_118670, HIEFFPLA_NET_0_118671, 
        HIEFFPLA_NET_0_118672, HIEFFPLA_NET_0_118673, 
        HIEFFPLA_NET_0_118674, HIEFFPLA_NET_0_118675, 
        HIEFFPLA_NET_0_118676, HIEFFPLA_NET_0_118677, 
        HIEFFPLA_NET_0_118678, HIEFFPLA_NET_0_118679, 
        HIEFFPLA_NET_0_118680, HIEFFPLA_NET_0_118681, 
        HIEFFPLA_NET_0_118682, HIEFFPLA_NET_0_118683, 
        HIEFFPLA_NET_0_118684, HIEFFPLA_NET_0_118685, 
        HIEFFPLA_NET_0_118686, HIEFFPLA_NET_0_118687, 
        HIEFFPLA_NET_0_118688, HIEFFPLA_NET_0_118689, 
        HIEFFPLA_NET_0_118690, HIEFFPLA_NET_0_118691, 
        HIEFFPLA_NET_0_118692, HIEFFPLA_NET_0_118693, 
        HIEFFPLA_NET_0_118694, HIEFFPLA_NET_0_118695, 
        HIEFFPLA_NET_0_118696, HIEFFPLA_NET_0_118697, 
        HIEFFPLA_NET_0_118698, HIEFFPLA_NET_0_118699, 
        HIEFFPLA_NET_0_118700, HIEFFPLA_NET_0_118701, 
        HIEFFPLA_NET_0_118702, HIEFFPLA_NET_0_118703, 
        HIEFFPLA_NET_0_118704, HIEFFPLA_NET_0_118705, 
        HIEFFPLA_NET_0_118706, HIEFFPLA_NET_0_118707, 
        HIEFFPLA_NET_0_118708, HIEFFPLA_NET_0_118709, 
        HIEFFPLA_NET_0_118710, HIEFFPLA_NET_0_118711, 
        HIEFFPLA_NET_0_118712, HIEFFPLA_NET_0_118713, 
        HIEFFPLA_NET_0_118714, HIEFFPLA_NET_0_118715, 
        HIEFFPLA_NET_0_118716, HIEFFPLA_NET_0_118717, 
        HIEFFPLA_NET_0_118718, HIEFFPLA_NET_0_118719, 
        HIEFFPLA_NET_0_118720, HIEFFPLA_NET_0_118721, 
        HIEFFPLA_NET_0_118722, HIEFFPLA_NET_0_118723, 
        HIEFFPLA_NET_0_118724, HIEFFPLA_NET_0_118725, 
        HIEFFPLA_NET_0_118726, HIEFFPLA_NET_0_118727, 
        HIEFFPLA_NET_0_118728, HIEFFPLA_NET_0_118729, 
        HIEFFPLA_NET_0_118730, HIEFFPLA_NET_0_118731, 
        HIEFFPLA_NET_0_118732, HIEFFPLA_NET_0_118733, 
        HIEFFPLA_NET_0_118734, HIEFFPLA_NET_0_118735, 
        HIEFFPLA_NET_0_118736, HIEFFPLA_NET_0_118737, 
        HIEFFPLA_NET_0_118738, HIEFFPLA_NET_0_118739, 
        HIEFFPLA_NET_0_118740, HIEFFPLA_NET_0_118741, 
        HIEFFPLA_NET_0_118742, HIEFFPLA_NET_0_118743, 
        HIEFFPLA_NET_0_118744, HIEFFPLA_NET_0_118745, 
        HIEFFPLA_NET_0_118746, HIEFFPLA_NET_0_118747, 
        HIEFFPLA_NET_0_118748, HIEFFPLA_NET_0_118749, 
        HIEFFPLA_NET_0_118750, HIEFFPLA_NET_0_118751, 
        HIEFFPLA_NET_0_118752, HIEFFPLA_NET_0_118753, 
        HIEFFPLA_NET_0_118754, HIEFFPLA_NET_0_118755, 
        HIEFFPLA_NET_0_118756, HIEFFPLA_NET_0_118757, 
        HIEFFPLA_NET_0_118758, HIEFFPLA_NET_0_118759, 
        HIEFFPLA_NET_0_118760, HIEFFPLA_NET_0_118761, 
        HIEFFPLA_NET_0_118762, HIEFFPLA_NET_0_118763, 
        HIEFFPLA_NET_0_118764, HIEFFPLA_NET_0_118765, 
        HIEFFPLA_NET_0_118766, HIEFFPLA_NET_0_118767, 
        HIEFFPLA_NET_0_118768, HIEFFPLA_NET_0_118769, 
        HIEFFPLA_NET_0_118770, HIEFFPLA_NET_0_118771, 
        HIEFFPLA_NET_0_118772, HIEFFPLA_NET_0_118773, 
        HIEFFPLA_NET_0_118774, HIEFFPLA_NET_0_118775, 
        HIEFFPLA_NET_0_118776, HIEFFPLA_NET_0_118777, 
        HIEFFPLA_NET_0_118778, HIEFFPLA_NET_0_118779, 
        HIEFFPLA_NET_0_118780, HIEFFPLA_NET_0_118781, 
        HIEFFPLA_NET_0_118782, HIEFFPLA_NET_0_118783, 
        HIEFFPLA_NET_0_118784, HIEFFPLA_NET_0_118785, 
        HIEFFPLA_NET_0_118786, HIEFFPLA_NET_0_118787, 
        HIEFFPLA_NET_0_118788, HIEFFPLA_NET_0_118789, 
        HIEFFPLA_NET_0_118790, HIEFFPLA_NET_0_118791, 
        HIEFFPLA_NET_0_118792, HIEFFPLA_NET_0_118793, 
        HIEFFPLA_NET_0_118794, HIEFFPLA_NET_0_118795, 
        HIEFFPLA_NET_0_118796, HIEFFPLA_NET_0_118797, 
        HIEFFPLA_NET_0_118798, HIEFFPLA_NET_0_118799, 
        HIEFFPLA_NET_0_118800, HIEFFPLA_NET_0_118801, 
        HIEFFPLA_NET_0_118802, HIEFFPLA_NET_0_118803, 
        HIEFFPLA_NET_0_118804, HIEFFPLA_NET_0_118805, 
        HIEFFPLA_NET_0_118806, HIEFFPLA_NET_0_118807, 
        HIEFFPLA_NET_0_118808, HIEFFPLA_NET_0_118809, 
        HIEFFPLA_NET_0_118810, HIEFFPLA_NET_0_118811, 
        HIEFFPLA_NET_0_118812, HIEFFPLA_NET_0_118813, 
        HIEFFPLA_NET_0_118814, HIEFFPLA_NET_0_118815, 
        HIEFFPLA_NET_0_118816, HIEFFPLA_NET_0_118817, 
        HIEFFPLA_NET_0_118818, HIEFFPLA_NET_0_118819, 
        HIEFFPLA_NET_0_118820, HIEFFPLA_NET_0_118821, 
        HIEFFPLA_NET_0_118822, HIEFFPLA_NET_0_118823, 
        HIEFFPLA_NET_0_118824, HIEFFPLA_NET_0_118825, 
        HIEFFPLA_NET_0_118826, HIEFFPLA_NET_0_118827, 
        HIEFFPLA_NET_0_118828, HIEFFPLA_NET_0_118829, 
        HIEFFPLA_NET_0_118830, HIEFFPLA_NET_0_118831, 
        HIEFFPLA_NET_0_118832, HIEFFPLA_NET_0_118833, 
        HIEFFPLA_NET_0_118834, HIEFFPLA_NET_0_118835, 
        HIEFFPLA_NET_0_118836, HIEFFPLA_NET_0_118837, 
        HIEFFPLA_NET_0_118838, HIEFFPLA_NET_0_118839, 
        HIEFFPLA_NET_0_118840, HIEFFPLA_NET_0_118841, 
        HIEFFPLA_NET_0_118842, HIEFFPLA_NET_0_118843, 
        HIEFFPLA_NET_0_118844, HIEFFPLA_NET_0_118845, 
        HIEFFPLA_NET_0_118846, HIEFFPLA_NET_0_118847, 
        HIEFFPLA_NET_0_118848, HIEFFPLA_NET_0_118849, 
        HIEFFPLA_NET_0_118850, HIEFFPLA_NET_0_118851, 
        HIEFFPLA_NET_0_118852, HIEFFPLA_NET_0_118853, 
        HIEFFPLA_NET_0_118854, HIEFFPLA_NET_0_118855, 
        HIEFFPLA_NET_0_118856, HIEFFPLA_NET_0_118857, 
        HIEFFPLA_NET_0_118858, HIEFFPLA_NET_0_118859, 
        HIEFFPLA_NET_0_118860, HIEFFPLA_NET_0_118861, 
        HIEFFPLA_NET_0_118862, HIEFFPLA_NET_0_118863, 
        HIEFFPLA_NET_0_118864, HIEFFPLA_NET_0_118865, 
        HIEFFPLA_NET_0_118866, HIEFFPLA_NET_0_118867, 
        HIEFFPLA_NET_0_118868, HIEFFPLA_NET_0_118869, 
        HIEFFPLA_NET_0_118870, HIEFFPLA_NET_0_118871, 
        HIEFFPLA_NET_0_118872, HIEFFPLA_NET_0_118873, 
        HIEFFPLA_NET_0_118874, HIEFFPLA_NET_0_118875, 
        HIEFFPLA_NET_0_118876, HIEFFPLA_NET_0_118877, 
        HIEFFPLA_NET_0_118878, HIEFFPLA_NET_0_118879, 
        HIEFFPLA_NET_0_118880, HIEFFPLA_NET_0_118881, 
        HIEFFPLA_NET_0_118882, HIEFFPLA_NET_0_118883, 
        HIEFFPLA_NET_0_118884, HIEFFPLA_NET_0_118885, 
        HIEFFPLA_NET_0_118886, HIEFFPLA_NET_0_118887, 
        HIEFFPLA_NET_0_118888, HIEFFPLA_NET_0_118889, 
        HIEFFPLA_NET_0_118890, HIEFFPLA_NET_0_118891, 
        HIEFFPLA_NET_0_118892, HIEFFPLA_NET_0_118893, 
        HIEFFPLA_NET_0_118894, HIEFFPLA_NET_0_118895, 
        HIEFFPLA_NET_0_118896, HIEFFPLA_NET_0_118897, 
        HIEFFPLA_NET_0_118898, HIEFFPLA_NET_0_118899, 
        HIEFFPLA_NET_0_118900, HIEFFPLA_NET_0_118901, 
        HIEFFPLA_NET_0_118902, HIEFFPLA_NET_0_118903, 
        HIEFFPLA_NET_0_118904, HIEFFPLA_NET_0_118905, 
        HIEFFPLA_NET_0_118906, HIEFFPLA_NET_0_118907, 
        HIEFFPLA_NET_0_118908, HIEFFPLA_NET_0_118909, 
        HIEFFPLA_NET_0_118910, HIEFFPLA_NET_0_118911, 
        HIEFFPLA_NET_0_118912, HIEFFPLA_NET_0_118913, 
        HIEFFPLA_NET_0_118914, HIEFFPLA_NET_0_118915, 
        HIEFFPLA_NET_0_118916, HIEFFPLA_NET_0_118917, 
        HIEFFPLA_NET_0_118918, HIEFFPLA_NET_0_118919, 
        HIEFFPLA_NET_0_118920, HIEFFPLA_NET_0_118921, 
        HIEFFPLA_NET_0_118922, HIEFFPLA_NET_0_118923, 
        HIEFFPLA_NET_0_118924, HIEFFPLA_NET_0_118925, 
        HIEFFPLA_NET_0_118926, HIEFFPLA_NET_0_118927, 
        HIEFFPLA_NET_0_118928, HIEFFPLA_NET_0_118929, 
        HIEFFPLA_NET_0_118930, HIEFFPLA_NET_0_118931, 
        HIEFFPLA_NET_0_118932, HIEFFPLA_NET_0_118933, 
        HIEFFPLA_NET_0_118934, HIEFFPLA_NET_0_118935, 
        HIEFFPLA_NET_0_118936, HIEFFPLA_NET_0_118937, 
        HIEFFPLA_NET_0_118938, HIEFFPLA_NET_0_118939, 
        HIEFFPLA_NET_0_118940, HIEFFPLA_NET_0_118941, 
        HIEFFPLA_NET_0_118942, HIEFFPLA_NET_0_118943, 
        HIEFFPLA_NET_0_118944, HIEFFPLA_NET_0_118945, 
        HIEFFPLA_NET_0_118946, HIEFFPLA_NET_0_118947, 
        HIEFFPLA_NET_0_118948, HIEFFPLA_NET_0_118949, 
        HIEFFPLA_NET_0_118950, HIEFFPLA_NET_0_118951, 
        HIEFFPLA_NET_0_118952, HIEFFPLA_NET_0_118953, 
        HIEFFPLA_NET_0_118954, HIEFFPLA_NET_0_118955, 
        HIEFFPLA_NET_0_118956, HIEFFPLA_NET_0_118957, 
        HIEFFPLA_NET_0_118958, HIEFFPLA_NET_0_118959, 
        HIEFFPLA_NET_0_118960, HIEFFPLA_NET_0_118961, 
        HIEFFPLA_NET_0_118962, HIEFFPLA_NET_0_118963, 
        HIEFFPLA_NET_0_118964, HIEFFPLA_NET_0_118965, 
        HIEFFPLA_NET_0_118966, HIEFFPLA_NET_0_118967, 
        HIEFFPLA_NET_0_118968, HIEFFPLA_NET_0_118969, 
        HIEFFPLA_NET_0_118970, HIEFFPLA_NET_0_118971, 
        HIEFFPLA_NET_0_118972, HIEFFPLA_NET_0_118973, 
        HIEFFPLA_NET_0_118974, HIEFFPLA_NET_0_118975, 
        HIEFFPLA_NET_0_118976, HIEFFPLA_NET_0_118977, 
        HIEFFPLA_NET_0_118978, HIEFFPLA_NET_0_118979, 
        HIEFFPLA_NET_0_118980, HIEFFPLA_NET_0_118981, 
        HIEFFPLA_NET_0_118982, HIEFFPLA_NET_0_118983, 
        HIEFFPLA_NET_0_118984, HIEFFPLA_NET_0_118985, 
        HIEFFPLA_NET_0_118986, HIEFFPLA_NET_0_118987, 
        HIEFFPLA_NET_0_118988, HIEFFPLA_NET_0_118989, 
        HIEFFPLA_NET_0_118990, HIEFFPLA_NET_0_118991, 
        HIEFFPLA_NET_0_118992, HIEFFPLA_NET_0_118993, 
        HIEFFPLA_NET_0_118994, HIEFFPLA_NET_0_118995, 
        HIEFFPLA_NET_0_118996, HIEFFPLA_NET_0_118997, 
        HIEFFPLA_NET_0_118998, HIEFFPLA_NET_0_118999, 
        HIEFFPLA_NET_0_119000, HIEFFPLA_NET_0_119001, 
        HIEFFPLA_NET_0_119002, HIEFFPLA_NET_0_119003, 
        HIEFFPLA_NET_0_119004, HIEFFPLA_NET_0_119005, 
        HIEFFPLA_NET_0_119006, HIEFFPLA_NET_0_119007, 
        HIEFFPLA_NET_0_119008, HIEFFPLA_NET_0_119009, 
        HIEFFPLA_NET_0_119010, HIEFFPLA_NET_0_119011, 
        HIEFFPLA_NET_0_119012, HIEFFPLA_NET_0_119013, 
        HIEFFPLA_NET_0_119014, HIEFFPLA_NET_0_119015, 
        HIEFFPLA_NET_0_119016, HIEFFPLA_NET_0_119017, 
        HIEFFPLA_NET_0_119018, HIEFFPLA_NET_0_119019, 
        HIEFFPLA_NET_0_119020, HIEFFPLA_NET_0_119021, 
        HIEFFPLA_NET_0_119022, HIEFFPLA_NET_0_119023, 
        HIEFFPLA_NET_0_119024, HIEFFPLA_NET_0_119025, 
        HIEFFPLA_NET_0_119026, HIEFFPLA_NET_0_119027, 
        HIEFFPLA_NET_0_119028, HIEFFPLA_NET_0_119029, 
        HIEFFPLA_NET_0_119030, HIEFFPLA_NET_0_119031, 
        HIEFFPLA_NET_0_119032, HIEFFPLA_NET_0_119033, 
        HIEFFPLA_NET_0_119034, HIEFFPLA_NET_0_119035, 
        HIEFFPLA_NET_0_119036, HIEFFPLA_NET_0_119037, 
        HIEFFPLA_NET_0_119038, HIEFFPLA_NET_0_119039, 
        HIEFFPLA_NET_0_119040, HIEFFPLA_NET_0_119041, 
        HIEFFPLA_NET_0_119042, HIEFFPLA_NET_0_119043, 
        HIEFFPLA_NET_0_119044, HIEFFPLA_NET_0_119045, 
        HIEFFPLA_NET_0_119046, HIEFFPLA_NET_0_119047, 
        HIEFFPLA_NET_0_119048, HIEFFPLA_NET_0_119049, 
        HIEFFPLA_NET_0_119050, HIEFFPLA_NET_0_119051, 
        HIEFFPLA_NET_0_119052, HIEFFPLA_NET_0_119053, 
        HIEFFPLA_NET_0_119054, HIEFFPLA_NET_0_119055, 
        HIEFFPLA_NET_0_119056, HIEFFPLA_NET_0_119057, 
        HIEFFPLA_NET_0_119058, HIEFFPLA_NET_0_119059, 
        HIEFFPLA_NET_0_119060, HIEFFPLA_NET_0_119061, 
        HIEFFPLA_NET_0_119062, HIEFFPLA_NET_0_119063, 
        HIEFFPLA_NET_0_119064, HIEFFPLA_NET_0_119065, 
        HIEFFPLA_NET_0_119066, HIEFFPLA_NET_0_119067, 
        HIEFFPLA_NET_0_119068, HIEFFPLA_NET_0_119069, 
        HIEFFPLA_NET_0_119070, HIEFFPLA_NET_0_119071, 
        HIEFFPLA_NET_0_119072, HIEFFPLA_NET_0_119073, 
        HIEFFPLA_NET_0_119074, HIEFFPLA_NET_0_119075, 
        HIEFFPLA_NET_0_119076, HIEFFPLA_NET_0_119077, 
        HIEFFPLA_NET_0_119078, HIEFFPLA_NET_0_119079, 
        HIEFFPLA_NET_0_119080, HIEFFPLA_NET_0_119081, 
        HIEFFPLA_NET_0_119082, HIEFFPLA_NET_0_119083, 
        HIEFFPLA_NET_0_119084, HIEFFPLA_NET_0_119085, 
        HIEFFPLA_NET_0_119086, HIEFFPLA_NET_0_119087, 
        HIEFFPLA_NET_0_119088, HIEFFPLA_NET_0_119089, 
        HIEFFPLA_NET_0_119090, HIEFFPLA_NET_0_119091, 
        HIEFFPLA_NET_0_119092, HIEFFPLA_NET_0_119093, 
        HIEFFPLA_NET_0_119094, HIEFFPLA_NET_0_119095, 
        HIEFFPLA_NET_0_119096, HIEFFPLA_NET_0_119097, 
        HIEFFPLA_NET_0_119098, HIEFFPLA_NET_0_119099, 
        HIEFFPLA_NET_0_119100, HIEFFPLA_NET_0_119101, 
        HIEFFPLA_NET_0_119102, HIEFFPLA_NET_0_119103, 
        HIEFFPLA_NET_0_119104, HIEFFPLA_NET_0_119105, 
        HIEFFPLA_NET_0_119106, HIEFFPLA_NET_0_119107, 
        HIEFFPLA_NET_0_119108, HIEFFPLA_NET_0_119109, 
        HIEFFPLA_NET_0_119110, HIEFFPLA_NET_0_119111, 
        HIEFFPLA_NET_0_119112, HIEFFPLA_NET_0_119113, 
        HIEFFPLA_NET_0_119114, HIEFFPLA_NET_0_119115, 
        HIEFFPLA_NET_0_119116, HIEFFPLA_NET_0_119117, 
        HIEFFPLA_NET_0_119118, HIEFFPLA_NET_0_119119, 
        HIEFFPLA_NET_0_119120, HIEFFPLA_NET_0_119121, 
        HIEFFPLA_NET_0_119122, HIEFFPLA_NET_0_119123, 
        HIEFFPLA_NET_0_119124, HIEFFPLA_NET_0_119125, 
        HIEFFPLA_NET_0_119126, HIEFFPLA_NET_0_119127, 
        HIEFFPLA_NET_0_119128, HIEFFPLA_NET_0_119129, 
        HIEFFPLA_NET_0_119130, HIEFFPLA_NET_0_119131, 
        HIEFFPLA_NET_0_119132, HIEFFPLA_NET_0_119133, 
        HIEFFPLA_NET_0_119134, HIEFFPLA_NET_0_119135, 
        HIEFFPLA_NET_0_119136, HIEFFPLA_NET_0_119137, 
        HIEFFPLA_NET_0_119138, HIEFFPLA_NET_0_119139, 
        HIEFFPLA_NET_0_119140, HIEFFPLA_NET_0_119141, 
        HIEFFPLA_NET_0_119142, HIEFFPLA_NET_0_119143, 
        HIEFFPLA_NET_0_119144, HIEFFPLA_NET_0_119145, 
        HIEFFPLA_NET_0_119146, HIEFFPLA_NET_0_119147, 
        HIEFFPLA_NET_0_119148, HIEFFPLA_NET_0_119149, 
        HIEFFPLA_NET_0_119150, HIEFFPLA_NET_0_119151, 
        HIEFFPLA_NET_0_119152, HIEFFPLA_NET_0_119153, 
        HIEFFPLA_NET_0_119154, HIEFFPLA_NET_0_119155, 
        HIEFFPLA_NET_0_119156, HIEFFPLA_NET_0_119157, 
        HIEFFPLA_NET_0_119158, HIEFFPLA_NET_0_119159, 
        HIEFFPLA_NET_0_119160, HIEFFPLA_NET_0_119161, 
        HIEFFPLA_NET_0_119162, HIEFFPLA_NET_0_119163, 
        HIEFFPLA_NET_0_119164, HIEFFPLA_NET_0_119165, 
        HIEFFPLA_NET_0_119166, HIEFFPLA_NET_0_119167, 
        HIEFFPLA_NET_0_119168, HIEFFPLA_NET_0_119169, 
        HIEFFPLA_NET_0_119170, HIEFFPLA_NET_0_119171, 
        HIEFFPLA_NET_0_119172, HIEFFPLA_NET_0_119173, 
        HIEFFPLA_NET_0_119174, HIEFFPLA_NET_0_119175, 
        HIEFFPLA_NET_0_119176, HIEFFPLA_NET_0_119177, 
        HIEFFPLA_NET_0_119178, HIEFFPLA_NET_0_119179, 
        HIEFFPLA_NET_0_119180, HIEFFPLA_NET_0_119181, 
        HIEFFPLA_NET_0_119182, HIEFFPLA_NET_0_119183, 
        HIEFFPLA_NET_0_119184, HIEFFPLA_NET_0_119185, 
        HIEFFPLA_NET_0_119186, HIEFFPLA_NET_0_119187, 
        HIEFFPLA_NET_0_119188, HIEFFPLA_NET_0_119189, 
        HIEFFPLA_NET_0_119190, HIEFFPLA_NET_0_119191, 
        HIEFFPLA_NET_0_119192, HIEFFPLA_NET_0_119193, 
        HIEFFPLA_NET_0_119194, HIEFFPLA_NET_0_119195, 
        HIEFFPLA_NET_0_119196, HIEFFPLA_NET_0_119197, 
        HIEFFPLA_NET_0_119198, HIEFFPLA_NET_0_119199, 
        HIEFFPLA_NET_0_119200, HIEFFPLA_NET_0_119201, 
        HIEFFPLA_NET_0_119202, HIEFFPLA_NET_0_119203, 
        HIEFFPLA_NET_0_119204, HIEFFPLA_NET_0_119205, 
        HIEFFPLA_NET_0_119206, HIEFFPLA_NET_0_119207, 
        HIEFFPLA_NET_0_119208, HIEFFPLA_NET_0_119209, 
        HIEFFPLA_NET_0_119210, HIEFFPLA_NET_0_119211, 
        HIEFFPLA_NET_0_119212, HIEFFPLA_NET_0_119213, 
        HIEFFPLA_NET_0_119214, HIEFFPLA_NET_0_119215, 
        HIEFFPLA_NET_0_119216, HIEFFPLA_NET_0_119217, 
        HIEFFPLA_NET_0_119218, HIEFFPLA_NET_0_119219, 
        HIEFFPLA_NET_0_119220, HIEFFPLA_NET_0_119221, 
        HIEFFPLA_NET_0_119222, HIEFFPLA_NET_0_119223, 
        HIEFFPLA_NET_0_119224, HIEFFPLA_NET_0_119225, 
        HIEFFPLA_NET_0_119226, HIEFFPLA_NET_0_119227, 
        HIEFFPLA_NET_0_119228, HIEFFPLA_NET_0_119229, 
        HIEFFPLA_NET_0_119230, HIEFFPLA_NET_0_119231, 
        HIEFFPLA_NET_0_119232, HIEFFPLA_NET_0_119233, 
        HIEFFPLA_NET_0_119234, HIEFFPLA_NET_0_119235, 
        HIEFFPLA_NET_0_119236, HIEFFPLA_NET_0_119237, 
        HIEFFPLA_NET_0_119238, HIEFFPLA_NET_0_119239, 
        HIEFFPLA_NET_0_119240, HIEFFPLA_NET_0_119241, 
        HIEFFPLA_NET_0_119242, HIEFFPLA_NET_0_119243, 
        HIEFFPLA_NET_0_119244, HIEFFPLA_NET_0_119245, 
        HIEFFPLA_NET_0_119246, HIEFFPLA_NET_0_119247, 
        HIEFFPLA_NET_0_119248, HIEFFPLA_NET_0_119249, 
        HIEFFPLA_NET_0_119250, HIEFFPLA_NET_0_119251, 
        HIEFFPLA_NET_0_119252, HIEFFPLA_NET_0_119253, 
        HIEFFPLA_NET_0_119254, HIEFFPLA_NET_0_119255, 
        HIEFFPLA_NET_0_119256, HIEFFPLA_NET_0_119257, 
        HIEFFPLA_NET_0_119258, HIEFFPLA_NET_0_119259, 
        HIEFFPLA_NET_0_119260, HIEFFPLA_NET_0_119261, 
        HIEFFPLA_NET_0_119262, HIEFFPLA_NET_0_119263, 
        HIEFFPLA_NET_0_119264, HIEFFPLA_NET_0_119265, 
        HIEFFPLA_NET_0_119266, HIEFFPLA_NET_0_119267, 
        HIEFFPLA_NET_0_119268, HIEFFPLA_NET_0_119269, 
        HIEFFPLA_NET_0_119270, HIEFFPLA_NET_0_119271, 
        HIEFFPLA_NET_0_119272, HIEFFPLA_NET_0_119273, 
        HIEFFPLA_NET_0_119274, HIEFFPLA_NET_0_119275, 
        HIEFFPLA_NET_0_119276, HIEFFPLA_NET_0_119277, 
        HIEFFPLA_NET_0_119278, HIEFFPLA_NET_0_119279, 
        HIEFFPLA_NET_0_119280, HIEFFPLA_NET_0_119281, 
        HIEFFPLA_NET_0_119282, HIEFFPLA_NET_0_119283, 
        HIEFFPLA_NET_0_119284, HIEFFPLA_NET_0_119285, 
        HIEFFPLA_NET_0_119286, HIEFFPLA_NET_0_119287, 
        HIEFFPLA_NET_0_119288, HIEFFPLA_NET_0_119289, 
        HIEFFPLA_NET_0_119290, HIEFFPLA_NET_0_119291, 
        HIEFFPLA_NET_0_119292, HIEFFPLA_NET_0_119293, 
        HIEFFPLA_NET_0_119294, HIEFFPLA_NET_0_119295, 
        HIEFFPLA_NET_0_119296, HIEFFPLA_NET_0_119297, 
        HIEFFPLA_NET_0_119298, HIEFFPLA_NET_0_119299, 
        HIEFFPLA_NET_0_119300, HIEFFPLA_NET_0_119301, 
        HIEFFPLA_NET_0_119302, HIEFFPLA_NET_0_119303, 
        HIEFFPLA_NET_0_119304, HIEFFPLA_NET_0_119305, 
        HIEFFPLA_NET_0_119306, HIEFFPLA_NET_0_119307, 
        HIEFFPLA_NET_0_119308, HIEFFPLA_NET_0_119309, 
        HIEFFPLA_NET_0_119310, HIEFFPLA_NET_0_119311, 
        HIEFFPLA_NET_0_119312, HIEFFPLA_NET_0_119313, 
        HIEFFPLA_NET_0_119314, HIEFFPLA_NET_0_119315, 
        HIEFFPLA_NET_0_119316, HIEFFPLA_NET_0_119317, 
        HIEFFPLA_NET_0_119318, HIEFFPLA_NET_0_119319, 
        HIEFFPLA_NET_0_119320, HIEFFPLA_NET_0_119321, 
        HIEFFPLA_NET_0_119322, HIEFFPLA_NET_0_119323, 
        HIEFFPLA_NET_0_119324, HIEFFPLA_NET_0_119325, 
        HIEFFPLA_NET_0_119326, HIEFFPLA_NET_0_119327, 
        HIEFFPLA_NET_0_119328, HIEFFPLA_NET_0_119329, 
        HIEFFPLA_NET_0_119330, HIEFFPLA_NET_0_119331, 
        HIEFFPLA_NET_0_119332, HIEFFPLA_NET_0_119333, 
        HIEFFPLA_NET_0_119334, HIEFFPLA_NET_0_119335, 
        HIEFFPLA_NET_0_119336, HIEFFPLA_NET_0_119337, 
        HIEFFPLA_NET_0_119338, HIEFFPLA_NET_0_119339, 
        HIEFFPLA_NET_0_119340, HIEFFPLA_NET_0_119341, 
        HIEFFPLA_NET_0_119342, HIEFFPLA_NET_0_119343, 
        HIEFFPLA_NET_0_119344, HIEFFPLA_NET_0_119345, 
        HIEFFPLA_NET_0_119346, HIEFFPLA_NET_0_119347, 
        HIEFFPLA_NET_0_119348, HIEFFPLA_NET_0_119349, 
        HIEFFPLA_NET_0_119350, HIEFFPLA_NET_0_119351, 
        HIEFFPLA_NET_0_119352, HIEFFPLA_NET_0_119353, 
        HIEFFPLA_NET_0_119354, HIEFFPLA_NET_0_119355, 
        HIEFFPLA_NET_0_119356, HIEFFPLA_NET_0_119357, 
        HIEFFPLA_NET_0_119358, HIEFFPLA_NET_0_119359, 
        HIEFFPLA_NET_0_119360, HIEFFPLA_NET_0_119361, 
        HIEFFPLA_NET_0_119362, HIEFFPLA_NET_0_119363, 
        HIEFFPLA_NET_0_119364, HIEFFPLA_NET_0_119365, 
        HIEFFPLA_NET_0_119366, HIEFFPLA_NET_0_119367, 
        HIEFFPLA_NET_0_119368, HIEFFPLA_NET_0_119369, 
        HIEFFPLA_NET_0_119370, HIEFFPLA_NET_0_119371, 
        HIEFFPLA_NET_0_119372, HIEFFPLA_NET_0_119373, 
        HIEFFPLA_NET_0_119374, HIEFFPLA_NET_0_119375, 
        HIEFFPLA_NET_0_119376, HIEFFPLA_NET_0_119377, 
        HIEFFPLA_NET_0_119378, HIEFFPLA_NET_0_119379, 
        HIEFFPLA_NET_0_119380, HIEFFPLA_NET_0_119381, 
        HIEFFPLA_NET_0_119382, HIEFFPLA_NET_0_119383, 
        HIEFFPLA_NET_0_119384, HIEFFPLA_NET_0_119385, 
        HIEFFPLA_NET_0_119386, HIEFFPLA_NET_0_119387, 
        HIEFFPLA_NET_0_119388, HIEFFPLA_NET_0_119389, 
        HIEFFPLA_NET_0_119390, HIEFFPLA_NET_0_119391, 
        HIEFFPLA_NET_0_119392, HIEFFPLA_NET_0_119393, 
        HIEFFPLA_NET_0_119394, HIEFFPLA_NET_0_119395, 
        HIEFFPLA_NET_0_119396, HIEFFPLA_NET_0_119397, 
        HIEFFPLA_NET_0_119398, HIEFFPLA_NET_0_119399, 
        HIEFFPLA_NET_0_119400, HIEFFPLA_NET_0_119401, 
        HIEFFPLA_NET_0_119402, HIEFFPLA_NET_0_119403, 
        HIEFFPLA_NET_0_119404, HIEFFPLA_NET_0_119405, 
        HIEFFPLA_NET_0_119406, HIEFFPLA_NET_0_119407, 
        HIEFFPLA_NET_0_119408, HIEFFPLA_NET_0_119409, 
        HIEFFPLA_NET_0_119410, HIEFFPLA_NET_0_119411, 
        HIEFFPLA_NET_0_119412, HIEFFPLA_NET_0_119413, 
        HIEFFPLA_NET_0_119414, HIEFFPLA_NET_0_119415, 
        HIEFFPLA_NET_0_119416, HIEFFPLA_NET_0_119417, 
        HIEFFPLA_NET_0_119418, HIEFFPLA_NET_0_119419, 
        HIEFFPLA_NET_0_119420, HIEFFPLA_NET_0_119421, 
        HIEFFPLA_NET_0_119422, HIEFFPLA_NET_0_119423, 
        HIEFFPLA_NET_0_119424, HIEFFPLA_NET_0_119425, 
        HIEFFPLA_NET_0_119426, HIEFFPLA_NET_0_119427, 
        HIEFFPLA_NET_0_119428, HIEFFPLA_NET_0_119429, 
        HIEFFPLA_NET_0_119430, HIEFFPLA_NET_0_119431, 
        HIEFFPLA_NET_0_119432, HIEFFPLA_NET_0_119433, 
        HIEFFPLA_NET_0_119434, HIEFFPLA_NET_0_119435, 
        HIEFFPLA_NET_0_119436, HIEFFPLA_NET_0_119437, 
        HIEFFPLA_NET_0_119438, HIEFFPLA_NET_0_119439, 
        HIEFFPLA_NET_0_119440, HIEFFPLA_NET_0_119441, 
        HIEFFPLA_NET_0_119442, HIEFFPLA_NET_0_119443, 
        HIEFFPLA_NET_0_119444, HIEFFPLA_NET_0_119445, 
        HIEFFPLA_NET_0_119446, HIEFFPLA_NET_0_119447, 
        HIEFFPLA_NET_0_119448, HIEFFPLA_NET_0_119449, 
        HIEFFPLA_NET_0_119450, HIEFFPLA_NET_0_119451, 
        HIEFFPLA_NET_0_119452, HIEFFPLA_NET_0_119453, 
        HIEFFPLA_NET_0_119454, HIEFFPLA_NET_0_119455, 
        HIEFFPLA_NET_0_119456, HIEFFPLA_NET_0_119457, 
        HIEFFPLA_NET_0_119458, HIEFFPLA_NET_0_119459, 
        HIEFFPLA_NET_0_119460, HIEFFPLA_NET_0_119461, 
        HIEFFPLA_NET_0_119462, HIEFFPLA_NET_0_119463, 
        HIEFFPLA_NET_0_119464, HIEFFPLA_NET_0_119465, 
        HIEFFPLA_NET_0_119466, HIEFFPLA_NET_0_119467, 
        HIEFFPLA_NET_0_119468, HIEFFPLA_NET_0_119469, 
        HIEFFPLA_NET_0_119470, HIEFFPLA_NET_0_119471, 
        HIEFFPLA_NET_0_119472, HIEFFPLA_NET_0_119473, 
        HIEFFPLA_NET_0_119474, HIEFFPLA_NET_0_119475, 
        HIEFFPLA_NET_0_119476, HIEFFPLA_NET_0_119477, 
        HIEFFPLA_NET_0_119478, HIEFFPLA_NET_0_119479, 
        HIEFFPLA_NET_0_119480, HIEFFPLA_NET_0_119481, 
        HIEFFPLA_NET_0_119482, HIEFFPLA_NET_0_119483, 
        HIEFFPLA_NET_0_119484, HIEFFPLA_NET_0_119485, 
        HIEFFPLA_NET_0_119486, HIEFFPLA_NET_0_119487, 
        HIEFFPLA_NET_0_119488, HIEFFPLA_NET_0_119489, 
        HIEFFPLA_NET_0_119490, HIEFFPLA_NET_0_119491, 
        HIEFFPLA_NET_0_119492, HIEFFPLA_NET_0_119493, 
        HIEFFPLA_NET_0_119494, HIEFFPLA_NET_0_119495, 
        HIEFFPLA_NET_0_119496, HIEFFPLA_NET_0_119497, 
        HIEFFPLA_NET_0_119498, HIEFFPLA_NET_0_119499, 
        HIEFFPLA_NET_0_119500, HIEFFPLA_NET_0_119501, 
        HIEFFPLA_NET_0_119502, HIEFFPLA_NET_0_119503, 
        HIEFFPLA_NET_0_119504, HIEFFPLA_NET_0_119505, 
        HIEFFPLA_NET_0_119506, HIEFFPLA_NET_0_119507, 
        HIEFFPLA_NET_0_119508, HIEFFPLA_NET_0_119509, 
        HIEFFPLA_NET_0_119510, HIEFFPLA_NET_0_119511, 
        HIEFFPLA_NET_0_119512, HIEFFPLA_NET_0_119513, 
        HIEFFPLA_NET_0_119514, HIEFFPLA_NET_0_119515, 
        HIEFFPLA_NET_0_119516, HIEFFPLA_NET_0_119517, 
        HIEFFPLA_NET_0_119518, HIEFFPLA_NET_0_119519, 
        HIEFFPLA_NET_0_119520, HIEFFPLA_NET_0_119521, 
        HIEFFPLA_NET_0_119522, HIEFFPLA_NET_0_119523, 
        HIEFFPLA_NET_0_119524, HIEFFPLA_NET_0_119525, 
        HIEFFPLA_NET_0_119526, HIEFFPLA_NET_0_119527, 
        HIEFFPLA_NET_0_119528, HIEFFPLA_NET_0_119529, 
        HIEFFPLA_NET_0_119530, HIEFFPLA_NET_0_119531, 
        HIEFFPLA_NET_0_119532, HIEFFPLA_NET_0_119533, 
        HIEFFPLA_NET_0_119534, HIEFFPLA_NET_0_119535, 
        HIEFFPLA_NET_0_119536, HIEFFPLA_NET_0_119537, 
        HIEFFPLA_NET_0_119538, HIEFFPLA_NET_0_119539, 
        HIEFFPLA_NET_0_119540, HIEFFPLA_NET_0_119541, 
        HIEFFPLA_NET_0_119542, HIEFFPLA_NET_0_119543, 
        HIEFFPLA_NET_0_119544, HIEFFPLA_NET_0_119545, 
        HIEFFPLA_NET_0_119546, HIEFFPLA_NET_0_119547, 
        HIEFFPLA_NET_0_119548, HIEFFPLA_NET_0_119549, 
        HIEFFPLA_NET_0_119550, HIEFFPLA_NET_0_119551, 
        HIEFFPLA_NET_0_119552, HIEFFPLA_NET_0_119553, 
        HIEFFPLA_NET_0_119554, HIEFFPLA_NET_0_119555, 
        HIEFFPLA_NET_0_119556, HIEFFPLA_NET_0_119557, 
        HIEFFPLA_NET_0_119558, HIEFFPLA_NET_0_119559, 
        HIEFFPLA_NET_0_119560, HIEFFPLA_NET_0_119561, 
        HIEFFPLA_NET_0_119562, HIEFFPLA_NET_0_119563, 
        HIEFFPLA_NET_0_119564, HIEFFPLA_NET_0_119565, 
        HIEFFPLA_NET_0_119566, HIEFFPLA_NET_0_119567, 
        HIEFFPLA_NET_0_119568, HIEFFPLA_NET_0_119569, 
        HIEFFPLA_NET_0_119570, HIEFFPLA_NET_0_119571, 
        HIEFFPLA_NET_0_119572, HIEFFPLA_NET_0_119573, 
        HIEFFPLA_NET_0_119574, HIEFFPLA_NET_0_119575, 
        HIEFFPLA_NET_0_119576, HIEFFPLA_NET_0_119577, 
        HIEFFPLA_NET_0_119578, HIEFFPLA_NET_0_119579, 
        HIEFFPLA_NET_0_119580, HIEFFPLA_NET_0_119581, 
        HIEFFPLA_NET_0_119582, HIEFFPLA_NET_0_119583, 
        HIEFFPLA_NET_0_119584, HIEFFPLA_NET_0_119585, 
        HIEFFPLA_NET_0_119586, HIEFFPLA_NET_0_119587, 
        HIEFFPLA_NET_0_119588, HIEFFPLA_NET_0_119589, 
        HIEFFPLA_NET_0_119590, HIEFFPLA_NET_0_119591, 
        HIEFFPLA_NET_0_119592, HIEFFPLA_NET_0_119593, 
        HIEFFPLA_NET_0_119594, HIEFFPLA_NET_0_119595, 
        HIEFFPLA_NET_0_119596, HIEFFPLA_NET_0_119597, 
        HIEFFPLA_NET_0_119598, HIEFFPLA_NET_0_119599, 
        HIEFFPLA_NET_0_119600, HIEFFPLA_NET_0_119601, 
        HIEFFPLA_NET_0_119602, HIEFFPLA_NET_0_119603, 
        HIEFFPLA_NET_0_119604, HIEFFPLA_NET_0_119605, 
        HIEFFPLA_NET_0_119606, HIEFFPLA_NET_0_119607, 
        HIEFFPLA_NET_0_119608, HIEFFPLA_NET_0_119609, 
        HIEFFPLA_NET_0_119610, HIEFFPLA_NET_0_119611, 
        HIEFFPLA_NET_0_119612, HIEFFPLA_NET_0_119613, 
        HIEFFPLA_NET_0_119614, HIEFFPLA_NET_0_119615, 
        HIEFFPLA_NET_0_119616, HIEFFPLA_NET_0_119617, 
        HIEFFPLA_NET_0_119618, HIEFFPLA_NET_0_119619, 
        HIEFFPLA_NET_0_119620, HIEFFPLA_NET_0_119621, 
        HIEFFPLA_NET_0_119622, HIEFFPLA_NET_0_119623, 
        HIEFFPLA_NET_0_119624, HIEFFPLA_NET_0_119625, 
        HIEFFPLA_NET_0_119626, HIEFFPLA_NET_0_119627, 
        HIEFFPLA_NET_0_119628, HIEFFPLA_NET_0_119629, 
        HIEFFPLA_NET_0_119630, HIEFFPLA_NET_0_119631, 
        HIEFFPLA_NET_0_119632, HIEFFPLA_NET_0_119633, 
        HIEFFPLA_NET_0_119634, HIEFFPLA_NET_0_119635, 
        HIEFFPLA_NET_0_119636, HIEFFPLA_NET_0_119637, 
        HIEFFPLA_NET_0_119638, HIEFFPLA_NET_0_119639, 
        HIEFFPLA_NET_0_119640, HIEFFPLA_NET_0_119641, 
        HIEFFPLA_NET_0_119642, HIEFFPLA_NET_0_119643, 
        HIEFFPLA_NET_0_119644, HIEFFPLA_NET_0_119645, 
        HIEFFPLA_NET_0_119646, HIEFFPLA_NET_0_119647, 
        HIEFFPLA_NET_0_119648, HIEFFPLA_NET_0_119649, 
        HIEFFPLA_NET_0_119650, HIEFFPLA_NET_0_119651, 
        HIEFFPLA_NET_0_119652, HIEFFPLA_NET_0_119653, 
        HIEFFPLA_NET_0_119654, HIEFFPLA_NET_0_119655, 
        HIEFFPLA_NET_0_119656, HIEFFPLA_NET_0_119657, 
        HIEFFPLA_NET_0_119658, HIEFFPLA_NET_0_119659, 
        HIEFFPLA_NET_0_119660, HIEFFPLA_NET_0_119661, 
        HIEFFPLA_NET_0_119662, HIEFFPLA_NET_0_119663, 
        HIEFFPLA_NET_0_119664, HIEFFPLA_NET_0_119665, 
        HIEFFPLA_NET_0_119666, HIEFFPLA_NET_0_119667, 
        HIEFFPLA_NET_0_119668, HIEFFPLA_NET_0_119669, 
        HIEFFPLA_NET_0_119670, HIEFFPLA_NET_0_119671, 
        HIEFFPLA_NET_0_119672, HIEFFPLA_NET_0_119673, 
        HIEFFPLA_NET_0_119674, HIEFFPLA_NET_0_119675, 
        HIEFFPLA_NET_0_119676, HIEFFPLA_NET_0_119677, 
        HIEFFPLA_NET_0_119678, HIEFFPLA_NET_0_119679, 
        HIEFFPLA_NET_0_119680, HIEFFPLA_NET_0_119681, 
        HIEFFPLA_NET_0_119682, HIEFFPLA_NET_0_119683, 
        HIEFFPLA_NET_0_119684, HIEFFPLA_NET_0_119685, 
        HIEFFPLA_NET_0_119686, HIEFFPLA_NET_0_119687, 
        HIEFFPLA_NET_0_119688, HIEFFPLA_NET_0_119689, 
        HIEFFPLA_NET_0_119690, HIEFFPLA_NET_0_119691, 
        HIEFFPLA_NET_0_119692, HIEFFPLA_NET_0_119693, 
        HIEFFPLA_NET_0_119694, HIEFFPLA_NET_0_119695, 
        HIEFFPLA_NET_0_119696, HIEFFPLA_NET_0_119697, 
        HIEFFPLA_NET_0_119698, HIEFFPLA_NET_0_119699, 
        HIEFFPLA_NET_0_119700, HIEFFPLA_NET_0_119701, 
        HIEFFPLA_NET_0_119702, HIEFFPLA_NET_0_119703, 
        HIEFFPLA_NET_0_119704, HIEFFPLA_NET_0_119705, 
        HIEFFPLA_NET_0_119706, HIEFFPLA_NET_0_119707, 
        HIEFFPLA_NET_0_119708, HIEFFPLA_NET_0_119709, 
        HIEFFPLA_NET_0_119710, HIEFFPLA_NET_0_119711, 
        HIEFFPLA_NET_0_119712, HIEFFPLA_NET_0_119713, 
        HIEFFPLA_NET_0_119714, HIEFFPLA_NET_0_119715, 
        HIEFFPLA_NET_0_119716, HIEFFPLA_NET_0_119717, 
        HIEFFPLA_NET_0_119718, HIEFFPLA_NET_0_119719, 
        HIEFFPLA_NET_0_119720, HIEFFPLA_NET_0_119721, 
        HIEFFPLA_NET_0_119722, HIEFFPLA_NET_0_119723, 
        HIEFFPLA_NET_0_119724, HIEFFPLA_NET_0_119725, 
        HIEFFPLA_NET_0_119726, HIEFFPLA_NET_0_119727, 
        HIEFFPLA_NET_0_119728, HIEFFPLA_NET_0_119729, 
        HIEFFPLA_NET_0_119730, HIEFFPLA_NET_0_119731, 
        HIEFFPLA_NET_0_119732, HIEFFPLA_NET_0_119733, 
        HIEFFPLA_NET_0_119734, HIEFFPLA_NET_0_119735, 
        HIEFFPLA_NET_0_119736, HIEFFPLA_NET_0_119737, 
        HIEFFPLA_NET_0_119738, HIEFFPLA_NET_0_119739, 
        HIEFFPLA_NET_0_119740, HIEFFPLA_NET_0_119741, 
        HIEFFPLA_NET_0_119742, HIEFFPLA_NET_0_119743, 
        HIEFFPLA_NET_0_119744, HIEFFPLA_NET_0_119745, 
        HIEFFPLA_NET_0_119746, HIEFFPLA_NET_0_119747, 
        HIEFFPLA_NET_0_119748, HIEFFPLA_NET_0_119749, 
        HIEFFPLA_NET_0_119750, HIEFFPLA_NET_0_119751, 
        HIEFFPLA_NET_0_119752, HIEFFPLA_NET_0_119753, 
        HIEFFPLA_NET_0_119754, HIEFFPLA_NET_0_119755, 
        HIEFFPLA_NET_0_119756, HIEFFPLA_NET_0_119757, 
        HIEFFPLA_NET_0_119758, HIEFFPLA_NET_0_119759, 
        HIEFFPLA_NET_0_119760, HIEFFPLA_NET_0_119761, 
        HIEFFPLA_NET_0_119762, HIEFFPLA_NET_0_119763, 
        HIEFFPLA_NET_0_119764, HIEFFPLA_NET_0_119765, 
        HIEFFPLA_NET_0_119766, HIEFFPLA_NET_0_119767, 
        HIEFFPLA_NET_0_119768, HIEFFPLA_NET_0_119769, 
        HIEFFPLA_NET_0_119770, HIEFFPLA_NET_0_119771, 
        HIEFFPLA_NET_0_119772, HIEFFPLA_NET_0_119773, 
        HIEFFPLA_NET_0_119774, HIEFFPLA_NET_0_119775, 
        HIEFFPLA_NET_0_119776, HIEFFPLA_NET_0_119777, 
        HIEFFPLA_NET_0_119778, HIEFFPLA_NET_0_119779, 
        HIEFFPLA_NET_0_119780, HIEFFPLA_NET_0_119781, 
        HIEFFPLA_NET_0_119782, HIEFFPLA_NET_0_119783, 
        HIEFFPLA_NET_0_119784, HIEFFPLA_NET_0_119785, 
        HIEFFPLA_NET_0_119786, HIEFFPLA_NET_0_119787, 
        HIEFFPLA_NET_0_119788, HIEFFPLA_NET_0_119789, 
        HIEFFPLA_NET_0_119790, HIEFFPLA_NET_0_119791, 
        HIEFFPLA_NET_0_119792, HIEFFPLA_NET_0_119793, 
        HIEFFPLA_NET_0_119794, HIEFFPLA_NET_0_119795, 
        HIEFFPLA_NET_0_119796, HIEFFPLA_NET_0_119797, 
        HIEFFPLA_NET_0_119798, HIEFFPLA_NET_0_119799, 
        HIEFFPLA_NET_0_119800, HIEFFPLA_NET_0_119801, 
        HIEFFPLA_NET_0_119802, HIEFFPLA_NET_0_119803, 
        HIEFFPLA_NET_0_119804, HIEFFPLA_NET_0_119805, 
        HIEFFPLA_NET_0_119806, HIEFFPLA_NET_0_119807, 
        HIEFFPLA_NET_0_119808, HIEFFPLA_NET_0_119809, 
        HIEFFPLA_NET_0_119810, HIEFFPLA_NET_0_119811, 
        HIEFFPLA_NET_0_119812, HIEFFPLA_NET_0_119813, 
        HIEFFPLA_NET_0_119814, HIEFFPLA_NET_0_119815, 
        HIEFFPLA_NET_0_119816, HIEFFPLA_NET_0_119817, 
        HIEFFPLA_NET_0_119818, HIEFFPLA_NET_0_119819, 
        HIEFFPLA_NET_0_119820, HIEFFPLA_NET_0_119821, 
        HIEFFPLA_NET_0_119822, HIEFFPLA_NET_0_119823, 
        HIEFFPLA_NET_0_119824, HIEFFPLA_NET_0_119825, 
        HIEFFPLA_NET_0_119826, HIEFFPLA_NET_0_119827, 
        HIEFFPLA_NET_0_119828, HIEFFPLA_NET_0_119829, 
        HIEFFPLA_NET_0_119830, HIEFFPLA_NET_0_119831, 
        HIEFFPLA_NET_0_119832, HIEFFPLA_NET_0_119833, 
        HIEFFPLA_NET_0_119834, HIEFFPLA_NET_0_119835, 
        HIEFFPLA_NET_0_119836, HIEFFPLA_NET_0_119837, 
        HIEFFPLA_NET_0_119838, HIEFFPLA_NET_0_119839, 
        HIEFFPLA_NET_0_119840, HIEFFPLA_NET_0_119841, 
        HIEFFPLA_NET_0_119842, HIEFFPLA_NET_0_119843, 
        HIEFFPLA_NET_0_119844, HIEFFPLA_NET_0_119845, 
        HIEFFPLA_NET_0_119846, HIEFFPLA_NET_0_119847, 
        HIEFFPLA_NET_0_119848, HIEFFPLA_NET_0_119849, 
        HIEFFPLA_NET_0_119850, HIEFFPLA_NET_0_119851, 
        HIEFFPLA_NET_0_119852, HIEFFPLA_NET_0_119853, 
        HIEFFPLA_NET_0_119854, HIEFFPLA_NET_0_119855, 
        HIEFFPLA_NET_0_119856, HIEFFPLA_NET_0_119857, 
        HIEFFPLA_NET_0_119858, HIEFFPLA_NET_0_119859, 
        HIEFFPLA_NET_0_119860, HIEFFPLA_NET_0_119861, 
        HIEFFPLA_NET_0_119862, HIEFFPLA_NET_0_119863, 
        HIEFFPLA_NET_0_119864, HIEFFPLA_NET_0_119865, 
        HIEFFPLA_NET_0_119866, HIEFFPLA_NET_0_119867, 
        HIEFFPLA_NET_0_119868, HIEFFPLA_NET_0_119869, 
        HIEFFPLA_NET_0_119870, HIEFFPLA_NET_0_119871, 
        HIEFFPLA_NET_0_119872, HIEFFPLA_NET_0_119873, 
        HIEFFPLA_NET_0_119874, HIEFFPLA_NET_0_119875, 
        HIEFFPLA_NET_0_119876, HIEFFPLA_NET_0_119877, 
        HIEFFPLA_NET_0_119878, HIEFFPLA_NET_0_119879, 
        HIEFFPLA_NET_0_119880, HIEFFPLA_NET_0_119881, 
        HIEFFPLA_NET_0_119882, HIEFFPLA_NET_0_119883, 
        HIEFFPLA_NET_0_119884, HIEFFPLA_NET_0_119885, 
        HIEFFPLA_NET_0_119886, HIEFFPLA_NET_0_119887, 
        HIEFFPLA_NET_0_119888, HIEFFPLA_NET_0_119889, 
        HIEFFPLA_NET_0_119890, HIEFFPLA_NET_0_119891, 
        HIEFFPLA_NET_0_119892, HIEFFPLA_NET_0_119893, 
        HIEFFPLA_NET_0_119894, HIEFFPLA_NET_0_119895, 
        HIEFFPLA_NET_0_119896, HIEFFPLA_NET_0_119897, 
        HIEFFPLA_NET_0_119898, HIEFFPLA_NET_0_119899, 
        HIEFFPLA_NET_0_119900, HIEFFPLA_NET_0_119901, 
        HIEFFPLA_NET_0_119902, HIEFFPLA_NET_0_119903, 
        HIEFFPLA_NET_0_119904, HIEFFPLA_NET_0_119905, 
        HIEFFPLA_NET_0_119906, HIEFFPLA_NET_0_119907, 
        HIEFFPLA_NET_0_119908, HIEFFPLA_NET_0_119909, 
        HIEFFPLA_NET_0_119910, HIEFFPLA_NET_0_119911, 
        HIEFFPLA_NET_0_119912, HIEFFPLA_NET_0_119913, 
        HIEFFPLA_NET_0_119914, HIEFFPLA_NET_0_119915, 
        HIEFFPLA_NET_0_119916, HIEFFPLA_NET_0_119917, 
        HIEFFPLA_NET_0_119918, HIEFFPLA_NET_0_119919, 
        HIEFFPLA_NET_0_119920, HIEFFPLA_NET_0_119921, 
        HIEFFPLA_NET_0_119922, HIEFFPLA_NET_0_119923, 
        HIEFFPLA_NET_0_119924, HIEFFPLA_NET_0_119925, 
        HIEFFPLA_NET_0_119926, HIEFFPLA_NET_0_119927, 
        HIEFFPLA_NET_0_119928, HIEFFPLA_NET_0_119929, 
        HIEFFPLA_NET_0_119930, HIEFFPLA_NET_0_119931, 
        HIEFFPLA_NET_0_119932, HIEFFPLA_NET_0_119933, 
        HIEFFPLA_NET_0_119934, HIEFFPLA_NET_0_119935, 
        HIEFFPLA_NET_0_119936, HIEFFPLA_NET_0_119937, 
        HIEFFPLA_NET_0_119938, HIEFFPLA_NET_0_119939, 
        HIEFFPLA_NET_0_119940, HIEFFPLA_NET_0_119941, 
        HIEFFPLA_NET_0_119942, HIEFFPLA_NET_0_119943, 
        HIEFFPLA_NET_0_119944, HIEFFPLA_NET_0_119945, 
        HIEFFPLA_NET_0_119946, HIEFFPLA_NET_0_119947, 
        HIEFFPLA_NET_0_119948, HIEFFPLA_NET_0_119949, 
        HIEFFPLA_NET_0_119950, HIEFFPLA_NET_0_119951, 
        HIEFFPLA_NET_0_119952, HIEFFPLA_NET_0_119953, 
        HIEFFPLA_NET_0_119954, HIEFFPLA_NET_0_119955, 
        HIEFFPLA_NET_0_119956, HIEFFPLA_NET_0_119957, 
        HIEFFPLA_NET_0_119958, HIEFFPLA_NET_0_119959, 
        HIEFFPLA_NET_0_119960, HIEFFPLA_NET_0_119961, 
        HIEFFPLA_NET_0_119962, HIEFFPLA_NET_0_119963, 
        HIEFFPLA_NET_0_119964, HIEFFPLA_NET_0_119965, 
        HIEFFPLA_NET_0_119966, HIEFFPLA_NET_0_119967, 
        HIEFFPLA_NET_0_119968, HIEFFPLA_NET_0_119969, 
        HIEFFPLA_NET_0_119970, HIEFFPLA_NET_0_119971, 
        HIEFFPLA_NET_0_119972, HIEFFPLA_NET_0_119973, 
        HIEFFPLA_NET_0_119974, HIEFFPLA_NET_0_119975, 
        HIEFFPLA_NET_0_119976, HIEFFPLA_NET_0_119977, 
        HIEFFPLA_NET_0_119978, HIEFFPLA_NET_0_119979, 
        HIEFFPLA_NET_0_119980, HIEFFPLA_NET_0_119981, 
        HIEFFPLA_NET_0_119982, HIEFFPLA_NET_0_119983, 
        HIEFFPLA_NET_0_119984, HIEFFPLA_NET_0_119985, 
        HIEFFPLA_NET_0_119986, HIEFFPLA_NET_0_119987, 
        HIEFFPLA_NET_0_119988, HIEFFPLA_NET_0_119989, 
        HIEFFPLA_NET_0_119990, HIEFFPLA_NET_0_119991, 
        HIEFFPLA_NET_0_119992, HIEFFPLA_NET_0_119993, 
        HIEFFPLA_NET_0_119994, HIEFFPLA_NET_0_119995, 
        HIEFFPLA_NET_0_119996, HIEFFPLA_NET_0_119997, 
        HIEFFPLA_NET_0_119998, HIEFFPLA_NET_0_119999, 
        HIEFFPLA_NET_0_120000, HIEFFPLA_NET_0_120001, 
        HIEFFPLA_NET_0_120002, HIEFFPLA_NET_0_120003, 
        HIEFFPLA_NET_0_120004, HIEFFPLA_NET_0_120005, 
        HIEFFPLA_NET_0_120006, HIEFFPLA_NET_0_120007, 
        HIEFFPLA_NET_0_120008, HIEFFPLA_NET_0_120009, 
        HIEFFPLA_NET_0_120010, HIEFFPLA_NET_0_120011, 
        HIEFFPLA_NET_0_120012, HIEFFPLA_NET_0_120013, 
        HIEFFPLA_NET_0_120014, HIEFFPLA_NET_0_120015, 
        HIEFFPLA_NET_0_120016, HIEFFPLA_NET_0_120017, 
        HIEFFPLA_NET_0_120018, HIEFFPLA_NET_0_120019, 
        HIEFFPLA_NET_0_120020, HIEFFPLA_NET_0_120021, 
        HIEFFPLA_NET_0_120022, HIEFFPLA_NET_0_120023, 
        HIEFFPLA_NET_0_120024, HIEFFPLA_NET_0_120025, 
        HIEFFPLA_NET_0_120026, HIEFFPLA_NET_0_120027, 
        HIEFFPLA_NET_0_120028, HIEFFPLA_NET_0_120029, 
        HIEFFPLA_NET_0_120030, HIEFFPLA_NET_0_120031, 
        HIEFFPLA_NET_0_120032, HIEFFPLA_NET_0_120033, 
        HIEFFPLA_NET_0_120034, HIEFFPLA_NET_0_120035, 
        HIEFFPLA_NET_0_120036, HIEFFPLA_NET_0_120037, 
        HIEFFPLA_NET_0_120038, HIEFFPLA_NET_0_120039, 
        HIEFFPLA_NET_0_120040, HIEFFPLA_NET_0_120041, 
        HIEFFPLA_NET_0_120042, HIEFFPLA_NET_0_120043, 
        HIEFFPLA_NET_0_120044, HIEFFPLA_NET_0_120045, 
        HIEFFPLA_NET_0_120046, HIEFFPLA_NET_0_120047, 
        HIEFFPLA_NET_0_120048, HIEFFPLA_NET_0_120049, 
        HIEFFPLA_NET_0_120050, HIEFFPLA_NET_0_120051, 
        HIEFFPLA_NET_0_120052, HIEFFPLA_NET_0_120053, 
        HIEFFPLA_NET_0_120054, HIEFFPLA_NET_0_120055, 
        HIEFFPLA_NET_0_120056, HIEFFPLA_NET_0_120057, 
        HIEFFPLA_NET_0_120058, HIEFFPLA_NET_0_120059, 
        HIEFFPLA_NET_0_120060, HIEFFPLA_NET_0_120061, 
        HIEFFPLA_NET_0_120062, HIEFFPLA_NET_0_120063, 
        HIEFFPLA_NET_0_120064, HIEFFPLA_NET_0_120065, 
        HIEFFPLA_NET_0_120066, HIEFFPLA_NET_0_120067, 
        HIEFFPLA_NET_0_120068, HIEFFPLA_NET_0_120069, 
        HIEFFPLA_NET_0_120070, HIEFFPLA_NET_0_120071, 
        HIEFFPLA_NET_0_120072, HIEFFPLA_NET_0_120073, 
        HIEFFPLA_NET_0_120074, HIEFFPLA_NET_0_120075, 
        HIEFFPLA_NET_0_120076, HIEFFPLA_NET_0_120077, 
        HIEFFPLA_NET_0_120078, HIEFFPLA_NET_0_120079, 
        HIEFFPLA_NET_0_120080, HIEFFPLA_NET_0_120081, 
        HIEFFPLA_NET_0_120082, HIEFFPLA_NET_0_120083, 
        HIEFFPLA_NET_0_120084, HIEFFPLA_NET_0_120085, 
        HIEFFPLA_NET_0_120086, HIEFFPLA_NET_0_120087, 
        HIEFFPLA_NET_0_120088, HIEFFPLA_NET_0_120089, 
        HIEFFPLA_NET_0_120090, HIEFFPLA_NET_0_120091, 
        HIEFFPLA_NET_0_120092, HIEFFPLA_NET_0_120093, 
        HIEFFPLA_NET_0_120094, HIEFFPLA_NET_0_120095, 
        HIEFFPLA_NET_0_120096, HIEFFPLA_NET_0_120097, 
        HIEFFPLA_NET_0_120098, HIEFFPLA_NET_0_120099, 
        HIEFFPLA_NET_0_120100, HIEFFPLA_NET_0_120101, 
        HIEFFPLA_NET_0_120102, HIEFFPLA_NET_0_120103, 
        HIEFFPLA_NET_0_120104, HIEFFPLA_NET_0_120105, 
        HIEFFPLA_NET_0_120106, HIEFFPLA_NET_0_120107, 
        HIEFFPLA_NET_0_120108, HIEFFPLA_NET_0_120109, 
        HIEFFPLA_NET_0_120110, HIEFFPLA_NET_0_120111, 
        HIEFFPLA_NET_0_120112, HIEFFPLA_NET_0_120113, 
        HIEFFPLA_NET_0_120114, HIEFFPLA_NET_0_120115, 
        HIEFFPLA_NET_0_120116, HIEFFPLA_NET_0_120117, 
        HIEFFPLA_NET_0_120118, HIEFFPLA_NET_0_120119, 
        HIEFFPLA_NET_0_120120, HIEFFPLA_NET_0_120121, 
        HIEFFPLA_NET_0_120122, HIEFFPLA_NET_0_120123, 
        HIEFFPLA_NET_0_120124, HIEFFPLA_NET_0_120125, 
        HIEFFPLA_NET_0_120126, HIEFFPLA_NET_0_120127, 
        HIEFFPLA_NET_0_120128, HIEFFPLA_NET_0_120129, 
        HIEFFPLA_NET_0_120130, HIEFFPLA_NET_0_120131, 
        HIEFFPLA_NET_0_120132, HIEFFPLA_NET_0_120133, 
        HIEFFPLA_NET_0_120134, HIEFFPLA_NET_0_120135, 
        HIEFFPLA_NET_0_120136, HIEFFPLA_NET_0_120137, 
        HIEFFPLA_NET_0_120138, HIEFFPLA_NET_0_120139, 
        HIEFFPLA_NET_0_120140, HIEFFPLA_NET_0_120141, 
        HIEFFPLA_NET_0_120142, HIEFFPLA_NET_0_120143, 
        HIEFFPLA_NET_0_120144, HIEFFPLA_NET_0_120145, 
        HIEFFPLA_NET_0_120146, HIEFFPLA_NET_0_120147, 
        HIEFFPLA_NET_0_120148, HIEFFPLA_NET_0_120149, 
        HIEFFPLA_NET_0_120150, HIEFFPLA_NET_0_120151, 
        HIEFFPLA_NET_0_120152, HIEFFPLA_NET_0_120153, 
        HIEFFPLA_NET_0_120154, HIEFFPLA_NET_0_120155, 
        HIEFFPLA_NET_0_120156, HIEFFPLA_NET_0_120157, 
        HIEFFPLA_NET_0_120158, HIEFFPLA_NET_0_120159, 
        HIEFFPLA_NET_0_120160, HIEFFPLA_NET_0_120161, 
        HIEFFPLA_NET_0_120162, HIEFFPLA_NET_0_120163, 
        HIEFFPLA_NET_0_120164, HIEFFPLA_NET_0_120165, 
        HIEFFPLA_NET_0_120166, HIEFFPLA_NET_0_120167, 
        HIEFFPLA_NET_0_120168, HIEFFPLA_NET_0_120169, 
        HIEFFPLA_NET_0_120170, HIEFFPLA_NET_0_120171, 
        HIEFFPLA_NET_0_120172, HIEFFPLA_NET_0_120173, 
        HIEFFPLA_NET_0_120174, HIEFFPLA_NET_0_120175, 
        HIEFFPLA_NET_0_120176, HIEFFPLA_NET_0_120177, 
        HIEFFPLA_NET_0_120178, HIEFFPLA_NET_0_120179, 
        HIEFFPLA_NET_0_120180, HIEFFPLA_NET_0_120181, 
        HIEFFPLA_NET_0_120182, HIEFFPLA_NET_0_120183, 
        HIEFFPLA_NET_0_120184, HIEFFPLA_NET_0_120185, 
        HIEFFPLA_NET_0_120186, HIEFFPLA_NET_0_120187, 
        HIEFFPLA_NET_0_120188, HIEFFPLA_NET_0_120189, 
        HIEFFPLA_NET_0_120190, HIEFFPLA_NET_0_120191, 
        HIEFFPLA_NET_0_120192, HIEFFPLA_NET_0_120193, 
        HIEFFPLA_NET_0_120194, HIEFFPLA_NET_0_120195, 
        HIEFFPLA_NET_0_120196, HIEFFPLA_NET_0_120197, 
        HIEFFPLA_NET_0_120198, HIEFFPLA_NET_0_120199, 
        HIEFFPLA_NET_0_120200, HIEFFPLA_NET_0_120201, 
        HIEFFPLA_NET_0_120202, HIEFFPLA_NET_0_120203, 
        HIEFFPLA_NET_0_120204, HIEFFPLA_NET_0_120205, 
        HIEFFPLA_NET_0_120206, HIEFFPLA_NET_0_120207, 
        HIEFFPLA_NET_0_120208, HIEFFPLA_NET_0_120209, 
        HIEFFPLA_NET_0_120210, HIEFFPLA_NET_0_120211, 
        HIEFFPLA_NET_0_120212, HIEFFPLA_NET_0_120213, 
        HIEFFPLA_NET_0_120214, HIEFFPLA_NET_0_120215, 
        HIEFFPLA_NET_0_120216, HIEFFPLA_NET_0_120217, 
        HIEFFPLA_NET_0_120218, HIEFFPLA_NET_0_120219, 
        HIEFFPLA_NET_0_120220, HIEFFPLA_NET_0_120221, 
        HIEFFPLA_NET_0_120222, HIEFFPLA_NET_0_120223, 
        HIEFFPLA_NET_0_120224, HIEFFPLA_NET_0_120225, 
        HIEFFPLA_NET_0_120226, HIEFFPLA_NET_0_120227, 
        HIEFFPLA_NET_0_120228, HIEFFPLA_NET_0_120229, 
        HIEFFPLA_NET_0_120230, HIEFFPLA_NET_0_120231, 
        HIEFFPLA_NET_0_120232, HIEFFPLA_NET_0_120233, 
        HIEFFPLA_NET_0_120234, HIEFFPLA_NET_0_120235, 
        HIEFFPLA_NET_0_120236, HIEFFPLA_NET_0_120237, 
        HIEFFPLA_NET_0_120238, HIEFFPLA_NET_0_120239, 
        HIEFFPLA_NET_0_120240, HIEFFPLA_NET_0_120241, 
        HIEFFPLA_NET_0_120242, HIEFFPLA_NET_0_120243, 
        HIEFFPLA_NET_0_120244, HIEFFPLA_NET_0_120245, 
        HIEFFPLA_NET_0_120246, HIEFFPLA_NET_0_120247, 
        HIEFFPLA_NET_0_120248, HIEFFPLA_NET_0_120249, 
        HIEFFPLA_NET_0_120250, HIEFFPLA_NET_0_120251, 
        HIEFFPLA_NET_0_120252, HIEFFPLA_NET_0_120253, 
        HIEFFPLA_NET_0_120254, HIEFFPLA_NET_0_120255, 
        HIEFFPLA_NET_0_120256, HIEFFPLA_NET_0_120257, 
        HIEFFPLA_NET_0_120258, HIEFFPLA_NET_0_120259, 
        HIEFFPLA_NET_0_120260, HIEFFPLA_NET_0_120261, 
        HIEFFPLA_NET_0_120262, HIEFFPLA_NET_0_120263, 
        HIEFFPLA_NET_0_120264, HIEFFPLA_NET_0_120265, 
        HIEFFPLA_NET_0_120266, HIEFFPLA_NET_0_120267, 
        HIEFFPLA_NET_0_120268, HIEFFPLA_NET_0_120269, 
        HIEFFPLA_NET_0_120270, HIEFFPLA_NET_0_120271, 
        HIEFFPLA_NET_0_120272, HIEFFPLA_NET_0_120273, 
        HIEFFPLA_NET_0_120274, HIEFFPLA_NET_0_120275, 
        HIEFFPLA_NET_0_120276, HIEFFPLA_NET_0_120277, 
        HIEFFPLA_NET_0_120278, HIEFFPLA_NET_0_120279, 
        HIEFFPLA_NET_0_120280, HIEFFPLA_NET_0_120281, 
        HIEFFPLA_NET_0_120282, HIEFFPLA_NET_0_120283, 
        HIEFFPLA_NET_0_120284, HIEFFPLA_NET_0_120285, 
        HIEFFPLA_NET_0_120286, HIEFFPLA_NET_0_120287, 
        HIEFFPLA_NET_0_120288, HIEFFPLA_NET_0_120289, 
        HIEFFPLA_NET_0_120290, HIEFFPLA_NET_0_120291, 
        HIEFFPLA_NET_0_120292, HIEFFPLA_NET_0_120293, 
        HIEFFPLA_NET_0_120294, HIEFFPLA_NET_0_120295, 
        HIEFFPLA_NET_0_120296, HIEFFPLA_NET_0_120297, 
        HIEFFPLA_NET_0_120298, HIEFFPLA_NET_0_120299, 
        HIEFFPLA_NET_0_120300, HIEFFPLA_NET_0_120301, 
        HIEFFPLA_NET_0_120302, HIEFFPLA_NET_0_120303, 
        HIEFFPLA_NET_0_120304, HIEFFPLA_NET_0_120305, 
        HIEFFPLA_NET_0_120306, HIEFFPLA_NET_0_120307, 
        HIEFFPLA_NET_0_120308, HIEFFPLA_NET_0_120309, 
        HIEFFPLA_NET_0_120310, HIEFFPLA_NET_0_120311, 
        HIEFFPLA_NET_0_120312, HIEFFPLA_NET_0_120313, 
        HIEFFPLA_NET_0_120314, HIEFFPLA_NET_0_120315, 
        HIEFFPLA_NET_0_120316, HIEFFPLA_NET_0_120317, 
        HIEFFPLA_NET_0_120318, HIEFFPLA_NET_0_120319, 
        HIEFFPLA_NET_0_120320, HIEFFPLA_NET_0_120321, 
        HIEFFPLA_NET_0_120322, HIEFFPLA_NET_0_120323, 
        HIEFFPLA_NET_0_120324, HIEFFPLA_NET_0_120325, 
        HIEFFPLA_NET_0_120326, HIEFFPLA_NET_0_120327, 
        HIEFFPLA_NET_0_120328, HIEFFPLA_NET_0_120329, 
        HIEFFPLA_NET_0_120330, HIEFFPLA_NET_0_120331, 
        HIEFFPLA_NET_0_120332, HIEFFPLA_NET_0_120333, 
        HIEFFPLA_NET_0_120334, HIEFFPLA_NET_0_120335, 
        HIEFFPLA_NET_0_120336, HIEFFPLA_NET_0_120337, 
        HIEFFPLA_NET_0_120338, HIEFFPLA_NET_0_120339, 
        HIEFFPLA_NET_0_120340, HIEFFPLA_NET_0_120341, 
        HIEFFPLA_NET_0_120342, HIEFFPLA_NET_0_120343, 
        HIEFFPLA_NET_0_120344, HIEFFPLA_NET_0_120345, 
        HIEFFPLA_NET_0_120346, HIEFFPLA_NET_0_120347, 
        HIEFFPLA_NET_0_120348, HIEFFPLA_NET_0_120349, 
        HIEFFPLA_NET_0_120350, HIEFFPLA_NET_0_120351, 
        HIEFFPLA_NET_0_120352, HIEFFPLA_NET_0_120353, 
        HIEFFPLA_NET_0_120354, HIEFFPLA_NET_0_120355, 
        HIEFFPLA_NET_0_120356, HIEFFPLA_NET_0_120357, 
        HIEFFPLA_NET_0_120358, HIEFFPLA_NET_0_120359, 
        HIEFFPLA_NET_0_120360, HIEFFPLA_NET_0_120361, 
        HIEFFPLA_NET_0_120362, HIEFFPLA_NET_0_120363, 
        HIEFFPLA_NET_0_120364, HIEFFPLA_NET_0_120365, 
        HIEFFPLA_NET_0_120366, HIEFFPLA_NET_0_120367, 
        HIEFFPLA_NET_0_120368, HIEFFPLA_NET_0_161278, 
        HIEFFPLA_NET_0_161279, HIEFFPLA_NET_0_161280, 
        HIEFFPLA_NET_0_161281, HIEFFPLA_NET_0_161282, 
        HIEFFPLA_NET_0_161283, HIEFFPLA_NET_0_161284, 
        HIEFFPLA_NET_0_161285, HIEFFPLA_NET_0_161286, 
        HIEFFPLA_NET_0_161287, HIEFFPLA_NET_0_161288, 
        HIEFFPLA_NET_0_161289, HIEFFPLA_NET_0_161290, 
        HIEFFPLA_NET_0_161291, HIEFFPLA_NET_0_161292, 
        HIEFFPLA_NET_0_161293, HIEFFPLA_NET_0_161294, 
        HIEFFPLA_NET_0_161295, HIEFFPLA_NET_0_161296, 
        HIEFFPLA_NET_0_161297, MASTER_SALT_POR_B_i_0_i, 
        MASTER_SALT_POR_B_i_0_i_0, MASTER_SALT_POR_B_i_0_i_1, 
        MASTER_SALT_POR_B_i_0_i_10, MASTER_SALT_POR_B_i_0_i_11, 
        MASTER_SALT_POR_B_i_0_i_12, MASTER_SALT_POR_B_i_0_i_13, 
        MASTER_SALT_POR_B_i_0_i_14, MASTER_SALT_POR_B_i_0_i_15, 
        MASTER_SALT_POR_B_i_0_i_16, MASTER_SALT_POR_B_i_0_i_17, 
        MASTER_SALT_POR_B_i_0_i_2, MASTER_SALT_POR_B_i_0_i_3, 
        MASTER_SALT_POR_B_i_0_i_4, MASTER_SALT_POR_B_i_0_i_5, 
        MASTER_SALT_POR_B_i_0_i_6, MASTER_SALT_POR_B_i_0_i_7, 
        MASTER_SALT_POR_B_i_0_i_8, MASTER_SALT_POR_B_i_0_i_9, 
        \OP_MODE[0]\, \OP_MODE[4]\, \OP_MODE_c_0[1]\, 
        \OP_MODE_c_1[1]\, \OP_MODE_c_2[1]\, \OP_MODE_c_3[1]\, 
        \OP_MODE_c_4[1]\, \OP_MODE_c_5[1]\, \OP_MODE_c_6[1]\, 
        P_MASTER_POR_B_c_0_0, P_MASTER_POR_B_c_1, 
        P_MASTER_POR_B_c_10, P_MASTER_POR_B_c_11, 
        P_MASTER_POR_B_c_12, P_MASTER_POR_B_c_13, 
        P_MASTER_POR_B_c_14, P_MASTER_POR_B_c_15, 
        P_MASTER_POR_B_c_16, P_MASTER_POR_B_c_16_0, 
        P_MASTER_POR_B_c_17, P_MASTER_POR_B_c_17_0, 
        P_MASTER_POR_B_c_18, P_MASTER_POR_B_c_19, 
        P_MASTER_POR_B_c_2, P_MASTER_POR_B_c_20, 
        P_MASTER_POR_B_c_21, P_MASTER_POR_B_c_22, 
        P_MASTER_POR_B_c_22_0, P_MASTER_POR_B_c_23, 
        P_MASTER_POR_B_c_24, P_MASTER_POR_B_c_24_0, 
        P_MASTER_POR_B_c_25, P_MASTER_POR_B_c_26, 
        P_MASTER_POR_B_c_27, P_MASTER_POR_B_c_27_0, 
        P_MASTER_POR_B_c_27_1, P_MASTER_POR_B_c_28, 
        P_MASTER_POR_B_c_29, P_MASTER_POR_B_c_3, 
        P_MASTER_POR_B_c_30, P_MASTER_POR_B_c_31, 
        P_MASTER_POR_B_c_31_0, P_MASTER_POR_B_c_32, 
        P_MASTER_POR_B_c_32_0, P_MASTER_POR_B_c_33, 
        P_MASTER_POR_B_c_34, P_MASTER_POR_B_c_34_0, 
        P_MASTER_POR_B_c_4, P_MASTER_POR_B_c_5, 
        P_MASTER_POR_B_c_6, P_MASTER_POR_B_c_7, 
        P_MASTER_POR_B_c_8, P_MASTER_POR_B_c_9, 
        P_USB_MASTER_EN_c_1, P_USB_MASTER_EN_c_10, 
        P_USB_MASTER_EN_c_11, P_USB_MASTER_EN_c_12, 
        P_USB_MASTER_EN_c_13, P_USB_MASTER_EN_c_14, 
        P_USB_MASTER_EN_c_15, P_USB_MASTER_EN_c_16, 
        P_USB_MASTER_EN_c_17, P_USB_MASTER_EN_c_18, 
        P_USB_MASTER_EN_c_19, P_USB_MASTER_EN_c_1_0, 
        P_USB_MASTER_EN_c_2, P_USB_MASTER_EN_c_20, 
        P_USB_MASTER_EN_c_21, P_USB_MASTER_EN_c_2_0, 
        P_USB_MASTER_EN_c_3, P_USB_MASTER_EN_c_4, 
        P_USB_MASTER_EN_c_5, P_USB_MASTER_EN_c_6, 
        P_USB_MASTER_EN_c_7, P_USB_MASTER_EN_c_8, 
        P_USB_MASTER_EN_c_9, \TFC_IN_F\, \TFC_IN_R\, 
        \TFC_STOP_ADDR[0]\, \TFC_STOP_ADDR[1]\, 
        \TFC_STOP_ADDR[2]\, \TFC_STOP_ADDR[3]\, 
        \TFC_STOP_ADDR[4]\, \TFC_STOP_ADDR[5]\, 
        \TFC_STOP_ADDR[6]\, \TFC_STOP_ADDR[7]\, 
        \TFC_STRT_ADDR[0]\, \TFC_STRT_ADDR[1]\, 
        \TFC_STRT_ADDR[2]\, \TFC_STRT_ADDR[3]\, 
        \TFC_STRT_ADDR[4]\, \TFC_STRT_ADDR[5]\, 
        \TFC_STRT_ADDR[6]\, \TFC_STRT_ADDR[7]\, 
        \U200A_TFC/GP_PG_SM[0]_net_1\, 
        \U200A_TFC/GP_PG_SM[10]_net_1\, 
        \U200A_TFC/GP_PG_SM[1]_net_1\, 
        \U200A_TFC/GP_PG_SM[2]_net_1\, 
        \U200A_TFC/GP_PG_SM[3]_net_1\, 
        \U200A_TFC/GP_PG_SM[4]_net_1\, 
        \U200A_TFC/GP_PG_SM[5]_net_1\, 
        \U200A_TFC/GP_PG_SM[6]_net_1\, 
        \U200A_TFC/GP_PG_SM[7]_net_1\, 
        \U200A_TFC/GP_PG_SM[8]_net_1\, 
        \U200A_TFC/GP_PG_SM[9]_net_1\, 
        \U200A_TFC/GP_PG_SM_0[10]_net_1\, 
        \U200A_TFC/LOC_STOP_ADDR[0]\, 
        \U200A_TFC/LOC_STOP_ADDR[1]\, 
        \U200A_TFC/LOC_STOP_ADDR[2]\, 
        \U200A_TFC/LOC_STOP_ADDR[3]\, 
        \U200A_TFC/LOC_STOP_ADDR[4]\, 
        \U200A_TFC/LOC_STOP_ADDR[5]\, 
        \U200A_TFC/LOC_STOP_ADDR[6]\, 
        \U200A_TFC/LOC_STOP_ADDR[7]\, 
        \U200A_TFC/LOC_STRT_ADDR[0]\, 
        \U200A_TFC/LOC_STRT_ADDR[1]\, 
        \U200A_TFC/LOC_STRT_ADDR[2]\, 
        \U200A_TFC/LOC_STRT_ADDR[3]\, 
        \U200A_TFC/LOC_STRT_ADDR[4]\, 
        \U200A_TFC/LOC_STRT_ADDR[5]\, 
        \U200A_TFC/LOC_STRT_ADDR[6]\, 
        \U200A_TFC/LOC_STRT_ADDR[7]\, \U200A_TFC/N_232_li\, 
        \U200A_TFC/RX_SER_WORD_1DEL[0]_net_1\, 
        \U200A_TFC/RX_SER_WORD_1DEL[1]_net_1\, 
        \U200A_TFC/RX_SER_WORD_1DEL[2]_net_1\, 
        \U200A_TFC/RX_SER_WORD_1DEL[3]_net_1\, 
        \U200A_TFC/RX_SER_WORD_1DEL[4]_net_1\, 
        \U200A_TFC/RX_SER_WORD_1DEL[5]_net_1\, 
        \U200A_TFC/RX_SER_WORD_1DEL[6]_net_1\, 
        \U200A_TFC/RX_SER_WORD_1DEL[7]_net_1\, 
        \U200A_TFC/RX_SER_WORD_2DEL[0]_net_1\, 
        \U200A_TFC/RX_SER_WORD_2DEL[1]_net_1\, 
        \U200A_TFC/RX_SER_WORD_2DEL[2]_net_1\, 
        \U200A_TFC/RX_SER_WORD_2DEL[3]_net_1\, 
        \U200A_TFC/RX_SER_WORD_2DEL[4]_net_1\, 
        \U200A_TFC/RX_SER_WORD_2DEL[5]_net_1\, 
        \U200A_TFC/RX_SER_WORD_2DEL[6]_net_1\, 
        \U200A_TFC/RX_SER_WORD_2DEL[7]_net_1\, 
        \U200A_TFC/RX_SER_WORD_3DEL[0]_net_1\, 
        \U200A_TFC/RX_SER_WORD_3DEL[4]_net_1\, 
        \U200A_TFC/RX_SER_WORD_3DEL[5]_net_1\, 
        \U200A_TFC/RX_SER_WORD_3DEL[6]_net_1\, 
        \U200A_TFC/RX_SER_WORD_3DEL_i_0[1]\, 
        \U200A_TFC/RX_SER_WORD_3DEL_i_0[2]\, 
        \U200A_TFC/RX_SER_WORD_3DEL_i_0[3]\, 
        \U200A_TFC/RX_SER_WORD_3DEL_i_0[7]\, 
        \U200B_ELINKS/GP_PG_SM[0]_net_1\, 
        \U200B_ELINKS/GP_PG_SM[10]_net_1\, 
        \U200B_ELINKS/GP_PG_SM[1]_net_1\, 
        \U200B_ELINKS/GP_PG_SM[2]_net_1\, 
        \U200B_ELINKS/GP_PG_SM[3]_net_1\, 
        \U200B_ELINKS/GP_PG_SM[4]_net_1\, 
        \U200B_ELINKS/GP_PG_SM[5]_net_1\, 
        \U200B_ELINKS/GP_PG_SM[6]_net_1\, 
        \U200B_ELINKS/GP_PG_SM[7]_net_1\, 
        \U200B_ELINKS/GP_PG_SM[8]_net_1\, 
        \U200B_ELINKS/GP_PG_SM[9]_net_1\, 
        \U200B_ELINKS/GP_PG_SM_0[10]_net_1\, 
        \U200B_ELINKS/LOC_STOP_ADDR[0]\, 
        \U200B_ELINKS/LOC_STOP_ADDR[1]\, 
        \U200B_ELINKS/LOC_STOP_ADDR[2]\, 
        \U200B_ELINKS/LOC_STOP_ADDR[3]\, 
        \U200B_ELINKS/LOC_STOP_ADDR[4]\, 
        \U200B_ELINKS/LOC_STOP_ADDR[5]\, 
        \U200B_ELINKS/LOC_STOP_ADDR[6]\, 
        \U200B_ELINKS/LOC_STOP_ADDR[7]\, 
        \U200B_ELINKS/LOC_STRT_ADDR[0]\, 
        \U200B_ELINKS/LOC_STRT_ADDR[1]\, 
        \U200B_ELINKS/LOC_STRT_ADDR[2]\, 
        \U200B_ELINKS/LOC_STRT_ADDR[3]\, 
        \U200B_ELINKS/LOC_STRT_ADDR[4]\, 
        \U200B_ELINKS/LOC_STRT_ADDR[5]\, 
        \U200B_ELINKS/LOC_STRT_ADDR[6]\, 
        \U200B_ELINKS/LOC_STRT_ADDR[7]\, \U200B_ELINKS/N_232_li\, 
        \U200B_ELINKS/RX_SER_WORD_1DEL[0]_net_1\, 
        \U200B_ELINKS/RX_SER_WORD_1DEL[1]_net_1\, 
        \U200B_ELINKS/RX_SER_WORD_1DEL[2]_net_1\, 
        \U200B_ELINKS/RX_SER_WORD_1DEL[3]_net_1\, 
        \U200B_ELINKS/RX_SER_WORD_1DEL[4]_net_1\, 
        \U200B_ELINKS/RX_SER_WORD_1DEL[5]_net_1\, 
        \U200B_ELINKS/RX_SER_WORD_1DEL[6]_net_1\, 
        \U200B_ELINKS/RX_SER_WORD_1DEL[7]_net_1\, 
        \U200B_ELINKS/RX_SER_WORD_2DEL[0]_net_1\, 
        \U200B_ELINKS/RX_SER_WORD_2DEL[1]_net_1\, 
        \U200B_ELINKS/RX_SER_WORD_2DEL[2]_net_1\, 
        \U200B_ELINKS/RX_SER_WORD_2DEL[3]_net_1\, 
        \U200B_ELINKS/RX_SER_WORD_2DEL[4]_net_1\, 
        \U200B_ELINKS/RX_SER_WORD_2DEL[5]_net_1\, 
        \U200B_ELINKS/RX_SER_WORD_2DEL[6]_net_1\, 
        \U200B_ELINKS/RX_SER_WORD_2DEL[7]_net_1\, 
        \U200B_ELINKS/RX_SER_WORD_3DEL[0]_net_1\, 
        \U200B_ELINKS/RX_SER_WORD_3DEL[4]_net_1\, 
        \U200B_ELINKS/RX_SER_WORD_3DEL[5]_net_1\, 
        \U200B_ELINKS/RX_SER_WORD_3DEL[6]_net_1\, 
        \U200B_ELINKS/RX_SER_WORD_3DEL_i_0[1]\, 
        \U200B_ELINKS/RX_SER_WORD_3DEL_i_0[2]\, 
        \U200B_ELINKS/RX_SER_WORD_3DEL_i_0[3]\, 
        \U200B_ELINKS/RX_SER_WORD_3DEL_i_0[7]\, 
        \U50_PATTERNS/CHKSUM[0]\, \U50_PATTERNS/CHKSUM[1]\, 
        \U50_PATTERNS/CHKSUM[2]\, \U50_PATTERNS/CHKSUM[3]\, 
        \U50_PATTERNS/CHKSUM[4]\, \U50_PATTERNS/CHKSUM[5]\, 
        \U50_PATTERNS/CHKSUM[6]\, \U50_PATTERNS/CHKSUM[7]\, 
        \U50_PATTERNS/ELINKS_STOP_ADDR[0]\, 
        \U50_PATTERNS/ELINKS_STOP_ADDR[1]\, 
        \U50_PATTERNS/ELINKS_STOP_ADDR[2]\, 
        \U50_PATTERNS/ELINKS_STOP_ADDR[3]\, 
        \U50_PATTERNS/ELINKS_STOP_ADDR[4]\, 
        \U50_PATTERNS/ELINKS_STOP_ADDR[5]\, 
        \U50_PATTERNS/ELINKS_STOP_ADDR[6]\, 
        \U50_PATTERNS/ELINKS_STOP_ADDR[7]\, 
        \U50_PATTERNS/ELINKS_STOP_ADDR_T[0]\, 
        \U50_PATTERNS/ELINKS_STOP_ADDR_T[1]\, 
        \U50_PATTERNS/ELINKS_STOP_ADDR_T[2]\, 
        \U50_PATTERNS/ELINKS_STOP_ADDR_T[3]\, 
        \U50_PATTERNS/ELINKS_STOP_ADDR_T[4]\, 
        \U50_PATTERNS/ELINKS_STOP_ADDR_T[5]\, 
        \U50_PATTERNS/ELINKS_STOP_ADDR_T[6]\, 
        \U50_PATTERNS/ELINKS_STOP_ADDR_T[7]\, 
        \U50_PATTERNS/ELINKS_STRT_ADDR[0]\, 
        \U50_PATTERNS/ELINKS_STRT_ADDR[1]\, 
        \U50_PATTERNS/ELINKS_STRT_ADDR[2]\, 
        \U50_PATTERNS/ELINKS_STRT_ADDR[3]\, 
        \U50_PATTERNS/ELINKS_STRT_ADDR[4]\, 
        \U50_PATTERNS/ELINKS_STRT_ADDR[5]\, 
        \U50_PATTERNS/ELINKS_STRT_ADDR[6]\, 
        \U50_PATTERNS/ELINKS_STRT_ADDR[7]\, 
        \U50_PATTERNS/ELINKS_STRT_ADDR_T[0]\, 
        \U50_PATTERNS/ELINKS_STRT_ADDR_T[1]\, 
        \U50_PATTERNS/ELINKS_STRT_ADDR_T[2]\, 
        \U50_PATTERNS/ELINKS_STRT_ADDR_T[3]\, 
        \U50_PATTERNS/ELINKS_STRT_ADDR_T[4]\, 
        \U50_PATTERNS/ELINKS_STRT_ADDR_T[5]\, 
        \U50_PATTERNS/ELINKS_STRT_ADDR_T[6]\, 
        \U50_PATTERNS/ELINKS_STRT_ADDR_T[7]\, 
        \U50_PATTERNS/ELK_N_ACTIVE_net_1\, 
        \U50_PATTERNS/OP_MODE[0]\, \U50_PATTERNS/OP_MODE[1]\, 
        \U50_PATTERNS/OP_MODE[2]\, \U50_PATTERNS/OP_MODE[3]\, 
        \U50_PATTERNS/OP_MODE[4]\, \U50_PATTERNS/OP_MODE[5]\, 
        \U50_PATTERNS/OP_MODE[6]\, \U50_PATTERNS/OP_MODE[7]\, 
        \U50_PATTERNS/OP_MODE_T[0]\, \U50_PATTERNS/OP_MODE_T[1]\, 
        \U50_PATTERNS/OP_MODE_T[2]\, \U50_PATTERNS/OP_MODE_T[3]\, 
        \U50_PATTERNS/OP_MODE_T[4]\, \U50_PATTERNS/OP_MODE_T[5]\, 
        \U50_PATTERNS/OP_MODE_T[6]\, \U50_PATTERNS/OP_MODE_T[7]\, 
        \U50_PATTERNS/RD_XFER_TYPE[0]_net_1\, 
        \U50_PATTERNS/RD_XFER_TYPE[1]_net_1\, 
        \U50_PATTERNS/RD_XFER_TYPE[2]_net_1\, 
        \U50_PATTERNS/RD_XFER_TYPE[3]_net_1\, 
        \U50_PATTERNS/RD_XFER_TYPE[4]_net_1\, 
        \U50_PATTERNS/RD_XFER_TYPE[5]_net_1\, 
        \U50_PATTERNS/RD_XFER_TYPE[6]_net_1\, 
        \U50_PATTERNS/RD_XFER_TYPE[7]_net_1\, 
        \U50_PATTERNS/REG_ADDR[0]\, \U50_PATTERNS/REG_ADDR[1]\, 
        \U50_PATTERNS/REG_ADDR[2]\, \U50_PATTERNS/REG_ADDR[3]\, 
        \U50_PATTERNS/REG_ADDR[4]\, \U50_PATTERNS/REG_ADDR[5]\, 
        \U50_PATTERNS/REG_ADDR[6]\, \U50_PATTERNS/REG_ADDR[7]\, 
        \U50_PATTERNS/REG_ADDR[8]\, 
        \U50_PATTERNS/REG_STATE[0]_net_1\, 
        \U50_PATTERNS/REG_STATE[1]_net_1\, 
        \U50_PATTERNS/REG_STATE[2]_net_1\, 
        \U50_PATTERNS/REG_STATE[3]_net_1\, 
        \U50_PATTERNS/REG_STATE[4]_net_1\, 
        \U50_PATTERNS/REG_STATE[5]_net_1\, 
        \U50_PATTERNS/REG_STATE_0[1]_net_1\, 
        \U50_PATTERNS/REG_STATE_0[2]_net_1\, 
        \U50_PATTERNS/REG_STATE_0[4]_net_1\, 
        \U50_PATTERNS/REG_STATE_0[5]_net_1\, 
        \U50_PATTERNS/SI_CNT[0]\, \U50_PATTERNS/SI_CNT[1]\, 
        \U50_PATTERNS/SI_CNT[2]\, \U50_PATTERNS/SI_CNT[3]\, 
        \U50_PATTERNS/SM_BANK_SEL[0]\, 
        \U50_PATTERNS/SM_BANK_SEL[10]\, 
        \U50_PATTERNS/SM_BANK_SEL[11]\, 
        \U50_PATTERNS/SM_BANK_SEL[12]\, 
        \U50_PATTERNS/SM_BANK_SEL[13]\, 
        \U50_PATTERNS/SM_BANK_SEL[14]\, 
        \U50_PATTERNS/SM_BANK_SEL[15]\, 
        \U50_PATTERNS/SM_BANK_SEL[16]\, 
        \U50_PATTERNS/SM_BANK_SEL[17]\, 
        \U50_PATTERNS/SM_BANK_SEL[18]\, 
        \U50_PATTERNS/SM_BANK_SEL[19]\, 
        \U50_PATTERNS/SM_BANK_SEL[1]\, 
        \U50_PATTERNS/SM_BANK_SEL[20]\, 
        \U50_PATTERNS/SM_BANK_SEL[21]\, 
        \U50_PATTERNS/SM_BANK_SEL[2]\, 
        \U50_PATTERNS/SM_BANK_SEL[3]\, 
        \U50_PATTERNS/SM_BANK_SEL[4]\, 
        \U50_PATTERNS/SM_BANK_SEL[5]\, 
        \U50_PATTERNS/SM_BANK_SEL[6]\, 
        \U50_PATTERNS/SM_BANK_SEL[7]\, 
        \U50_PATTERNS/SM_BANK_SEL[8]\, 
        \U50_PATTERNS/SM_BANK_SEL[9]\, 
        \U50_PATTERNS/SM_BANK_SEL_0[20]\, 
        \U50_PATTERNS/SM_BANK_SEL_0[21]\, 
        \U50_PATTERNS/TFC_STOP_ADDR[0]\, 
        \U50_PATTERNS/TFC_STOP_ADDR[1]\, 
        \U50_PATTERNS/TFC_STOP_ADDR[2]\, 
        \U50_PATTERNS/TFC_STOP_ADDR[3]\, 
        \U50_PATTERNS/TFC_STOP_ADDR[4]\, 
        \U50_PATTERNS/TFC_STOP_ADDR[5]\, 
        \U50_PATTERNS/TFC_STOP_ADDR[6]\, 
        \U50_PATTERNS/TFC_STOP_ADDR[7]\, 
        \U50_PATTERNS/TFC_STOP_ADDR_T[0]\, 
        \U50_PATTERNS/TFC_STOP_ADDR_T[1]\, 
        \U50_PATTERNS/TFC_STOP_ADDR_T[2]\, 
        \U50_PATTERNS/TFC_STOP_ADDR_T[3]\, 
        \U50_PATTERNS/TFC_STOP_ADDR_T[4]\, 
        \U50_PATTERNS/TFC_STOP_ADDR_T[5]\, 
        \U50_PATTERNS/TFC_STOP_ADDR_T[6]\, 
        \U50_PATTERNS/TFC_STOP_ADDR_T[7]\, 
        \U50_PATTERNS/TFC_STRT_ADDR[0]\, 
        \U50_PATTERNS/TFC_STRT_ADDR[1]\, 
        \U50_PATTERNS/TFC_STRT_ADDR[2]\, 
        \U50_PATTERNS/TFC_STRT_ADDR[3]\, 
        \U50_PATTERNS/TFC_STRT_ADDR[4]\, 
        \U50_PATTERNS/TFC_STRT_ADDR[5]\, 
        \U50_PATTERNS/TFC_STRT_ADDR[6]\, 
        \U50_PATTERNS/TFC_STRT_ADDR[7]\, 
        \U50_PATTERNS/TFC_STRT_ADDR_T[0]\, 
        \U50_PATTERNS/TFC_STRT_ADDR_T[1]\, 
        \U50_PATTERNS/TFC_STRT_ADDR_T[2]\, 
        \U50_PATTERNS/TFC_STRT_ADDR_T[3]\, 
        \U50_PATTERNS/TFC_STRT_ADDR_T[4]\, 
        \U50_PATTERNS/TFC_STRT_ADDR_T[5]\, 
        \U50_PATTERNS/TFC_STRT_ADDR_T[6]\, 
        \U50_PATTERNS/TFC_STRT_ADDR_T[7]\, 
        \U50_PATTERNS/U4A_REGCROSS/DELCNT[0]_net_1\, 
        \U50_PATTERNS/U4A_REGCROSS/DELCNT[1]_net_1\, 
        \U50_PATTERNS/U4A_REGCROSS/SAMP_ONE[0]_net_1\, 
        \U50_PATTERNS/U4A_REGCROSS/SAMP_ONE[1]_net_1\, 
        \U50_PATTERNS/U4A_REGCROSS/SAMP_ONE[2]_net_1\, 
        \U50_PATTERNS/U4A_REGCROSS/SAMP_ONE[3]_net_1\, 
        \U50_PATTERNS/U4A_REGCROSS/SAMP_ONE[4]_net_1\, 
        \U50_PATTERNS/U4A_REGCROSS/SAMP_ONE[5]_net_1\, 
        \U50_PATTERNS/U4A_REGCROSS/SAMP_ONE[6]_net_1\, 
        \U50_PATTERNS/U4A_REGCROSS/SAMP_ONE[7]_net_1\, 
        \U50_PATTERNS/U4A_REGCROSS/SAMP_TWO[0]_net_1\, 
        \U50_PATTERNS/U4A_REGCROSS/SAMP_TWO[1]_net_1\, 
        \U50_PATTERNS/U4A_REGCROSS/SAMP_TWO[2]_net_1\, 
        \U50_PATTERNS/U4A_REGCROSS/SAMP_TWO[3]_net_1\, 
        \U50_PATTERNS/U4A_REGCROSS/SAMP_TWO[4]_net_1\, 
        \U50_PATTERNS/U4A_REGCROSS/SAMP_TWO[5]_net_1\, 
        \U50_PATTERNS/U4A_REGCROSS/SAMP_TWO[6]_net_1\, 
        \U50_PATTERNS/U4A_REGCROSS/SAMP_TWO[7]_net_1\, 
        \U50_PATTERNS/U4A_REGCROSS/SYNC_SM[0]_net_1\, 
        \U50_PATTERNS/U4B_REGCROSS/DELCNT[0]_net_1\, 
        \U50_PATTERNS/U4B_REGCROSS/DELCNT[1]_net_1\, 
        \U50_PATTERNS/U4B_REGCROSS/SAMP_ONE[0]_net_1\, 
        \U50_PATTERNS/U4B_REGCROSS/SAMP_ONE[1]_net_1\, 
        \U50_PATTERNS/U4B_REGCROSS/SAMP_ONE[2]_net_1\, 
        \U50_PATTERNS/U4B_REGCROSS/SAMP_ONE[3]_net_1\, 
        \U50_PATTERNS/U4B_REGCROSS/SAMP_ONE[4]_net_1\, 
        \U50_PATTERNS/U4B_REGCROSS/SAMP_ONE[5]_net_1\, 
        \U50_PATTERNS/U4B_REGCROSS/SAMP_ONE[6]_net_1\, 
        \U50_PATTERNS/U4B_REGCROSS/SAMP_ONE[7]_net_1\, 
        \U50_PATTERNS/U4B_REGCROSS/SAMP_TWO[0]_net_1\, 
        \U50_PATTERNS/U4B_REGCROSS/SAMP_TWO[1]_net_1\, 
        \U50_PATTERNS/U4B_REGCROSS/SAMP_TWO[2]_net_1\, 
        \U50_PATTERNS/U4B_REGCROSS/SAMP_TWO[3]_net_1\, 
        \U50_PATTERNS/U4B_REGCROSS/SAMP_TWO[4]_net_1\, 
        \U50_PATTERNS/U4B_REGCROSS/SAMP_TWO[5]_net_1\, 
        \U50_PATTERNS/U4B_REGCROSS/SAMP_TWO[6]_net_1\, 
        \U50_PATTERNS/U4B_REGCROSS/SAMP_TWO[7]_net_1\, 
        \U50_PATTERNS/U4B_REGCROSS/SYNC_SM[0]_net_1\, 
        \U50_PATTERNS/U4C_REGCROSS/DELCNT[0]_net_1\, 
        \U50_PATTERNS/U4C_REGCROSS/DELCNT[1]_net_1\, 
        \U50_PATTERNS/U4C_REGCROSS/SAMP_ONE[0]_net_1\, 
        \U50_PATTERNS/U4C_REGCROSS/SAMP_ONE[1]_net_1\, 
        \U50_PATTERNS/U4C_REGCROSS/SAMP_ONE[2]_net_1\, 
        \U50_PATTERNS/U4C_REGCROSS/SAMP_ONE[3]_net_1\, 
        \U50_PATTERNS/U4C_REGCROSS/SAMP_ONE[4]_net_1\, 
        \U50_PATTERNS/U4C_REGCROSS/SAMP_ONE[5]_net_1\, 
        \U50_PATTERNS/U4C_REGCROSS/SAMP_ONE[6]_net_1\, 
        \U50_PATTERNS/U4C_REGCROSS/SAMP_ONE[7]_net_1\, 
        \U50_PATTERNS/U4C_REGCROSS/SAMP_TWO[0]_net_1\, 
        \U50_PATTERNS/U4C_REGCROSS/SAMP_TWO[1]_net_1\, 
        \U50_PATTERNS/U4C_REGCROSS/SAMP_TWO[2]_net_1\, 
        \U50_PATTERNS/U4C_REGCROSS/SAMP_TWO[3]_net_1\, 
        \U50_PATTERNS/U4C_REGCROSS/SAMP_TWO[4]_net_1\, 
        \U50_PATTERNS/U4C_REGCROSS/SAMP_TWO[5]_net_1\, 
        \U50_PATTERNS/U4C_REGCROSS/SAMP_TWO[6]_net_1\, 
        \U50_PATTERNS/U4C_REGCROSS/SAMP_TWO[7]_net_1\, 
        \U50_PATTERNS/U4C_REGCROSS/SYNC_SM[0]_net_1\, 
        \U50_PATTERNS/U4D_REGCROSS/DELCNT[0]_net_1\, 
        \U50_PATTERNS/U4D_REGCROSS/DELCNT[1]_net_1\, 
        \U50_PATTERNS/U4D_REGCROSS/SAMP_ONE[0]_net_1\, 
        \U50_PATTERNS/U4D_REGCROSS/SAMP_ONE[1]_net_1\, 
        \U50_PATTERNS/U4D_REGCROSS/SAMP_ONE[2]_net_1\, 
        \U50_PATTERNS/U4D_REGCROSS/SAMP_ONE[3]_net_1\, 
        \U50_PATTERNS/U4D_REGCROSS/SAMP_ONE[4]_net_1\, 
        \U50_PATTERNS/U4D_REGCROSS/SAMP_ONE[5]_net_1\, 
        \U50_PATTERNS/U4D_REGCROSS/SAMP_ONE[6]_net_1\, 
        \U50_PATTERNS/U4D_REGCROSS/SAMP_ONE[7]_net_1\, 
        \U50_PATTERNS/U4D_REGCROSS/SAMP_TWO[0]_net_1\, 
        \U50_PATTERNS/U4D_REGCROSS/SAMP_TWO[1]_net_1\, 
        \U50_PATTERNS/U4D_REGCROSS/SAMP_TWO[2]_net_1\, 
        \U50_PATTERNS/U4D_REGCROSS/SAMP_TWO[3]_net_1\, 
        \U50_PATTERNS/U4D_REGCROSS/SAMP_TWO[4]_net_1\, 
        \U50_PATTERNS/U4D_REGCROSS/SAMP_TWO[5]_net_1\, 
        \U50_PATTERNS/U4D_REGCROSS/SAMP_TWO[6]_net_1\, 
        \U50_PATTERNS/U4D_REGCROSS/SAMP_TWO[7]_net_1\, 
        \U50_PATTERNS/U4D_REGCROSS/SYNC_SM[0]_net_1\, 
        \U50_PATTERNS/U4E_REGCROSS/DELCNT[0]_net_1\, 
        \U50_PATTERNS/U4E_REGCROSS/DELCNT[1]_net_1\, 
        \U50_PATTERNS/U4E_REGCROSS/LOCAL_REG_VAL[3]\, 
        \U50_PATTERNS/U4E_REGCROSS/LOCAL_REG_VAL[7]\, 
        \U50_PATTERNS/U4E_REGCROSS/SAMP_ONE[0]_net_1\, 
        \U50_PATTERNS/U4E_REGCROSS/SAMP_ONE[1]_net_1\, 
        \U50_PATTERNS/U4E_REGCROSS/SAMP_ONE[2]_net_1\, 
        \U50_PATTERNS/U4E_REGCROSS/SAMP_ONE[3]_net_1\, 
        \U50_PATTERNS/U4E_REGCROSS/SAMP_ONE[4]_net_1\, 
        \U50_PATTERNS/U4E_REGCROSS/SAMP_ONE[5]_net_1\, 
        \U50_PATTERNS/U4E_REGCROSS/SAMP_ONE[6]_net_1\, 
        \U50_PATTERNS/U4E_REGCROSS/SAMP_ONE[7]_net_1\, 
        \U50_PATTERNS/U4E_REGCROSS/SAMP_TWO[0]_net_1\, 
        \U50_PATTERNS/U4E_REGCROSS/SAMP_TWO[1]_net_1\, 
        \U50_PATTERNS/U4E_REGCROSS/SAMP_TWO[2]_net_1\, 
        \U50_PATTERNS/U4E_REGCROSS/SAMP_TWO[3]_net_1\, 
        \U50_PATTERNS/U4E_REGCROSS/SAMP_TWO[4]_net_1\, 
        \U50_PATTERNS/U4E_REGCROSS/SAMP_TWO[5]_net_1\, 
        \U50_PATTERNS/U4E_REGCROSS/SAMP_TWO[6]_net_1\, 
        \U50_PATTERNS/U4E_REGCROSS/SAMP_TWO[7]_net_1\, 
        \U50_PATTERNS/U4E_REGCROSS/SYNC_SM[0]_net_1\, 
        \U50_PATTERNS/WR_XFER_TYPE[0]_net_1\, 
        \U50_PATTERNS/WR_XFER_TYPE[1]_net_1\, 
        \U50_PATTERNS/WR_XFER_TYPE[2]_net_1\, 
        \U50_PATTERNS/WR_XFER_TYPE[3]_net_1\, 
        \U50_PATTERNS/WR_XFER_TYPE[4]_net_1\, 
        \U50_PATTERNS/WR_XFER_TYPE[5]_net_1\, 
        \U50_PATTERNS/WR_XFER_TYPE[7]_net_1\, 
        \U_ELK0_CMD_TX/CLK40M_GEN_DEL0_net_1\, 
        \U_ELK0_CMD_TX/SER_CMD_WORD_F[0]_net_1\, 
        \U_ELK0_CMD_TX/SER_CMD_WORD_F[1]_net_1\, 
        \U_ELK0_CMD_TX/SER_CMD_WORD_F[3]_net_1\, 
        \U_ELK0_CMD_TX/SER_CMD_WORD_R[0]_net_1\, 
        \U_ELK0_CMD_TX/SER_CMD_WORD_R[1]_net_1\, 
        \U_ELK0_CMD_TX/SER_CMD_WORD_R[2]_net_1\, 
        \U_ELK0_CMD_TX/SER_CMD_WORD_R[3]_net_1\, 
        \U_ELK0_CMD_TX/SER_OUT_FI_i\, 
        \U_ELK0_CMD_TX/SER_OUT_RI_i\, 
        \U_ELK0_CMD_TX/START_RISE_net_1\, 
        \U_ELK10_CH/ELK_TX_DAT[0]\, \U_ELK10_CH/ELK_TX_DAT[1]\, 
        \U_ELK10_CH/ELK_TX_DAT[2]\, \U_ELK10_CH/ELK_TX_DAT[3]\, 
        \U_ELK10_CH/ELK_TX_DAT[4]\, \U_ELK10_CH/ELK_TX_DAT[5]\, 
        \U_ELK10_CH/ELK_TX_DAT[6]\, \U_ELK10_CH/ELK_TX_DAT[7]\, 
        \U_ELK10_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0_net_1\, 
        \U_ELK10_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]_net_1\, 
        \U_ELK10_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]_net_1\, 
        \U_ELK10_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]_net_1\, 
        \U_ELK10_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]_net_1\, 
        \U_ELK10_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]_net_1\, 
        \U_ELK10_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]_net_1\, 
        \U_ELK10_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]_net_1\, 
        \U_ELK10_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]_net_1\, 
        \U_ELK10_CH/U_ELK1_CMD_TX/SER_OUT_FI_net_1\, 
        \U_ELK10_CH/U_ELK1_CMD_TX/SER_OUT_RI_net_1\, 
        \U_ELK10_CH/U_ELK1_CMD_TX/START_RISE_net_1\, 
        \U_ELK11_CH/ELK_TX_DAT[0]\, \U_ELK11_CH/ELK_TX_DAT[1]\, 
        \U_ELK11_CH/ELK_TX_DAT[2]\, \U_ELK11_CH/ELK_TX_DAT[3]\, 
        \U_ELK11_CH/ELK_TX_DAT[4]\, \U_ELK11_CH/ELK_TX_DAT[5]\, 
        \U_ELK11_CH/ELK_TX_DAT[6]\, \U_ELK11_CH/ELK_TX_DAT[7]\, 
        \U_ELK11_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0_net_1\, 
        \U_ELK11_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]_net_1\, 
        \U_ELK11_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]_net_1\, 
        \U_ELK11_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]_net_1\, 
        \U_ELK11_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]_net_1\, 
        \U_ELK11_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]_net_1\, 
        \U_ELK11_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]_net_1\, 
        \U_ELK11_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]_net_1\, 
        \U_ELK11_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]_net_1\, 
        \U_ELK11_CH/U_ELK1_CMD_TX/SER_OUT_FI_net_1\, 
        \U_ELK11_CH/U_ELK1_CMD_TX/SER_OUT_RI_net_1\, 
        \U_ELK11_CH/U_ELK1_CMD_TX/START_RISE_net_1\, 
        \U_ELK12_CH/ELK_TX_DAT[0]\, \U_ELK12_CH/ELK_TX_DAT[1]\, 
        \U_ELK12_CH/ELK_TX_DAT[2]\, \U_ELK12_CH/ELK_TX_DAT[3]\, 
        \U_ELK12_CH/ELK_TX_DAT[4]\, \U_ELK12_CH/ELK_TX_DAT[5]\, 
        \U_ELK12_CH/ELK_TX_DAT[6]\, \U_ELK12_CH/ELK_TX_DAT[7]\, 
        \U_ELK12_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0_net_1\, 
        \U_ELK12_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]_net_1\, 
        \U_ELK12_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]_net_1\, 
        \U_ELK12_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]_net_1\, 
        \U_ELK12_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]_net_1\, 
        \U_ELK12_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]_net_1\, 
        \U_ELK12_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]_net_1\, 
        \U_ELK12_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]_net_1\, 
        \U_ELK12_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]_net_1\, 
        \U_ELK12_CH/U_ELK1_CMD_TX/SER_OUT_FI_net_1\, 
        \U_ELK12_CH/U_ELK1_CMD_TX/SER_OUT_RI_net_1\, 
        \U_ELK12_CH/U_ELK1_CMD_TX/START_RISE_net_1\, 
        \U_ELK13_CH/ELK_TX_DAT[0]\, \U_ELK13_CH/ELK_TX_DAT[1]\, 
        \U_ELK13_CH/ELK_TX_DAT[2]\, \U_ELK13_CH/ELK_TX_DAT[3]\, 
        \U_ELK13_CH/ELK_TX_DAT[4]\, \U_ELK13_CH/ELK_TX_DAT[5]\, 
        \U_ELK13_CH/ELK_TX_DAT[6]\, \U_ELK13_CH/ELK_TX_DAT[7]\, 
        \U_ELK13_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0_net_1\, 
        \U_ELK13_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]_net_1\, 
        \U_ELK13_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]_net_1\, 
        \U_ELK13_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]_net_1\, 
        \U_ELK13_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]_net_1\, 
        \U_ELK13_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]_net_1\, 
        \U_ELK13_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]_net_1\, 
        \U_ELK13_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]_net_1\, 
        \U_ELK13_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]_net_1\, 
        \U_ELK13_CH/U_ELK1_CMD_TX/SER_OUT_FI_net_1\, 
        \U_ELK13_CH/U_ELK1_CMD_TX/SER_OUT_RI_net_1\, 
        \U_ELK13_CH/U_ELK1_CMD_TX/START_RISE_net_1\, 
        \U_ELK14_CH/ELK_TX_DAT[0]\, \U_ELK14_CH/ELK_TX_DAT[1]\, 
        \U_ELK14_CH/ELK_TX_DAT[2]\, \U_ELK14_CH/ELK_TX_DAT[3]\, 
        \U_ELK14_CH/ELK_TX_DAT[4]\, \U_ELK14_CH/ELK_TX_DAT[5]\, 
        \U_ELK14_CH/ELK_TX_DAT[6]\, \U_ELK14_CH/ELK_TX_DAT[7]\, 
        \U_ELK14_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0_net_1\, 
        \U_ELK14_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]_net_1\, 
        \U_ELK14_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]_net_1\, 
        \U_ELK14_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]_net_1\, 
        \U_ELK14_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]_net_1\, 
        \U_ELK14_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]_net_1\, 
        \U_ELK14_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]_net_1\, 
        \U_ELK14_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]_net_1\, 
        \U_ELK14_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]_net_1\, 
        \U_ELK14_CH/U_ELK1_CMD_TX/SER_OUT_FI_net_1\, 
        \U_ELK14_CH/U_ELK1_CMD_TX/SER_OUT_RI_net_1\, 
        \U_ELK14_CH/U_ELK1_CMD_TX/START_RISE_net_1\, 
        \U_ELK15_CH/ELK_TX_DAT[0]\, \U_ELK15_CH/ELK_TX_DAT[1]\, 
        \U_ELK15_CH/ELK_TX_DAT[2]\, \U_ELK15_CH/ELK_TX_DAT[3]\, 
        \U_ELK15_CH/ELK_TX_DAT[4]\, \U_ELK15_CH/ELK_TX_DAT[5]\, 
        \U_ELK15_CH/ELK_TX_DAT[6]\, \U_ELK15_CH/ELK_TX_DAT[7]\, 
        \U_ELK15_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0_net_1\, 
        \U_ELK15_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]_net_1\, 
        \U_ELK15_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]_net_1\, 
        \U_ELK15_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]_net_1\, 
        \U_ELK15_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]_net_1\, 
        \U_ELK15_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]_net_1\, 
        \U_ELK15_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]_net_1\, 
        \U_ELK15_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]_net_1\, 
        \U_ELK15_CH/U_ELK1_CMD_TX/SER_OUT_FI_net_1\, 
        \U_ELK15_CH/U_ELK1_CMD_TX/SER_OUT_RI_net_1\, 
        \U_ELK15_CH/U_ELK1_CMD_TX/START_RISE_net_1\, 
        \U_ELK16_CH/ELK_TX_DAT[0]\, \U_ELK16_CH/ELK_TX_DAT[1]\, 
        \U_ELK16_CH/ELK_TX_DAT[2]\, \U_ELK16_CH/ELK_TX_DAT[3]\, 
        \U_ELK16_CH/ELK_TX_DAT[4]\, \U_ELK16_CH/ELK_TX_DAT[5]\, 
        \U_ELK16_CH/ELK_TX_DAT[6]\, \U_ELK16_CH/ELK_TX_DAT[7]\, 
        \U_ELK16_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0_net_1\, 
        \U_ELK16_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]_net_1\, 
        \U_ELK16_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]_net_1\, 
        \U_ELK16_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]_net_1\, 
        \U_ELK16_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]_net_1\, 
        \U_ELK16_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]_net_1\, 
        \U_ELK16_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]_net_1\, 
        \U_ELK16_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]_net_1\, 
        \U_ELK16_CH/U_ELK1_CMD_TX/SER_OUT_FI_net_1\, 
        \U_ELK16_CH/U_ELK1_CMD_TX/SER_OUT_RI_net_1\, 
        \U_ELK16_CH/U_ELK1_CMD_TX/START_RISE_net_1\, 
        \U_ELK17_CH/ELK_TX_DAT[0]\, \U_ELK17_CH/ELK_TX_DAT[1]\, 
        \U_ELK17_CH/ELK_TX_DAT[2]\, \U_ELK17_CH/ELK_TX_DAT[3]\, 
        \U_ELK17_CH/ELK_TX_DAT[4]\, \U_ELK17_CH/ELK_TX_DAT[5]\, 
        \U_ELK17_CH/ELK_TX_DAT[6]\, \U_ELK17_CH/ELK_TX_DAT[7]\, 
        \U_ELK17_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0_net_1\, 
        \U_ELK17_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]_net_1\, 
        \U_ELK17_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]_net_1\, 
        \U_ELK17_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]_net_1\, 
        \U_ELK17_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]_net_1\, 
        \U_ELK17_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]_net_1\, 
        \U_ELK17_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]_net_1\, 
        \U_ELK17_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]_net_1\, 
        \U_ELK17_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]_net_1\, 
        \U_ELK17_CH/U_ELK1_CMD_TX/SER_OUT_FI_net_1\, 
        \U_ELK17_CH/U_ELK1_CMD_TX/SER_OUT_RI_net_1\, 
        \U_ELK17_CH/U_ELK1_CMD_TX/START_RISE_net_1\, 
        \U_ELK18_CH/ELK_TX_DAT[0]\, \U_ELK18_CH/ELK_TX_DAT[1]\, 
        \U_ELK18_CH/ELK_TX_DAT[2]\, \U_ELK18_CH/ELK_TX_DAT[3]\, 
        \U_ELK18_CH/ELK_TX_DAT[4]\, \U_ELK18_CH/ELK_TX_DAT[5]\, 
        \U_ELK18_CH/ELK_TX_DAT[6]\, \U_ELK18_CH/ELK_TX_DAT[7]\, 
        \U_ELK18_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0_net_1\, 
        \U_ELK18_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]_net_1\, 
        \U_ELK18_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]_net_1\, 
        \U_ELK18_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]_net_1\, 
        \U_ELK18_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]_net_1\, 
        \U_ELK18_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]_net_1\, 
        \U_ELK18_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]_net_1\, 
        \U_ELK18_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]_net_1\, 
        \U_ELK18_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]_net_1\, 
        \U_ELK18_CH/U_ELK1_CMD_TX/SER_OUT_FI_net_1\, 
        \U_ELK18_CH/U_ELK1_CMD_TX/SER_OUT_RI_net_1\, 
        \U_ELK18_CH/U_ELK1_CMD_TX/START_RISE_net_1\, 
        \U_ELK19_CH/ELK_TX_DAT[0]\, \U_ELK19_CH/ELK_TX_DAT[1]\, 
        \U_ELK19_CH/ELK_TX_DAT[2]\, \U_ELK19_CH/ELK_TX_DAT[3]\, 
        \U_ELK19_CH/ELK_TX_DAT[4]\, \U_ELK19_CH/ELK_TX_DAT[5]\, 
        \U_ELK19_CH/ELK_TX_DAT[6]\, \U_ELK19_CH/ELK_TX_DAT[7]\, 
        \U_ELK19_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0_net_1\, 
        \U_ELK19_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]_net_1\, 
        \U_ELK19_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]_net_1\, 
        \U_ELK19_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]_net_1\, 
        \U_ELK19_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]_net_1\, 
        \U_ELK19_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]_net_1\, 
        \U_ELK19_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]_net_1\, 
        \U_ELK19_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]_net_1\, 
        \U_ELK19_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]_net_1\, 
        \U_ELK19_CH/U_ELK1_CMD_TX/SER_OUT_FI_net_1\, 
        \U_ELK19_CH/U_ELK1_CMD_TX/SER_OUT_RI_net_1\, 
        \U_ELK19_CH/U_ELK1_CMD_TX/START_RISE_net_1\, 
        \U_ELK1_CH/ELK_TX_DAT[0]\, \U_ELK1_CH/ELK_TX_DAT[1]\, 
        \U_ELK1_CH/ELK_TX_DAT[2]\, \U_ELK1_CH/ELK_TX_DAT[3]\, 
        \U_ELK1_CH/ELK_TX_DAT[4]\, \U_ELK1_CH/ELK_TX_DAT[5]\, 
        \U_ELK1_CH/ELK_TX_DAT[6]\, \U_ELK1_CH/ELK_TX_DAT[7]\, 
        \U_ELK1_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0_net_1\, 
        \U_ELK1_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]_net_1\, 
        \U_ELK1_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]_net_1\, 
        \U_ELK1_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]_net_1\, 
        \U_ELK1_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]_net_1\, 
        \U_ELK1_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]_net_1\, 
        \U_ELK1_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]_net_1\, 
        \U_ELK1_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]_net_1\, 
        \U_ELK1_CH/U_ELK1_CMD_TX/SER_OUT_FI_i\, 
        \U_ELK1_CH/U_ELK1_CMD_TX/SER_OUT_RI_i\, 
        \U_ELK1_CH/U_ELK1_CMD_TX/START_RISE_net_1\, 
        \U_ELK2_CH/ELK_TX_DAT[0]\, \U_ELK2_CH/ELK_TX_DAT[1]\, 
        \U_ELK2_CH/ELK_TX_DAT[2]\, \U_ELK2_CH/ELK_TX_DAT[3]\, 
        \U_ELK2_CH/ELK_TX_DAT[4]\, \U_ELK2_CH/ELK_TX_DAT[5]\, 
        \U_ELK2_CH/ELK_TX_DAT[6]\, \U_ELK2_CH/ELK_TX_DAT[7]\, 
        \U_ELK2_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0_net_1\, 
        \U_ELK2_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]_net_1\, 
        \U_ELK2_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]_net_1\, 
        \U_ELK2_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]_net_1\, 
        \U_ELK2_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]_net_1\, 
        \U_ELK2_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]_net_1\, 
        \U_ELK2_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]_net_1\, 
        \U_ELK2_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]_net_1\, 
        \U_ELK2_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]_net_1\, 
        \U_ELK2_CH/U_ELK1_CMD_TX/SER_OUT_FI_net_1\, 
        \U_ELK2_CH/U_ELK1_CMD_TX/SER_OUT_RI_net_1\, 
        \U_ELK2_CH/U_ELK1_CMD_TX/START_RISE_net_1\, 
        \U_ELK3_CH/ELK_TX_DAT[0]\, \U_ELK3_CH/ELK_TX_DAT[1]\, 
        \U_ELK3_CH/ELK_TX_DAT[2]\, \U_ELK3_CH/ELK_TX_DAT[3]\, 
        \U_ELK3_CH/ELK_TX_DAT[4]\, \U_ELK3_CH/ELK_TX_DAT[5]\, 
        \U_ELK3_CH/ELK_TX_DAT[6]\, \U_ELK3_CH/ELK_TX_DAT[7]\, 
        \U_ELK3_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0_net_1\, 
        \U_ELK3_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]_net_1\, 
        \U_ELK3_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]_net_1\, 
        \U_ELK3_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]_net_1\, 
        \U_ELK3_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]_net_1\, 
        \U_ELK3_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]_net_1\, 
        \U_ELK3_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]_net_1\, 
        \U_ELK3_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]_net_1\, 
        \U_ELK3_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]_net_1\, 
        \U_ELK3_CH/U_ELK1_CMD_TX/SER_OUT_FI_i\, 
        \U_ELK3_CH/U_ELK1_CMD_TX/SER_OUT_RI_i\, 
        \U_ELK3_CH/U_ELK1_CMD_TX/START_RISE_net_1\, 
        \U_ELK4_CH/ELK_TX_DAT[0]\, \U_ELK4_CH/ELK_TX_DAT[1]\, 
        \U_ELK4_CH/ELK_TX_DAT[2]\, \U_ELK4_CH/ELK_TX_DAT[3]\, 
        \U_ELK4_CH/ELK_TX_DAT[4]\, \U_ELK4_CH/ELK_TX_DAT[5]\, 
        \U_ELK4_CH/ELK_TX_DAT[6]\, \U_ELK4_CH/ELK_TX_DAT[7]\, 
        \U_ELK4_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0_net_1\, 
        \U_ELK4_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]_net_1\, 
        \U_ELK4_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]_net_1\, 
        \U_ELK4_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]_net_1\, 
        \U_ELK4_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]_net_1\, 
        \U_ELK4_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]_net_1\, 
        \U_ELK4_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]_net_1\, 
        \U_ELK4_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]_net_1\, 
        \U_ELK4_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]_net_1\, 
        \U_ELK4_CH/U_ELK1_CMD_TX/SER_OUT_FI_i\, 
        \U_ELK4_CH/U_ELK1_CMD_TX/SER_OUT_RI_i\, 
        \U_ELK4_CH/U_ELK1_CMD_TX/START_RISE_net_1\, 
        \U_ELK5_CH/ELK_TX_DAT[0]\, \U_ELK5_CH/ELK_TX_DAT[1]\, 
        \U_ELK5_CH/ELK_TX_DAT[2]\, \U_ELK5_CH/ELK_TX_DAT[3]\, 
        \U_ELK5_CH/ELK_TX_DAT[4]\, \U_ELK5_CH/ELK_TX_DAT[5]\, 
        \U_ELK5_CH/ELK_TX_DAT[6]\, \U_ELK5_CH/ELK_TX_DAT[7]\, 
        \U_ELK5_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0_net_1\, 
        \U_ELK5_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]_net_1\, 
        \U_ELK5_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]_net_1\, 
        \U_ELK5_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]_net_1\, 
        \U_ELK5_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]_net_1\, 
        \U_ELK5_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]_net_1\, 
        \U_ELK5_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]_net_1\, 
        \U_ELK5_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]_net_1\, 
        \U_ELK5_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]_net_1\, 
        \U_ELK5_CH/U_ELK1_CMD_TX/SER_OUT_FI_net_1\, 
        \U_ELK5_CH/U_ELK1_CMD_TX/SER_OUT_RI_net_1\, 
        \U_ELK5_CH/U_ELK1_CMD_TX/START_RISE_net_1\, 
        \U_ELK6_CH/ELK_TX_DAT[0]\, \U_ELK6_CH/ELK_TX_DAT[1]\, 
        \U_ELK6_CH/ELK_TX_DAT[2]\, \U_ELK6_CH/ELK_TX_DAT[3]\, 
        \U_ELK6_CH/ELK_TX_DAT[4]\, \U_ELK6_CH/ELK_TX_DAT[5]\, 
        \U_ELK6_CH/ELK_TX_DAT[6]\, \U_ELK6_CH/ELK_TX_DAT[7]\, 
        \U_ELK6_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0_net_1\, 
        \U_ELK6_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]_net_1\, 
        \U_ELK6_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]_net_1\, 
        \U_ELK6_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]_net_1\, 
        \U_ELK6_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]_net_1\, 
        \U_ELK6_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]_net_1\, 
        \U_ELK6_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]_net_1\, 
        \U_ELK6_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]_net_1\, 
        \U_ELK6_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]_net_1\, 
        \U_ELK6_CH/U_ELK1_CMD_TX/SER_OUT_FI_net_1\, 
        \U_ELK6_CH/U_ELK1_CMD_TX/SER_OUT_RI_net_1\, 
        \U_ELK6_CH/U_ELK1_CMD_TX/START_RISE_net_1\, 
        \U_ELK7_CH/ELK_TX_DAT[0]\, \U_ELK7_CH/ELK_TX_DAT[1]\, 
        \U_ELK7_CH/ELK_TX_DAT[2]\, \U_ELK7_CH/ELK_TX_DAT[3]\, 
        \U_ELK7_CH/ELK_TX_DAT[4]\, \U_ELK7_CH/ELK_TX_DAT[5]\, 
        \U_ELK7_CH/ELK_TX_DAT[6]\, \U_ELK7_CH/ELK_TX_DAT[7]\, 
        \U_ELK7_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0_net_1\, 
        \U_ELK7_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]_net_1\, 
        \U_ELK7_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]_net_1\, 
        \U_ELK7_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]_net_1\, 
        \U_ELK7_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]_net_1\, 
        \U_ELK7_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]_net_1\, 
        \U_ELK7_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]_net_1\, 
        \U_ELK7_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]_net_1\, 
        \U_ELK7_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]_net_1\, 
        \U_ELK7_CH/U_ELK1_CMD_TX/SER_OUT_FI_net_1\, 
        \U_ELK7_CH/U_ELK1_CMD_TX/SER_OUT_RI_net_1\, 
        \U_ELK7_CH/U_ELK1_CMD_TX/START_RISE_net_1\, 
        \U_ELK8_CH/ELK_TX_DAT[0]\, \U_ELK8_CH/ELK_TX_DAT[1]\, 
        \U_ELK8_CH/ELK_TX_DAT[2]\, \U_ELK8_CH/ELK_TX_DAT[3]\, 
        \U_ELK8_CH/ELK_TX_DAT[4]\, \U_ELK8_CH/ELK_TX_DAT[5]\, 
        \U_ELK8_CH/ELK_TX_DAT[6]\, \U_ELK8_CH/ELK_TX_DAT[7]\, 
        \U_ELK8_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0_net_1\, 
        \U_ELK8_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]_net_1\, 
        \U_ELK8_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]_net_1\, 
        \U_ELK8_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]_net_1\, 
        \U_ELK8_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]_net_1\, 
        \U_ELK8_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]_net_1\, 
        \U_ELK8_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]_net_1\, 
        \U_ELK8_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]_net_1\, 
        \U_ELK8_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]_net_1\, 
        \U_ELK8_CH/U_ELK1_CMD_TX/SER_OUT_FI_net_1\, 
        \U_ELK8_CH/U_ELK1_CMD_TX/SER_OUT_RI_net_1\, 
        \U_ELK8_CH/U_ELK1_CMD_TX/START_RISE_net_1\, 
        \U_ELK9_CH/ELK_TX_DAT[0]\, \U_ELK9_CH/ELK_TX_DAT[1]\, 
        \U_ELK9_CH/ELK_TX_DAT[2]\, \U_ELK9_CH/ELK_TX_DAT[3]\, 
        \U_ELK9_CH/ELK_TX_DAT[4]\, \U_ELK9_CH/ELK_TX_DAT[5]\, 
        \U_ELK9_CH/ELK_TX_DAT[6]\, \U_ELK9_CH/ELK_TX_DAT[7]\, 
        \U_ELK9_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0_net_1\, 
        \U_ELK9_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]_net_1\, 
        \U_ELK9_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]_net_1\, 
        \U_ELK9_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]_net_1\, 
        \U_ELK9_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]_net_1\, 
        \U_ELK9_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]_net_1\, 
        \U_ELK9_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]_net_1\, 
        \U_ELK9_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]_net_1\, 
        \U_ELK9_CH/U_ELK1_CMD_TX/SER_OUT_FI_net_1\, 
        \U_ELK9_CH/U_ELK1_CMD_TX/SER_OUT_RI_net_1\, 
        \U_ELK9_CH/U_ELK1_CMD_TX/START_RISE_net_1\, 
        \U_EXEC_MASTER/CCC_1_LOCK_STAT_0D_net_1\, 
        \U_EXEC_MASTER/CCC_1_LOCK_STAT_1D_net_1\, 
        \U_EXEC_MASTER/DEL_CNT[0]\, \U_EXEC_MASTER/DEL_CNT[1]\, 
        \U_EXEC_MASTER/DEL_CNT[2]\, \U_EXEC_MASTER/DEL_CNT[3]\, 
        \U_EXEC_MASTER/DEL_CNT[4]\, \U_EXEC_MASTER/DEL_CNT[5]\, 
        \U_EXEC_MASTER/DEL_CNT[6]\, \U_EXEC_MASTER/DEL_CNT[7]\, 
        \U_EXEC_MASTER/DEV_RST_0B_net_1\, 
        \U_EXEC_MASTER/DEV_RST_1B_i\, \U_EXEC_MASTER/PRESCALE[0]\, 
        \U_EXEC_MASTER/PRESCALE[1]\, \U_EXEC_MASTER/PRESCALE[2]\, 
        \U_EXEC_MASTER/PRESCALE[3]\, 
        \U_EXEC_MASTER/P_MASTER_POR_B_c_0\, 
        \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i\, 
        \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_0\, 
        \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_1\, 
        \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_2\, 
        \U_EXEC_MASTER/USB_MASTER_EN/CNT_EN_40M_net_1\, 
        \U_EXEC_MASTER/USB_MASTER_EN/CNT_EN_60M0S_net_1\, 
        \U_EXEC_MASTER/USB_MASTER_EN/CNT_EN_60M1S_net_1\, 
        \U_EXEC_MASTER/USB_MASTER_EN/CNT_EN_60M2S_net_1\, 
        \U_EXEC_MASTER/USB_MASTER_EN/TERMCNT_FG40M0S_net_1\, 
        \U_EXEC_MASTER/USB_MASTER_EN/TERMCNT_FG40M1S_net_1\, 
        \U_EXEC_MASTER/USB_MASTER_EN/TERMCNT_FG40M2S_net_1\, 
        \U_EXEC_MASTER/USB_MASTER_EN/TERMCNT_FG60M_net_1\, 
        \U_EXEC_MASTER/USB_MASTER_EN/TEST_SM[0]_net_1\, 
        \U_EXEC_MASTER/USB_MASTER_EN/TEST_SM[1]_net_1\, 
        \U_EXEC_MASTER/USB_MASTER_EN/TEST_SM[3]_net_1\, 
        \U_EXEC_MASTER/USB_MASTER_EN/TEST_SM[4]_net_1\, 
        \U_EXEC_MASTER/USB_MASTER_EN/TEST_SM_i_0[2]\, 
        \U_EXEC_MASTER/USB_MASTER_EN/T_CNT60M[0]_net_1\, 
        \U_EXEC_MASTER/USB_MASTER_EN/T_CNT60M[1]_net_1\, 
        \U_EXEC_MASTER/USB_MASTER_EN/T_CNT60M[2]_net_1\, 
        \U_EXEC_MASTER/USB_MASTER_EN/T_CNT60M[3]_net_1\, 
        \U_EXEC_MASTER/USB_MASTER_EN/T_CNT60M[4]_net_1\, 
        \U_EXEC_MASTER/USB_MASTER_EN/T_CNT60M[5]_net_1\, 
        \U_EXEC_MASTER/USB_MASTER_EN/T_CNT60M[6]_net_1\, 
        \U_EXEC_MASTER/USB_MASTER_EN/T_CNT60M[7]_net_1\, 
        \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_40M_net_1\, 
        \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_1S_net_1\, 
        \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_1S_0_net_1\, 
        \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_S_net_1\, 
        \U_GEN_REF_CLK/GEN_40M_REFCNT[0]_net_1\, 
        \U_GEN_REF_CLK/GEN_40M_REFCNT[1]_net_1\, 
        \U_GEN_REF_CLK/GEN_40M_REFCNT[2]_net_1\, 
        \U_MASTER_DES/CCC2_CONFIG_TRIG\, 
        \U_MASTER_DES/PHASE_ADJ_160_L[0]\, 
        \U_MASTER_DES/PHASE_ADJ_160_L[1]\, 
        \U_MASTER_DES/PHASE_ADJ_160_L[2]\, 
        \U_MASTER_DES/PHASE_ADJ_160_L[3]\, 
        \U_MASTER_DES/PHASE_ADJ_160_L[4]\, 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[0]_net_1\, 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[10]_net_1\, 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[11]_net_1\, 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[1]_net_1\, 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[2]_net_1\, 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[31]_net_1\, 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[34]_net_1\, 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[37]_net_1\, 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[39]_net_1\, 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[40]_net_1\, 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[41]_net_1\, 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[42]_net_1\, 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[44]_net_1\, 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[46]\, 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[47]\, 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[48]\, 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[49]\, 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[50]\, 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[71]_net_1\, 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[72]_net_1\, 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[73]_net_1\, 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[76]_net_1\, 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[77]_net_1\, 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[78]_net_1\, 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[79]_net_1\, 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[7]_net_1\, 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[8]_net_1\, 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[9]_net_1\, 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[0]\, 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[1]\, 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[2]\, 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[3]\, 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[4]\, 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[5]\, 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[6]\, 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[7]\, 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM[0]_net_1\, 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM[1]_net_1\, 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM[2]_net_1\, 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM[3]_net_1\, 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM[4]_net_1\, 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM[5]_net_1\, 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM[6]_net_1\, 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM_0[4]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[0]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[10]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[11]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[12]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[13]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[14]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[1]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[2]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[3]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[4]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[5]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[6]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[7]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[8]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[9]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_SER_IN_F_1DEL_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_SER_IN_R_1DEL_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[0]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[10]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[11]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[12]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[13]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[14]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[1]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[2]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[3]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[4]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[5]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[6]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[7]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[8]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[9]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_WRD_40M_FIXED[0]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_WRD_40M_FIXED[10]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_WRD_40M_FIXED[11]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_WRD_40M_FIXED[12]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_WRD_40M_FIXED[13]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_WRD_40M_FIXED[14]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_WRD_40M_FIXED[1]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_WRD_40M_FIXED[2]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_WRD_40M_FIXED[3]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_WRD_40M_FIXED[4]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_WRD_40M_FIXED[5]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_WRD_40M_FIXED[6]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_WRD_40M_FIXED[7]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_WRD_40M_FIXED[8]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_WRD_40M_FIXED[9]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_BIT_OS_VAL[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_BIT_OS_VAL[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_BIT_OS_VAL[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_BIT_OS_VAL[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_CLKPHASE[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_CLKPHASE[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_CLKPHASE[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_CLKPHASE[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_CLKPHASE[4]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_SEQCNT[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_SEQCNT[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_SEQCNT[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_SEQCNT[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_SEQCNT[4]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_0[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_0[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_0[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_0[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_0[4]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_0[5]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_0[6]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_0[7]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_0[8]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_1[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_1[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_1[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_1[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_1[4]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_1[5]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_1[6]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_1[7]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_1[8]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_2[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_2[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_2[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_2[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_2[4]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_2[5]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_2[6]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_2[7]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_2[8]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_3[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_3[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_3[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_3[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_3[4]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_3[5]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_3[6]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_3[7]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_3[8]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_4[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_4[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_4[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_4[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_4[4]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_4[5]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_4[6]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_4[7]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_4[8]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_5[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_5[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_5[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_5[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_5[4]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_5[5]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_5[6]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_5[7]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_5[8]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_6[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_6[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_6[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_6[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_6[4]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_6[5]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_6[6]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_6[7]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_6[8]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_7[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_7[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_7[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_7[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_7[4]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_7[5]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_7[6]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_7[7]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_7[8]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_SEL[3]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_0[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_0[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_0[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_0[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_10[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_10[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_10[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_10[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_11[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_11[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_11[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_11[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_12[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_12[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_12[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_12[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_13[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_13[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_13[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_13[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_14[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_14[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_14[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_14[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_15[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_15[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_15[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_15[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_16[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_16[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_16[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_16[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_17[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_17[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_17[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_17[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_18[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_18[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_18[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_18[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_19[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_19[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_19[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_19[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_1[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_1[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_1[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_1[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_20[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_20[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_20[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_20[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_21[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_21[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_21[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_21[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_22[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_22[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_22[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_22[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_23[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_23[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_23[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_23[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_24[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_24[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_24[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_24[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_25[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_25[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_25[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_25[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_26[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_26[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_26[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_26[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_27[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_27[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_27[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_27[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_28[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_28[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_28[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_28[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_29[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_29[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_29[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_29[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_2[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_2[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_2[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_2[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_30[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_30[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_30[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_30[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_31[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_31[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_31[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_31[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_3[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_3[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_3[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_3[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_4[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_4[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_4[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_4[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_5[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_5[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_5[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_5[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_6[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_6[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_6[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_6[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_7[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_7[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_7[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_7[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_8[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_8[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_8[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_8[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_9[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_9[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_9[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_9[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[0]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[1]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[2]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[3]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[4]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[0]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[1]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[2]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[3]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[4]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_1[3]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_1[4]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_2[3]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_2[4]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_3[4]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_4[4]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_5[4]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[0]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[1]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[2]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[3]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[4]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[5]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[6]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[7]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[8]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_0[6]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_0[8]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_1[6]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_2[6]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_3[6]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[4]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_1[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_1[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_2[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_2[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_3[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_4[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/MAX_CNT[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/MAX_CNT[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/MAX_CNT[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/MAX_CNT[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/MAX_CNT[4]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/MAX_CNT[5]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/MAX_CNT[6]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/MAX_CNT[7]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/MAX_CNT[8]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/Q[0]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/Q[10]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/Q[11]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/Q[12]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/Q[13]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/Q[14]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/Q[1]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/Q[2]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/Q[3]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/Q[4]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/Q[5]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/Q[6]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/Q[7]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/Q[8]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/Q[9]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/RECD_SER_WORD[0]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/RECD_SER_WORD[1]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/RECD_SER_WORD[2]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/RECD_SER_WORD[3]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/RECD_SER_WORD[4]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/RECD_SER_WORD[5]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/RECD_SER_WORD[6]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/RECD_SER_WORD[7]_net_1\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_10[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_10[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_10[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_10[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_10[4]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_11[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_11[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_11[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_11[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_11[4]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_12[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_12[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_12[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_12[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_12[4]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_13[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_13[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_13[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_13[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_13[4]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_14[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_14[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_14[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_14[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_14[4]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_15[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_15[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_15[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_15[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_15[4]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_16[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_16[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_16[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_16[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_16[4]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_17[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_17[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_17[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_17[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_17[4]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_18[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_18[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_18[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_18[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_18[4]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_19[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_19[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_19[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_19[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_19[4]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_1[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_1[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_1[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_1[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_1[4]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_20[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_20[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_20[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_20[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_20[4]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_21[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_21[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_21[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_21[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_21[4]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_22[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_22[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_22[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_22[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_22[4]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_23[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_23[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_23[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_23[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_23[4]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_24[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_24[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_24[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_24[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_24[4]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_25[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_25[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_25[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_25[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_25[4]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_26[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_26[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_26[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_26[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_26[4]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_27[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_27[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_27[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_27[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_27[4]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_28[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_28[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_28[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_28[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_28[4]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_29[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_29[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_29[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_29[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_29[4]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_2[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_2[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_2[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_2[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_2[4]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_30[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_30[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_30[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_30[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_30[4]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_31[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_31[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_31[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_31[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_31[4]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_3[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_3[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_3[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_3[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_3[4]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_4[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_4[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_4[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_4[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_4[4]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_5[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_5[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_5[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_5[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_5[4]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_6[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_6[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_6[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_6[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_6[4]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_7[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_7[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_7[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_7[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_7[4]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_8[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_8[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_8[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_8[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_8[4]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_9[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_9[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_9[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_9[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_9[4]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/TUNE_CLKPHASE[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/TUNE_CLKPHASE[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/TUNE_CLKPHASE[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/TUNE_CLKPHASE[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/TUNE_CLKPHASE[4]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[0]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[10]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[11]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[12]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[13]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[1]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[2]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[3]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[4]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[5]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[6]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[7]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[8]\, 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[9]\, AFLSDF_VCC, 
        AFLSDF_GND, \AFLSDF_INV_0\, \AFLSDF_INV_1\, 
        \AFLSDF_INV_2\, \AFLSDF_INV_3\, \AFLSDF_INV_4\, 
        \AFLSDF_INV_5\, \AFLSDF_INV_6\, \AFLSDF_INV_7\, 
        \AFLSDF_INV_8\, \AFLSDF_INV_9\, \AFLSDF_INV_10\, 
        \AFLSDF_INV_11\, \AFLSDF_INV_12\, \AFLSDF_INV_13\, 
        \AFLSDF_INV_14\, \AFLSDF_INV_15\, \AFLSDF_INV_16\, 
        \AFLSDF_INV_17\, \AFLSDF_INV_18\, \AFLSDF_INV_19\, 
        \AFLSDF_INV_20\, \AFLSDF_INV_21\, \AFLSDF_INV_22\, 
        \AFLSDF_INV_23\, \AFLSDF_INV_24\, \AFLSDF_INV_25\, 
        \AFLSDF_INV_26\, \AFLSDF_INV_27\, \AFLSDF_INV_28\, 
        \AFLSDF_INV_29\, \AFLSDF_INV_30\, \AFLSDF_INV_31\, 
        \AFLSDF_INV_32\, \AFLSDF_INV_33\, \AFLSDF_INV_34\, 
        \AFLSDF_INV_35\, \AFLSDF_INV_36\, \AFLSDF_INV_37\, 
        \AFLSDF_INV_38\, \AFLSDF_INV_39\, \AFLSDF_INV_40\, 
        \AFLSDF_INV_41\, \AFLSDF_INV_42\, \AFLSDF_INV_43\, 
        \AFLSDF_INV_44\, \AFLSDF_INV_45\, \AFLSDF_INV_46\, 
        \AFLSDF_INV_47\, \AFLSDF_INV_48\, \AFLSDF_INV_49\, 
        \AFLSDF_INV_50\, \AFLSDF_INV_51\, \AFLSDF_INV_52\, 
        \AFLSDF_INV_53\, \AFLSDF_INV_54\, \AFLSDF_INV_55\, 
        \AFLSDF_INV_56\, \AFLSDF_INV_57\, \AFLSDF_INV_58\, 
        \AFLSDF_INV_59\, \AFLSDF_INV_60\, \AFLSDF_INV_61\, 
        \AFLSDF_INV_62\, \AFLSDF_INV_63\, \AFLSDF_INV_64\, 
        \AFLSDF_INV_65\, \AFLSDF_INV_66\, \AFLSDF_INV_67\, 
        \AFLSDF_INV_68\ : std_logic;
    signal GND_power_net1 : std_logic;
    signal VCC_power_net1 : std_logic;

begin 

    AFLSDF_GND <= GND_power_net1;
    \GND\ <= GND_power_net1;
    \VCC\ <= VCC_power_net1;
    AFLSDF_VCC <= VCC_power_net1;

    \U_ELK10_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118650, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_6, Q => 
        \U_ELK10_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]_net_1\);
    
    HIEFFPLA_INST_0_61841 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_27[0]\, B => 
        HIEFFPLA_NET_0_117096, S => HIEFFPLA_NET_0_117196, Y => 
        HIEFFPLA_NET_0_116070);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_3[4]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116721, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_7, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_3[4]\);
    
    \U_ELK19_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]\ : DFN1C0
      port map(D => \U_ELK19_CH/U_SLAVE_1ELK/Q[14]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]_net_1\);
    
    \DCB_SALT_SEL_pad/U0/U1\ : IOIN_IB
      port map(YIN => \DCB_SALT_SEL_pad/U0/NET1\, Y => 
        DCB_SALT_SEL_c);
    
    \U50_PATTERNS/U4C_REGCROSS/SAMP_ONE[6]\ : DFN1C0
      port map(D => \U50_PATTERNS/ELINKS_STRT_ADDR[6]\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_33, Q => 
        \U50_PATTERNS/U4C_REGCROSS/SAMP_ONE[6]_net_1\);
    
    HIEFFPLA_INST_0_58396 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_14[1]\, B => 
        HIEFFPLA_NET_0_116677, S => HIEFFPLA_NET_0_117159, Y => 
        HIEFFPLA_NET_0_116527);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_3[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116337, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_19, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_3[2]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117044, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_17, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[1]\);
    
    HIEFFPLA_INST_0_55296 : AND3
      port map(A => HIEFFPLA_NET_0_115951, B => 
        HIEFFPLA_NET_0_117027, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[4]_net_1\, Y => 
        HIEFFPLA_NET_0_117068);
    
    HIEFFPLA_INST_0_53716 : AO1D
      port map(A => HIEFFPLA_NET_0_116678, B => 
        HIEFFPLA_NET_0_116593, C => HIEFFPLA_NET_0_117396, Y => 
        HIEFFPLA_NET_0_117367);
    
    HIEFFPLA_INST_0_55206 : AND2A
      port map(A => HIEFFPLA_NET_0_117207, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[6]_net_1\, Y => 
        HIEFFPLA_NET_0_117091);
    
    HIEFFPLA_INST_0_54021 : AO1B
      port map(A => HIEFFPLA_NET_0_117147, B => 
        HIEFFPLA_NET_0_117335, C => HIEFFPLA_NET_0_117086, Y => 
        HIEFFPLA_NET_0_117319);
    
    HIEFFPLA_INST_0_43663 : NAND2B
      port map(A => \U50_PATTERNS/SM_BANK_SEL[21]\, B => 
        \U50_PATTERNS/SM_BANK_SEL[5]\, Y => HIEFFPLA_NET_0_119249);
    
    HIEFFPLA_INST_0_61517 : MX2
      port map(A => HIEFFPLA_NET_0_117166, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_23[4]\, S => 
        HIEFFPLA_NET_0_117151, Y => HIEFFPLA_NET_0_116116);
    
    \U_ELK7_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U1\ : IOBI_ID_OD_EB
      port map(DR => \U_ELK7_CH/ELK_OUT_R\, DF => 
        \U_ELK7_CH/ELK_OUT_F\, CLR => \GND\, E => \AFLSDF_INV_46\, 
        ICLK => CCC_160M_ADJ, OCLK => CCC_160M_FXD, YIN => 
        \U_ELK7_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\, DOUT => 
        \U_ELK7_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, EOUT => 
        \U_ELK7_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET2\, YR => 
        \U_ELK7_CH/ELK_IN_DDR_R\, YF => \U_ELK7_CH/ELK_IN_DDR_F\);
    
    \U_ELK2_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL\ : DFN1C0
      port map(D => \U_ELK2_CH/ELK_IN_R_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL_net_1\);
    
    HIEFFPLA_INST_0_43076 : AND3
      port map(A => HIEFFPLA_NET_0_119389, B => 
        \U50_PATTERNS/REG_STATE[0]_net_1\, C => 
        HIEFFPLA_NET_0_119511, Y => HIEFFPLA_NET_0_119386);
    
    \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[13]\ : DFN1C0
      port map(D => 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]_net_1\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[13]_net_1\);
    
    HIEFFPLA_INST_0_43671 : AND2A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/SM_BANK_SEL[16]\, Y => 
        HIEFFPLA_NET_0_119246);
    
    HIEFFPLA_INST_0_37958 : MX2
      port map(A => \U200B_ELINKS/LOC_STOP_ADDR[4]\, B => 
        \ELKS_STOP_ADDR[4]\, S => 
        \U200B_ELINKS/GP_PG_SM_0[10]_net_1\, Y => 
        HIEFFPLA_NET_0_120183);
    
    HIEFFPLA_INST_0_111663 : AOI1
      port map(A => HIEFFPLA_NET_0_115834, B => 
        HIEFFPLA_NET_0_117684, C => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[5]\, Y => 
        HIEFFPLA_NET_0_117666);
    
    HIEFFPLA_INST_0_58902 : AND2A
      port map(A => HIEFFPLA_NET_0_117203, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_3[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116460);
    
    HIEFFPLA_INST_0_47523 : MX2
      port map(A => HIEFFPLA_NET_0_118498, B => 
        HIEFFPLA_NET_0_118495, S => \BIT_OS_SEL_4[0]\, Y => 
        \U_ELK13_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[4]\);
    
    \U_ELK17_CH/U_ELK1_CMD_TX/SER_OUT_RI\ : DFN1C0
      port map(D => 
        \U_ELK17_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_0, Q => 
        \U_ELK17_CH/U_ELK1_CMD_TX/SER_OUT_RI_net_1\);
    
    \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[11]\ : DFN1C0
      port map(D => \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\);
    
    HIEFFPLA_INST_0_48784 : MX2
      port map(A => HIEFFPLA_NET_0_118261, B => 
        HIEFFPLA_NET_0_118275, S => \BIT_OS_SEL_2[0]\, Y => 
        \U_ELK18_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[6]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_1[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117023, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_16_0, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_1[0]\);
    
    \U50_PATTERNS/REG_ADDR[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119529, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_10, Q => \U50_PATTERNS/REG_ADDR[4]\);
    
    \U50_PATTERNS/ELINK_ADDRA_3[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119991, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_1, Q => 
        \U50_PATTERNS/ELINK_ADDRA_3[0]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_24[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116431, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_18, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_24[3]\);
    
    HIEFFPLA_INST_0_46833 : AND2
      port map(A => \U_ELK11_CH/ELK_TX_DAT[0]\, B => 
        \U_ELK11_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118607);
    
    \U_ELK5_CH/U_ELK1_SERDAT_SOURCE/SERDAT[4]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118009, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i, Q => 
        \U_ELK5_CH/ELK_TX_DAT[4]\);
    
    \U_ELK7_CH/U_SLAVE_1ELK/RECD_SER_WORD[1]\ : DFN1C0
      port map(D => \U_ELK7_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[1]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_7[1]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_3[4]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_115935, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_24_0, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_3[4]_net_1\);
    
    \U_ELK13_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U1\ : IOBI_ID_OD_EB
      port map(DR => \U_ELK13_CH/ELK_OUT_R\, DF => 
        \U_ELK13_CH/ELK_OUT_F\, CLR => \GND\, E => 
        \AFLSDF_INV_20\, ICLK => CCC_160M_ADJ, OCLK => 
        CCC_160M_FXD, YIN => 
        \U_ELK13_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\, DOUT => 
        \U_ELK13_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, EOUT => 
        \U_ELK13_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET2\, YR => 
        \U_ELK13_CH/ELK_IN_DDR_R\, YF => 
        \U_ELK13_CH/ELK_IN_DDR_F\);
    
    \U50_PATTERNS/ELINK_DINA_0[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119868, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_5, Q => 
        \U50_PATTERNS/ELINK_DINA_0[3]\);
    
    HIEFFPLA_INST_0_50852 : MX2
      port map(A => 
        \U_ELK8_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]_net_1\, B => 
        \U_ELK8_CH/ELK_TX_DAT[7]\, S => 
        \U_ELK8_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_117880);
    
    HIEFFPLA_INST_0_47625 : AND2A
      port map(A => \OP_MODE_c_2[1]\, B => \PATT_ELK_DAT_14[6]\, 
        Y => HIEFFPLA_NET_0_118457);
    
    HIEFFPLA_INST_0_41296 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_4[6]\, B => 
        HIEFFPLA_NET_0_119566, S => HIEFFPLA_NET_0_119284, Y => 
        HIEFFPLA_NET_0_119753);
    
    HIEFFPLA_INST_0_41233 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_3[7]\, B => 
        HIEFFPLA_NET_0_119560, S => HIEFFPLA_NET_0_119247, Y => 
        HIEFFPLA_NET_0_119760);
    
    HIEFFPLA_INST_0_49115 : NAND2B
      port map(A => \OP_MODE_c_5[1]\, B => \PATT_ELK_DAT_1[2]\, Y
         => HIEFFPLA_NET_0_118191);
    
    AFLSDF_INV_36 : INV
      port map(A => DCB_SALT_SEL_c, Y => \AFLSDF_INV_36\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_15[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116518, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_15, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_15[2]\);
    
    HIEFFPLA_INST_0_56556 : AND3
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[6]_net_1\, B => 
        HIEFFPLA_NET_0_117426, C => HIEFFPLA_NET_0_117425, Y => 
        HIEFFPLA_NET_0_116839);
    
    HIEFFPLA_INST_0_49539 : MX2
      port map(A => HIEFFPLA_NET_0_118132, B => 
        HIEFFPLA_NET_0_118115, S => \BIT_OS_SEL_1[0]\, Y => 
        \U_ELK2_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[7]\);
    
    \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[10]\ : DFN1C0
      port map(D => 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\);
    
    \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[1]\ : DFN1C0
      port map(D => 
        \U_ELK5_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[8]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[6]_net_1\, CLK => 
        CCC_160M_ADJ, CLR => P_MASTER_POR_B_c_34_0, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[8]_net_1\);
    
    \U_ELK8_CH/U_ELK1_SERDAT_SOURCE/SERDAT[7]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117871, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_5, Q => 
        \U_ELK8_CH/ELK_TX_DAT[7]\);
    
    \U50_PATTERNS/ELINK_ADDRA_8[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119949, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_8, Q => 
        \U50_PATTERNS/ELINK_ADDRA_8[2]\);
    
    \U50_PATTERNS/U4B_REGCROSS/SAMP_ONE[0]\ : DFN1C0
      port map(D => \U50_PATTERNS/TFC_STOP_ADDR[0]\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_24_0, Q => 
        \U50_PATTERNS/U4B_REGCROSS/SAMP_ONE[0]_net_1\);
    
    \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[14]\ : DFN1C0
      port map(D => \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[14]_net_1\);
    
    \U_ELK17_CH/U_SLAVE_1ELK/Q[10]\ : DFN1C0
      port map(D => \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/Q[10]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_28[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116055, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_15, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_28[0]\);
    
    HIEFFPLA_INST_0_53046 : MX2
      port map(A => HIEFFPLA_NET_0_117564, B => 
        HIEFFPLA_NET_0_117560, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[2]\, Y => 
        HIEFFPLA_NET_0_117472);
    
    \U_ELK10_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]\ : DFN1C0
      port map(D => \U_ELK10_CH/U_SLAVE_1ELK/Q[12]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]_net_1\);
    
    \U_ELK18_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]\ : DFN1C0
      port map(D => \U_ELK18_CH/U_SLAVE_1ELK/Q[12]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]_net_1\);
    
    HIEFFPLA_INST_0_47682 : MX2
      port map(A => HIEFFPLA_NET_0_118455, B => 
        HIEFFPLA_NET_0_118452, S => \BIT_OS_SEL_2[1]\, Y => 
        HIEFFPLA_NET_0_118447);
    
    HIEFFPLA_INST_0_41838 : OA1A
      port map(A => HIEFFPLA_NET_0_119235, B => 
        \U50_PATTERNS/ELINK_RWA[14]\, C => HIEFFPLA_NET_0_119656, 
        Y => HIEFFPLA_NET_0_119686);
    
    HIEFFPLA_INST_0_62689 : XNOR3
      port map(A => HIEFFPLA_NET_0_115960, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_CLKPHASE[1]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_SEQCNT[2]\, Y => 
        HIEFFPLA_NET_0_115957);
    
    HIEFFPLA_INST_0_59770 : MX2
      port map(A => HIEFFPLA_NET_0_116586, B => 
        HIEFFPLA_NET_0_116346, S => HIEFFPLA_NET_0_117357, Y => 
        HIEFFPLA_NET_0_116350);
    
    HIEFFPLA_INST_0_48366 : AND2A
      port map(A => \OP_MODE_c_6[1]\, B => \PATT_ELK_DAT_17[0]\, 
        Y => HIEFFPLA_NET_0_118328);
    
    HIEFFPLA_INST_0_46752 : MX2
      port map(A => HIEFFPLA_NET_0_118632, B => 
        HIEFFPLA_NET_0_118629, S => \BIT_OS_SEL_0[0]\, Y => 
        \U_ELK10_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[1]\);
    
    HIEFFPLA_INST_0_44791 : XO1
      port map(A => \U50_PATTERNS/U4E_REGCROSS/SAMP_TWO[4]_net_1\, 
        B => \OP_MODE[4]\, C => HIEFFPLA_NET_0_119047, Y => 
        HIEFFPLA_NET_0_119049);
    
    HIEFFPLA_INST_0_42342 : NAND2
      port map(A => \U50_PATTERNS/RD_USB_ADBUS[1]\, B => 
        \U50_PATTERNS/RD_USB_ADBUS[0]\, Y => 
        HIEFFPLA_NET_0_119565);
    
    \U_ELK5_CH/U_SLAVE_1ELK/Q[6]\ : DFN1C0
      port map(D => \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/Q[6]_net_1\);
    
    \U_ELK1_CH/U_SLAVE_1ELK/RECD_SER_WORD[4]\ : DFN1C0
      port map(D => \U_ELK1_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[4]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_1[4]\);
    
    HIEFFPLA_INST_0_63001 : AND3
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[9]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[10]\, C => 
        HIEFFPLA_NET_0_115915, Y => HIEFFPLA_NET_0_115919);
    
    HIEFFPLA_INST_0_42365 : AND2A
      port map(A => \U50_PATTERNS/RD_XFER_TYPE[1]_net_1\, B => 
        \U50_PATTERNS/RD_XFER_TYPE[0]_net_1\, Y => 
        HIEFFPLA_NET_0_119554);
    
    \U50_PATTERNS/U3_USB_DAT_BUS/_BIBUF_F_24U[1]_/U0/U1\ : 
        IOBI_IRC_OB_EB
      port map(D => \U50_PATTERNS/WR_USB_ADBUS[1]\, CLR => 
        \AFLSDF_INV_5\, E => \U50_PATTERNS/TrienAux\, ICLK => 
        CLK60MHZ, YIN => 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[1]\\\\/U0/NET3\, 
        DOUT => 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[1]\\\\/U0/NET1\, 
        EOUT => 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[1]\\\\/U0/NET2\, 
        Y => \U50_PATTERNS/RD_USB_ADBUS[1]\);
    
    HIEFFPLA_INST_0_54645 : AO1C
      port map(A => HIEFFPLA_NET_0_117219, B => 
        HIEFFPLA_NET_0_117116, C => HIEFFPLA_NET_0_117086, Y => 
        HIEFFPLA_NET_0_117228);
    
    HIEFFPLA_INST_0_43100 : AND2B
      port map(A => \U50_PATTERNS/REG_STATE[1]_net_1\, B => 
        \U50_PATTERNS/REG_STATE[0]_net_1\, Y => 
        HIEFFPLA_NET_0_119377);
    
    HIEFFPLA_INST_0_59880 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_3[0]\, B => 
        HIEFFPLA_NET_0_116680, S => HIEFFPLA_NET_0_117091, Y => 
        HIEFFPLA_NET_0_116339);
    
    \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[9]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117699, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_31, Q => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[9]_net_1\);
    
    \U50_PATTERNS/ELINK_ADDRA_11[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120073, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_2, Q => 
        \U50_PATTERNS/ELINK_ADDRA_11[6]\);
    
    HIEFFPLA_INST_0_61253 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_4[4]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_20[4]\, S
         => \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_5[4]_net_1\, 
        Y => HIEFFPLA_NET_0_116153);
    
    \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[37]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117714, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_33, Q => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[37]_net_1\);
    
    HIEFFPLA_INST_0_48580 : MX2
      port map(A => 
        \U_ELK18_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]_net_1\, B => 
        \U_ELK18_CH/ELK_TX_DAT[2]\, S => 
        \U_ELK18_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118291);
    
    HIEFFPLA_INST_0_51505 : AND3
      port map(A => \U_EXEC_MASTER/CCC_1_LOCK_STAT_1D_net_1\, B
         => HIEFFPLA_NET_0_117764, C => HIEFFPLA_NET_0_117760, Y
         => HIEFFPLA_NET_0_117761);
    
    \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[9]\ : DFN1C0
      port map(D => \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\);
    
    \U_ELK14_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118470, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_5, Q => 
        \U_ELK14_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]_net_1\);
    
    \U63_TS_SIWU_BUF/\\\\TRIBUFF_F_24U[0]\\\\/U0/U0\ : 
        IOPAD_TRI_U
      port map(D => 
        \U63_TS_SIWU_BUF/\\\\TRIBUFF_F_24U[0]\\\\/U0/NET1\, E => 
        \U63_TS_SIWU_BUF/\\\\TRIBUFF_F_24U[0]\\\\/U0/NET2\, PAD
         => USB_SIWU_B);
    
    HIEFFPLA_INST_0_61040 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_2[0]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_18[0]\, S
         => \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_4[4]_net_1\, 
        Y => HIEFFPLA_NET_0_116181);
    
    \U_MASTER_DES/U13C_MASTER_DESER/RECD_SER_WORD[5]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_116899, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_30, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/RECD_SER_WORD[5]_net_1\);
    
    HIEFFPLA_INST_0_55127 : NAND3C
      port map(A => HIEFFPLA_NET_0_117123, B => 
        HIEFFPLA_NET_0_117339, C => HIEFFPLA_NET_0_117110, Y => 
        HIEFFPLA_NET_0_117116);
    
    \U_ELK4_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL\ : DFN1C0
      port map(D => 
        \U_ELK4_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL_net_1\);
    
    HIEFFPLA_INST_0_57160 : XA1B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_2[7]\, B => 
        HIEFFPLA_NET_0_116737, C => HIEFFPLA_NET_0_117179, Y => 
        HIEFFPLA_NET_0_116728);
    
    HIEFFPLA_INST_0_45618 : NAND3C
      port map(A => HIEFFPLA_NET_0_118713, B => 
        HIEFFPLA_NET_0_118723, C => HIEFFPLA_NET_0_118731, Y => 
        HIEFFPLA_NET_0_118879);
    
    HIEFFPLA_INST_0_45399 : NAND2A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_19[2]\, Y => 
        HIEFFPLA_NET_0_118921);
    
    \U_ELK16_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]\ : DFN1C0
      port map(D => \U_ELK16_CH/U_SLAVE_1ELK/Q[5]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]_net_1\);
    
    \U50_PATTERNS/U4D_REGCROSS/DELCNT[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119073, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_26, Q => 
        \U50_PATTERNS/U4D_REGCROSS/DELCNT[1]_net_1\);
    
    \U50_PATTERNS/ELINK_ADDRA_18[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120023, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_12, Q => 
        \U50_PATTERNS/ELINK_ADDRA_18[0]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_27[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116391, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_2, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_27[3]\);
    
    HIEFFPLA_INST_0_55196 : AND2B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[8]_net_1\, B => 
        HIEFFPLA_NET_0_117338, Y => HIEFFPLA_NET_0_117096);
    
    \U50_PATTERNS/TFC_DINA[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119193, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_4, Q => \U50_PATTERNS/TFC_DINA[4]\);
    
    HIEFFPLA_INST_0_161270 : DFN1C0
      port map(D => \U_ELK16_CH/ELK_TX_DAT[7]\, CLK => 
        CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_10, Q => 
        HIEFFPLA_NET_0_161285);
    
    \U200A_TFC/RX_SER_WORD_1DEL[4]\ : DFN1C0
      port map(D => \TFC_RX_SER_WORD[4]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_31, Q => 
        \U200A_TFC/RX_SER_WORD_1DEL[4]_net_1\);
    
    HIEFFPLA_INST_0_47098 : MX2
      port map(A => 
        \U_ELK12_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]_net_1\, B => 
        \U_ELK12_CH/ELK_TX_DAT[6]\, S => 
        \U_ELK12_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118559);
    
    HIEFFPLA_INST_0_39002 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_16[0]\, B => 
        HIEFFPLA_NET_0_119524, S => HIEFFPLA_NET_0_119257, Y => 
        HIEFFPLA_NET_0_120039);
    
    \U50_PATTERNS/U4D_REGCROSS/LOCAL_REG_VAL[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119090, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_3, Q => \ELKS_STOP_ADDR[1]\);
    
    \U_ELK7_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL\ : DFN1C0
      port map(D => \U_ELK7_CH/ELK_IN_F_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL_net_1\);
    
    HIEFFPLA_INST_0_62203 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_14[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_30[1]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[4]_net_1\, Y => 
        HIEFFPLA_NET_0_116023);
    
    HIEFFPLA_INST_0_50361 : NAND2B
      port map(A => \OP_MODE_c_0[1]\, B => \PATT_ELK_DAT_6[3]\, Y
         => HIEFFPLA_NET_0_117965);
    
    AFLSDF_INV_51 : INV
      port map(A => DCB_SALT_SEL_c, Y => \AFLSDF_INV_51\);
    
    HIEFFPLA_INST_0_56234 : AND2
      port map(A => DCB_SALT_SEL_c, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/RECD_SER_WORD[0]_net_1\, 
        Y => \ELK_RX_SER_WORD_0[0]\);
    
    HIEFFPLA_INST_0_55201 : AND3A
      port map(A => HIEFFPLA_NET_0_117247, B => 
        HIEFFPLA_NET_0_117242, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[6]_net_1\, Y => 
        HIEFFPLA_NET_0_117094);
    
    HIEFFPLA_INST_0_50053 : MX2
      port map(A => HIEFFPLA_NET_0_118039, B => 
        HIEFFPLA_NET_0_118023, S => \BIT_OS_SEL_0[1]\, Y => 
        HIEFFPLA_NET_0_118025);
    
    HIEFFPLA_INST_0_47740 : MX2
      port map(A => HIEFFPLA_NET_0_118431, B => 
        HIEFFPLA_NET_0_118447, S => \BIT_OS_SEL_4[0]\, Y => 
        \U_ELK14_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[0]\);
    
    \U50_PATTERNS/U4E_REGCROSS/LOCAL_REG_VAL_1[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119061, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_1, Q => \OP_MODE_c_1[1]\);
    
    HIEFFPLA_INST_0_46324 : NAND3C
      port map(A => HIEFFPLA_NET_0_119618, B => 
        HIEFFPLA_NET_0_119623, C => HIEFFPLA_NET_0_118882, Y => 
        HIEFFPLA_NET_0_118717);
    
    \U_MASTER_DES/U13C_MASTER_DESER/ARB_WRD_40M_FIXED[4]\ : 
        DFN1C0
      port map(D => \U_MASTER_DES/U13C_MASTER_DESER/Q[4]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_26, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_WRD_40M_FIXED[4]_net_1\);
    
    \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[6]\ : DFN1C0
      port map(D => 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\);
    
    HIEFFPLA_INST_0_45854 : AO1
      port map(A => HIEFFPLA_NET_0_119283, B => 
        \U50_PATTERNS/ELINK_DOUTA_13[1]\, C => 
        HIEFFPLA_NET_0_118780, Y => HIEFFPLA_NET_0_118827);
    
    \U_TFC_CMD_TX/SER_OUT_RDEL\ : DFN1C0
      port map(D => \U_TFC_CMD_TX/SER_OUT_RI_net_1\, CLK => 
        CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        TFC_OUT_R);
    
    \U50_PATTERNS/U4D_REGCROSS/SAMP_TWO[6]\ : DFN1C0
      port map(D => \U50_PATTERNS/U4D_REGCROSS/SAMP_ONE[6]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_30, Q => 
        \U50_PATTERNS/U4D_REGCROSS/SAMP_TWO[6]_net_1\);
    
    HIEFFPLA_INST_0_57467 : AND3A
      port map(A => HIEFFPLA_NET_0_116686, B => 
        HIEFFPLA_NET_0_116708, C => HIEFFPLA_NET_0_116620, Y => 
        HIEFFPLA_NET_0_116676);
    
    \U_ELK11_CH/U_ELK1_CMD_TX/SER_OUT_RI\ : DFN1C0
      port map(D => 
        \U_ELK11_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_2, Q => 
        \U_ELK11_CH/U_ELK1_CMD_TX/SER_OUT_RI_net_1\);
    
    HIEFFPLA_INST_0_50362 : AND2A
      port map(A => \OP_MODE_c_0[1]\, B => \PATT_ELK_DAT_6[4]\, Y
         => HIEFFPLA_NET_0_117964);
    
    HIEFFPLA_INST_0_46553 : MX2
      port map(A => HIEFFPLA_NET_0_118667, B => \ELK0_TX_DAT[6]\, 
        S => \U_ELK0_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118666);
    
    HIEFFPLA_INST_0_39641 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_5[7]\, B => 
        HIEFFPLA_NET_0_119516, S => HIEFFPLA_NET_0_119251, Y => 
        HIEFFPLA_NET_0_119968);
    
    \U_ELK6_CH/U_SLAVE_1ELK/Q[8]\ : DFN1C0
      port map(D => \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/Q[8]_net_1\);
    
    \U_ELK3_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]\ : DFN1C0
      port map(D => \U_ELK3_CH/U_SLAVE_1ELK/Q[10]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]_net_1\);
    
    HIEFFPLA_INST_0_61490 : MX2
      port map(A => HIEFFPLA_NET_0_117167, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_23[1]\, S => 
        HIEFFPLA_NET_0_117151, Y => HIEFFPLA_NET_0_116119);
    
    HIEFFPLA_INST_0_50067 : MX2
      port map(A => \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\, 
        B => \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[14]_net_1\, S => 
        \BIT_OS_SEL[2]\, Y => HIEFFPLA_NET_0_118023);
    
    HIEFFPLA_INST_0_50883 : MX2
      port map(A => HIEFFPLA_NET_0_117864, B => 
        HIEFFPLA_NET_0_117862, S => \BIT_OS_SEL_3[1]\, Y => 
        HIEFFPLA_NET_0_117868);
    
    HIEFFPLA_INST_0_39857 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_8[7]\, B => 
        HIEFFPLA_NET_0_119516, S => HIEFFPLA_NET_0_119291, Y => 
        HIEFFPLA_NET_0_119944);
    
    \U50_PATTERNS/ELINK_ADDRA_1[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120004, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_20, Q => 
        \U50_PATTERNS/ELINK_ADDRA_1[3]\);
    
    HIEFFPLA_INST_0_55152 : AO1
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[8]_net_1\, B => 
        \OP_MODE_c[5]\, C => HIEFFPLA_NET_0_117068, Y => 
        HIEFFPLA_NET_0_117111);
    
    \U_EXEC_MASTER/MPOR_DCB_B\ : DFI1P0
      port map(D => HIEFFPLA_NET_0_117769, CLK => CLK_40M_GL, PRE
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i\, QN => 
        \U_EXEC_MASTER/MPOR_DCB_B_net_1\);
    
    \U_ELK13_CH/U_SLAVE_1ELK/Q[11]\ : DFN1C0
      port map(D => \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/Q[11]_net_1\);
    
    HIEFFPLA_INST_0_37758 : AOI1
      port map(A => \U200B_ELINKS/GP_PG_SM[0]_net_1\, B => 
        HIEFFPLA_NET_0_120204, C => HIEFFPLA_NET_0_120197, Y => 
        HIEFFPLA_NET_0_120214);
    
    \U_ELK9_CH/U_SLAVE_1ELK/Q[11]\ : DFN1C0
      port map(D => \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/Q[11]_net_1\);
    
    \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[2]\ : DFN1C0
      port map(D => 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[2]_net_1\);
    
    \U200A_TFC/RX_SER_WORD_3DEL[2]\ : DFN1P0
      port map(D => \AFLSDF_INV_53\, CLK => CLK_40M_GL, PRE => 
        P_MASTER_POR_B_c_24, Q => 
        \U200A_TFC/RX_SER_WORD_3DEL_i_0[2]\);
    
    HIEFFPLA_INST_0_56809 : XA1C
      port map(A => HIEFFPLA_NET_0_116789, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_0[8]\, C => 
        HIEFFPLA_NET_0_117179, Y => HIEFFPLA_NET_0_116792);
    
    HIEFFPLA_INST_0_59936 : MX2
      port map(A => HIEFFPLA_NET_0_116687, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_3[2]\, S => 
        HIEFFPLA_NET_0_117207, Y => HIEFFPLA_NET_0_116331);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_5[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_115993, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_15, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_5[2]\);
    
    HIEFFPLA_INST_0_57087 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_2[8]\, B => 
        HIEFFPLA_NET_0_116727, S => HIEFFPLA_NET_0_117601, Y => 
        HIEFFPLA_NET_0_116747);
    
    HIEFFPLA_INST_0_55898 : MX2
      port map(A => HIEFFPLA_NET_0_116964, B => 
        HIEFFPLA_NET_0_116988, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[1]\, Y => 
        HIEFFPLA_NET_0_116976);
    
    HIEFFPLA_INST_0_49365 : NAND2B
      port map(A => \OP_MODE_c_1[1]\, B => \PATT_ELK_DAT_2[3]\, Y
         => HIEFFPLA_NET_0_118145);
    
    HIEFFPLA_INST_0_39758 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_7[4]\, B => 
        HIEFFPLA_NET_0_119519, S => HIEFFPLA_NET_0_119289, Y => 
        HIEFFPLA_NET_0_119955);
    
    HIEFFPLA_INST_0_43139 : AO1A
      port map(A => HIEFFPLA_NET_0_119387, B => 
        HIEFFPLA_NET_0_119347, C => HIEFFPLA_NET_0_119349, Y => 
        HIEFFPLA_NET_0_119362);
    
    HIEFFPLA_INST_0_63159 : XOR2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[1]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[0]\, Y => 
        HIEFFPLA_NET_0_115872);
    
    \U_TFC_CMD_TX/SER_OUT_FI\ : DFN1C0
      port map(D => \U_TFC_CMD_TX/SER_CMD_WORD_F[3]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_TFC_CMD_TX/SER_OUT_FI_net_1\);
    
    \U_ELK10_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118647, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_3, Q => 
        \U_ELK10_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]_net_1\);
    
    \U_ELK6_CH/U_SLAVE_1ELK/Q[4]\ : DFN1C0
      port map(D => \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/Q[4]_net_1\);
    
    HIEFFPLA_INST_0_44633 : XO1
      port map(A => \U50_PATTERNS/U4D_REGCROSS/SAMP_TWO[0]_net_1\, 
        B => \ELKS_STOP_ADDR[0]\, C => HIEFFPLA_NET_0_119076, Y
         => HIEFFPLA_NET_0_119080);
    
    \U50_PATTERNS/U4C_REGCROSS/LOCAL_REG_VAL[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119112, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_21, Q => \ELKS_STRT_ADDR[0]\);
    
    \U50_PATTERNS/ELINK_DINA_4[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119754, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_13, Q => 
        \U50_PATTERNS/ELINK_DINA_4[5]\);
    
    HIEFFPLA_INST_0_57687 : AOI1
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_5[0]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_5[1]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_5[2]\, Y => 
        HIEFFPLA_NET_0_116635);
    
    HIEFFPLA_INST_0_46263 : AO1
      port map(A => HIEFFPLA_NET_0_119476, B => 
        \U50_PATTERNS/CHKSUM[4]\, C => HIEFFPLA_NET_0_118901, Y
         => HIEFFPLA_NET_0_118729);
    
    HIEFFPLA_INST_0_43042 : OR3B
      port map(A => HIEFFPLA_NET_0_119600, B => 
        HIEFFPLA_NET_0_119586, C => HIEFFPLA_NET_0_119581, Y => 
        HIEFFPLA_NET_0_119394);
    
    HIEFFPLA_INST_0_46718 : MX2
      port map(A => \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[1]_net_1\, 
        B => \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\, S => 
        \BIT_OS_SEL_5[2]\, Y => HIEFFPLA_NET_0_118623);
    
    HIEFFPLA_INST_0_56834 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_1[1]\, B => 
        HIEFFPLA_NET_0_116767, S => HIEFFPLA_NET_0_117600, Y => 
        HIEFFPLA_NET_0_116787);
    
    HIEFFPLA_INST_0_59621 : MX2
      port map(A => HIEFFPLA_NET_0_116687, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_29[2]\, S => 
        HIEFFPLA_NET_0_117395, Y => HIEFFPLA_NET_0_116369);
    
    HIEFFPLA_INST_0_52526 : MX2
      port map(A => HIEFFPLA_NET_0_117492, B => 
        HIEFFPLA_NET_0_117488, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_2[3]\, Y => 
        HIEFFPLA_NET_0_117552);
    
    HIEFFPLA_INST_0_52134 : NAND3A
      port map(A => HIEFFPLA_NET_0_117624, B => 
        HIEFFPLA_NET_0_117626, C => HIEFFPLA_NET_0_117623, Y => 
        HIEFFPLA_NET_0_117629);
    
    HIEFFPLA_INST_0_38434 : MX2
      port map(A => \U50_PATTERNS/ELINKS_STRT_ADDR_T[0]\, B => 
        \U50_PATTERNS/RD_USB_ADBUS[0]\, S => 
        HIEFFPLA_NET_0_119493, Y => HIEFFPLA_NET_0_120103);
    
    HIEFFPLA_INST_0_57648 : AND3B
      port map(A => HIEFFPLA_NET_0_117085, B => 
        HIEFFPLA_NET_0_116635, C => HIEFFPLA_NET_0_116650, Y => 
        HIEFFPLA_NET_0_116643);
    
    HIEFFPLA_INST_0_47555 : MX2
      port map(A => HIEFFPLA_NET_0_118474, B => 
        HIEFFPLA_NET_0_118500, S => \BIT_OS_SEL_3[1]\, Y => 
        HIEFFPLA_NET_0_118476);
    
    HIEFFPLA_INST_0_39083 : MX2
      port map(A => HIEFFPLA_NET_0_119523, B => 
        \U50_PATTERNS/ELINK_ADDRA_17[1]\, S => 
        HIEFFPLA_NET_0_119260, Y => HIEFFPLA_NET_0_120030);
    
    HIEFFPLA_INST_0_39650 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_6[0]\, B => 
        HIEFFPLA_NET_0_119524, S => HIEFFPLA_NET_0_119258, Y => 
        HIEFFPLA_NET_0_119967);
    
    \U_EXEC_MASTER/MPOR_B_3\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117787, CLK => CLK_40M_GL, CLR
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_2\, Q => 
        P_MASTER_POR_B_c_3);
    
    \U_ELK16_CH/U_SLAVE_1ELK/Q[13]\ : DFN1C0
      port map(D => \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[13]_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/Q[13]_net_1\);
    
    HIEFFPLA_INST_0_59193 : MX2B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_24[3]\, B => 
        HIEFFPLA_NET_0_116774, S => HIEFFPLA_NET_0_117208, Y => 
        HIEFFPLA_NET_0_116422);
    
    HIEFFPLA_INST_0_44525 : XO1
      port map(A => \U50_PATTERNS/U4C_REGCROSS/SAMP_TWO[2]_net_1\, 
        B => \ELKS_STRT_ADDR[2]\, C => HIEFFPLA_NET_0_119098, Y
         => HIEFFPLA_NET_0_119102);
    
    HIEFFPLA_INST_0_56880 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_1[6]\, B => 
        HIEFFPLA_NET_0_116761, S => HIEFFPLA_NET_0_117600, Y => 
        HIEFFPLA_NET_0_116782);
    
    HIEFFPLA_INST_0_42693 : AOI1D
      port map(A => HIEFFPLA_NET_0_119396, B => 
        HIEFFPLA_NET_0_119465, C => HIEFFPLA_NET_0_119558, Y => 
        HIEFFPLA_NET_0_119481);
    
    \U_ELK18_CH/U_SLAVE_1ELK/Q[9]\ : DFN1C0
      port map(D => \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/Q[9]_net_1\);
    
    HIEFFPLA_INST_0_46492 : AND3C
      port map(A => \U50_PATTERNS/RD_USB_ADBUS[2]\, B => 
        HIEFFPLA_NET_0_119596, C => HIEFFPLA_NET_0_119571, Y => 
        HIEFFPLA_NET_0_118679);
    
    HIEFFPLA_INST_0_49555 : MX2
      port map(A => HIEFFPLA_NET_0_118128, B => 
        HIEFFPLA_NET_0_118113, S => \BIT_OS_SEL_1[1]\, Y => 
        HIEFFPLA_NET_0_118115);
    
    HIEFFPLA_INST_0_47967 : MX2
      port map(A => \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\, 
        B => \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[13]_net_1\, S => 
        \BIT_OS_SEL_2[2]\, Y => HIEFFPLA_NET_0_118397);
    
    HIEFFPLA_INST_0_161276 : DFN1C0
      port map(D => \ELK0_TX_DAT[4]\, CLK => CCC_160M_FXD, CLR
         => MASTER_SALT_POR_B_i_0_i_17, Q => 
        HIEFFPLA_NET_0_161279);
    
    HIEFFPLA_INST_0_46868 : MX2
      port map(A => 
        \U_ELK11_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]_net_1\, B => 
        \U_ELK11_CH/ELK_TX_DAT[7]\, S => 
        \U_ELK11_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118600);
    
    HIEFFPLA_INST_0_54586 : MX2
      port map(A => HIEFFPLA_NET_0_116497, B => 
        HIEFFPLA_NET_0_116278, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[3]_net_1\, Y => 
        HIEFFPLA_NET_0_117239);
    
    HIEFFPLA_INST_0_42656 : OA1A
      port map(A => HIEFFPLA_NET_0_119379, B => 
        HIEFFPLA_NET_0_119471, C => HIEFFPLA_NET_0_119393, Y => 
        HIEFFPLA_NET_0_119490);
    
    HIEFFPLA_INST_0_37175 : AND3C
      port map(A => \U200A_TFC/GP_PG_SM[6]_net_1\, B => 
        \U200A_TFC/GP_PG_SM[7]_net_1\, C => 
        \U200A_TFC/GP_PG_SM[8]_net_1\, Y => HIEFFPLA_NET_0_120333);
    
    HIEFFPLA_INST_0_54582 : AND3B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[3]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[1]_net_1\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[0]_net_1\, Y => 
        HIEFFPLA_NET_0_117240);
    
    HIEFFPLA_INST_0_42722 : NAND3
      port map(A => HIEFFPLA_NET_0_119431, B => 
        HIEFFPLA_NET_0_119371, C => 
        \U50_PATTERNS/REG_STATE_0[1]_net_1\, Y => 
        HIEFFPLA_NET_0_119475);
    
    \U_ELK4_CH/U_SLAVE_1ELK/Q[11]\ : DFN1C0
      port map(D => \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/Q[11]_net_1\);
    
    \U_ELK15_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118422, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_6, Q => 
        \U_ELK15_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]_net_1\);
    
    HIEFFPLA_INST_0_45988 : NAND2B
      port map(A => HIEFFPLA_NET_0_118795, B => 
        HIEFFPLA_NET_0_118696, Y => HIEFFPLA_NET_0_118796);
    
    \U_ELK11_CH/U_SLAVE_1ELK/Q[1]\ : DFN1C0
      port map(D => \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/Q[1]_net_1\);
    
    HIEFFPLA_INST_0_37072 : XO1A
      port map(A => HIEFFPLA_NET_0_120334, B => \TFC_ADDRB[0]\, C
         => \U200A_TFC/GP_PG_SM[10]_net_1\, Y => 
        HIEFFPLA_NET_0_120353);
    
    HIEFFPLA_INST_0_43377 : MX2
      port map(A => \U50_PATTERNS/SM_BANK_SEL[13]\, B => 
        HIEFFPLA_NET_0_119224, S => HIEFFPLA_NET_0_118691, Y => 
        HIEFFPLA_NET_0_119318);
    
    HIEFFPLA_INST_0_42581 : XA1B
      port map(A => \U50_PATTERNS/REG_ADDR[2]\, B => 
        HIEFFPLA_NET_0_119500, C => HIEFFPLA_NET_0_119452, Y => 
        HIEFFPLA_NET_0_119507);
    
    \U_ELK7_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]\ : DFN1C0
      port map(D => \U_ELK7_CH/U_SLAVE_1ELK/Q[12]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]_net_1\);
    
    \U200A_TFC/RX_SER_WORD_2DEL[1]\ : DFN1C0
      port map(D => \U200A_TFC/RX_SER_WORD_1DEL[1]_net_1\, CLK
         => CLK_40M_GL, CLR => P_MASTER_POR_B_c, Q => 
        \U200A_TFC/RX_SER_WORD_2DEL[1]_net_1\);
    
    HIEFFPLA_INST_0_49618 : NAND2B
      port map(A => \OP_MODE_c_5[1]\, B => \PATT_ELK_DAT_3[7]\, Y
         => HIEFFPLA_NET_0_118096);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_20[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116157, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_2, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_20[3]\);
    
    \U_ELK10_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]\ : DFN1C0
      port map(D => \U_ELK10_CH/U_SLAVE_1ELK/Q[14]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]_net_1\);
    
    HIEFFPLA_INST_0_57621 : NAND3
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_5[0]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_5[2]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_5[1]\, Y => 
        HIEFFPLA_NET_0_116650);
    
    HIEFFPLA_INST_0_55078 : AND3
      port map(A => HIEFFPLA_NET_0_117603, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[7]_net_1\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[6]_net_1\, Y => 
        HIEFFPLA_NET_0_117126);
    
    \U_ELK7_CH/U_ELK1_SERDAT_SOURCE/SERDAT[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117920, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_3, Q => 
        \U_ELK7_CH/ELK_TX_DAT[3]\);
    
    \U_ELK2_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]\ : DFN1C0
      port map(D => \U_ELK2_CH/U_SLAVE_1ELK/Q[8]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]_net_1\);
    
    \U_ELK18_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]\ : DFN1C0
      port map(D => \U_ELK18_CH/U_SLAVE_1ELK/Q[14]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]_net_1\);
    
    HIEFFPLA_INST_0_59202 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_24[0]\, B => 
        HIEFFPLA_NET_0_116774, S => HIEFFPLA_NET_0_117208, Y => 
        HIEFFPLA_NET_0_116421);
    
    \U_MASTER_DES/U13C_MASTER_DESER/ADJ_SER_IN_F_1DEL\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117611, CLK => CCC_160M_ADJ, 
        CLR => P_MASTER_POR_B_c_32, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_SER_IN_F_1DEL_net_1\);
    
    HIEFFPLA_INST_0_57769 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_6[7]\, B => 
        HIEFFPLA_NET_0_116608, S => HIEFFPLA_NET_0_117599, Y => 
        HIEFFPLA_NET_0_116625);
    
    \U_ELK6_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117972, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_6, Q => 
        \U_ELK6_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]_net_1\);
    
    \U_ELK1_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]\ : DFN1C0
      port map(D => \U_ELK1_CH/U_SLAVE_1ELK/Q[11]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]_net_1\);
    
    \U50_PATTERNS/ELINK_DINA_19[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119786, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_1, Q => 
        \U50_PATTERNS/ELINK_DINA_19[5]\);
    
    HIEFFPLA_INST_0_45637 : NAND3C
      port map(A => HIEFFPLA_NET_0_118900, B => 
        HIEFFPLA_NET_0_118728, C => HIEFFPLA_NET_0_118875, Y => 
        HIEFFPLA_NET_0_118876);
    
    \U_ELK8_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL\ : DFN1C0
      port map(D => \U_ELK8_CH/ELK_IN_R_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL_net_1\);
    
    \U_ELK18_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]\ : DFN1C0
      port map(D => \U_ELK18_CH/U_SLAVE_1ELK/Q[9]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]_net_1\);
    
    HIEFFPLA_INST_0_53030 : MX2
      port map(A => HIEFFPLA_NET_0_117454, B => 
        HIEFFPLA_NET_0_117566, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[2]\, Y => 
        HIEFFPLA_NET_0_117474);
    
    HIEFFPLA_INST_0_39987 : MX2
      port map(A => HIEFFPLA_NET_0_119902, B => 
        \U50_PATTERNS/ELINK_BLKA[16]\, S => 
        \U50_PATTERNS/SM_BANK_SEL[20]\, Y => 
        HIEFFPLA_NET_0_119928);
    
    HIEFFPLA_INST_0_53313 : AND3C
      port map(A => \BIT_OS_SEL_1[2]\, B => \BIT_OS_SEL_1[0]\, C
         => \BIT_OS_SEL_1[1]\, Y => HIEFFPLA_NET_0_117432);
    
    HIEFFPLA_INST_0_48792 : MX2
      port map(A => HIEFFPLA_NET_0_118275, B => 
        HIEFFPLA_NET_0_118250, S => \BIT_OS_SEL_2[0]\, Y => 
        \U_ELK18_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[7]\);
    
    HIEFFPLA_INST_0_47812 : MX2
      port map(A => HIEFFPLA_NET_0_118444, B => 
        HIEFFPLA_NET_0_118428, S => \BIT_OS_SEL_4[1]\, Y => 
        HIEFFPLA_NET_0_118430);
    
    \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[8]\ : DFN1C0
      port map(D => \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\);
    
    HIEFFPLA_INST_0_51057 : MX2
      port map(A => \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[0]_net_1\, B
         => \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\, S => 
        \BIT_OS_SEL_3[2]\, Y => HIEFFPLA_NET_0_117844);
    
    HIEFFPLA_INST_0_49997 : MX2
      port map(A => HIEFFPLA_NET_0_118035, B => 
        HIEFFPLA_NET_0_118049, S => \BIT_OS_SEL_0[0]\, Y => 
        \U_ELK4_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[2]\);
    
    HIEFFPLA_INST_0_63237 : AND2A
      port map(A => \OP_MODE_c_0[1]\, B => \PATT_TFC_DAT[0]\, Y
         => \U_TFC_SERDAT_SOURCE/N_SERDAT[0]\);
    
    HIEFFPLA_INST_0_50142 : MX2
      port map(A => HIEFFPLA_NET_0_118000, B => 
        HIEFFPLA_NET_0_117998, S => \BIT_OS_SEL_6[1]\, Y => 
        HIEFFPLA_NET_0_118002);
    
    \U_MASTER_DES/U13C_MASTER_DESER/ADJ_SER_IN_R_1DEL\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117610, CLK => CCC_160M_ADJ, 
        CLR => P_MASTER_POR_B_c_27_1, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_SER_IN_R_1DEL_net_1\);
    
    \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[31]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117716, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_33, Q => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[31]_net_1\);
    
    HIEFFPLA_INST_0_50859 : NAND2B
      port map(A => \OP_MODE_c_0[1]\, B => \PATT_ELK_DAT_8[3]\, Y
         => HIEFFPLA_NET_0_117875);
    
    \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_SEL[3]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_BIT_OS_VAL[3]\, CLK
         => CLK_40M_GL, CLR => P_MASTER_POR_B_c_27_1, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_SEL[3]_net_1\);
    
    \U50_PATTERNS/ELINK_DINA_5[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119747, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_14, Q => 
        \U50_PATTERNS/ELINK_DINA_5[4]\);
    
    HIEFFPLA_INST_0_62030 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_29[1]\, B => 
        HIEFFPLA_NET_0_117114, S => HIEFFPLA_NET_0_117072, Y => 
        HIEFFPLA_NET_0_116044);
    
    HIEFFPLA_INST_0_55379 : NAND3
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[2]_net_1\, B => 
        \U_MASTER_DES/CCC_RX_CLK_LOCK\, C => 
        HIEFFPLA_NET_0_115918, Y => HIEFFPLA_NET_0_117046);
    
    \U_TFC_SERDAT_SOURCE/SERDAT[2]\ : DFN1C0
      port map(D => \U_TFC_SERDAT_SOURCE/N_SERDAT[2]\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \TFC_TX_DAT[2]\);
    
    \U_ELK17_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118337, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_17, Q => 
        \U_ELK17_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]_net_1\);
    
    HIEFFPLA_INST_0_55648 : AO1
      port map(A => HIEFFPLA_NET_0_117087, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_2[3]\, C => 
        HIEFFPLA_NET_0_117008, Y => HIEFFPLA_NET_0_117009);
    
    HIEFFPLA_INST_0_47603 : MX2
      port map(A => 
        \U_ELK14_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]_net_1\, B => 
        \U_ELK14_CH/ELK_TX_DAT[3]\, S => 
        \U_ELK14_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118467);
    
    HIEFFPLA_INST_0_44518 : NAND3C
      port map(A => HIEFFPLA_NET_0_119100, B => 
        HIEFFPLA_NET_0_119101, C => HIEFFPLA_NET_0_119102, Y => 
        HIEFFPLA_NET_0_119103);
    
    HIEFFPLA_INST_0_61376 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_21[2]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_22[2]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_3[0]\, Y => 
        HIEFFPLA_NET_0_116135);
    
    HIEFFPLA_INST_0_42523 : OA1A
      port map(A => HIEFFPLA_NET_0_119433, B => 
        HIEFFPLA_NET_0_119010, C => \U50_PATTERNS/REG_ADDR[2]\, Y
         => HIEFFPLA_NET_0_119522);
    
    \U_ELK3_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118112, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_16, Q => 
        \U_ELK3_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]_net_1\);
    
    HIEFFPLA_INST_0_50335 : MX2
      port map(A => 
        \U_ELK6_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]_net_1\, B => 
        \U_ELK6_CH/ELK_TX_DAT[6]\, S => 
        \U_ELK6_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_117974);
    
    \U_EXEC_MASTER/MPOR_DCB_B_RNIPFG8\ : CLKINT
      port map(A => \U_EXEC_MASTER/MPOR_DCB_B_net_1\, Y => 
        MASTER_DCB_POR_B_i_0_i);
    
    HIEFFPLA_INST_0_52630 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_13[0]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_14[0]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_2[0]\, Y => 
        HIEFFPLA_NET_0_117536);
    
    HIEFFPLA_INST_0_47435 : MX2
      port map(A => HIEFFPLA_NET_0_118493, B => 
        HIEFFPLA_NET_0_118489, S => \BIT_OS_SEL_3[1]\, Y => 
        HIEFFPLA_NET_0_118492);
    
    HIEFFPLA_INST_0_41197 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_3[3]\, B => 
        HIEFFPLA_NET_0_119574, S => HIEFFPLA_NET_0_119247, Y => 
        HIEFFPLA_NET_0_119764);
    
    HIEFFPLA_INST_0_52370 : MX2
      port map(A => HIEFFPLA_NET_0_117528, B => 
        HIEFFPLA_NET_0_117484, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[1]\, Y => 
        HIEFFPLA_NET_0_117572);
    
    HIEFFPLA_INST_0_52007 : MX2C
      port map(A => \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[48]\, B
         => \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[49]\, S => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[0]\, Y => 
        HIEFFPLA_NET_0_117654);
    
    \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[13]\ : DFN1C0
      port map(D => \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\, 
        CLK => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[13]_net_1\);
    
    \U_EXEC_MASTER/USB_MASTER_EN/T_CNT60M[6]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117737, CLK => CLK60MHZ, CLR
         => P_MASTER_POR_B_c_28, Q => 
        \U_EXEC_MASTER/USB_MASTER_EN/T_CNT60M[6]_net_1\);
    
    HIEFFPLA_INST_0_45592 : AO1A
      port map(A => HIEFFPLA_NET_0_119428, B => 
        \U50_PATTERNS/ELINKS_STRT_ADDR[5]\, C => 
        HIEFFPLA_NET_0_118789, Y => HIEFFPLA_NET_0_118884);
    
    HIEFFPLA_INST_0_45502 : AND3A
      port map(A => HIEFFPLA_NET_0_119437, B => 
        \U50_PATTERNS/WR_XFER_TYPE[4]_net_1\, C => 
        HIEFFPLA_NET_0_119367, Y => HIEFFPLA_NET_0_118901);
    
    \U50_PATTERNS/ELINK_ADDRA_10[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120081, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_22, Q => 
        \U50_PATTERNS/ELINK_ADDRA_10[6]\);
    
    HIEFFPLA_INST_0_51160 : MX2
      port map(A => \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[2]_net_1\, B
         => \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\, S => 
        \BIT_OS_SEL_2[2]\, Y => HIEFFPLA_NET_0_117819);
    
    \U_EXEC_MASTER/MPOR_B_6\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117787, CLK => CLK_40M_GL, CLR
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_1\, Q => 
        P_MASTER_POR_B_c_6);
    
    \U_ELK13_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118512, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_16, Q => 
        \U_ELK13_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]_net_1\);
    
    HIEFFPLA_INST_0_48875 : MX2
      port map(A => HIEFFPLA_NET_0_118220, B => 
        HIEFFPLA_NET_0_118217, S => \BIT_OS_SEL_0[1]\, Y => 
        HIEFFPLA_NET_0_118230);
    
    \U_ELK19_CH/U_SLAVE_1ELK/RECD_SER_WORD[4]\ : DFN1C0
      port map(D => \U_ELK19_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[4]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_19[4]\);
    
    HIEFFPLA_INST_0_44931 : AND3A
      port map(A => \U50_PATTERNS/REG_STATE[5]_net_1\, B => 
        \U50_PATTERNS/REG_STATE[2]_net_1\, C => 
        \U50_PATTERNS/USB_RXF_B\, Y => HIEFFPLA_NET_0_119014);
    
    \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_SEL[1]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_BIT_OS_VAL[1]\, CLK
         => CLK_40M_GL, CLR => P_MASTER_POR_B_c_27_1, Q => 
        \BIT_OS_SEL[1]\);
    
    \U_ELK8_CH/U_SLAVE_1ELK/RECD_SER_WORD[2]\ : DFN1C0
      port map(D => \U_ELK8_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[2]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_8[2]\);
    
    HIEFFPLA_INST_0_42625 : NOR2A
      port map(A => \U50_PATTERNS/REG_ADDR[7]\, B => 
        HIEFFPLA_NET_0_119509, Y => HIEFFPLA_NET_0_119497);
    
    \U_ELK8_CH/U_SLAVE_1ELK/Q[8]\ : DFN1C0
      port map(D => \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/Q[8]_net_1\);
    
    HIEFFPLA_INST_0_60980 : MX2
      port map(A => HIEFFPLA_NET_0_117167, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_18[1]\, S => 
        HIEFFPLA_NET_0_117134, Y => HIEFFPLA_NET_0_116189);
    
    \U50_PATTERNS/ELINK_ADDRA_14[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120048, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_5, Q => 
        \U50_PATTERNS/ELINK_ADDRA_14[7]\);
    
    \U200A_TFC/LOC_STRT_ADDR[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120282, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_4, Q => \U200A_TFC/LOC_STRT_ADDR[0]\);
    
    HIEFFPLA_INST_0_42033 : AND2
      port map(A => \U50_PATTERNS/ELK_N_ACTIVE_net_1\, B => 
        HIEFFPLA_NET_0_119020, Y => HIEFFPLA_NET_0_119627);
    
    \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[3]\ : DFN1C0
      port map(D => 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[3]_net_1\);
    
    \U50_PATTERNS/ELINK_DINA_18[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119798, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_21, Q => 
        \U50_PATTERNS/ELINK_DINA_18[1]\);
    
    HIEFFPLA_INST_0_63240 : NAND2B
      port map(A => \OP_MODE_c_0[1]\, B => \PATT_TFC_DAT[3]\, Y
         => \U_TFC_SERDAT_SOURCE/N_SERDAT[3]\);
    
    AFLSDF_INV_62 : INV
      port map(A => \U_DDR_ELK0/ELK0_IN_DDR_R\, Y => 
        \AFLSDF_INV_62\);
    
    \U200B_ELINKS/R_RWB/U1\ : DFN1P0
      port map(D => HIEFFPLA_NET_0_120151, CLK => CLK_40M_GL, PRE
         => P_MASTER_POR_B_c_12, Q => ELKS_RWB);
    
    HIEFFPLA_INST_0_43189 : AND2B
      port map(A => \U50_PATTERNS/REG_STATE[4]_net_1\, B => 
        \U50_PATTERNS/REG_STATE[5]_net_1\, Y => 
        HIEFFPLA_NET_0_119351);
    
    HIEFFPLA_INST_0_42682 : AND3A
      port map(A => HIEFFPLA_NET_0_118996, B => 
        HIEFFPLA_NET_0_119424, C => 
        \U50_PATTERNS/REG_STATE_0[1]_net_1\, Y => 
        HIEFFPLA_NET_0_119484);
    
    HIEFFPLA_INST_0_37039 : AOI1A
      port map(A => \TFC_STRT_ADDR[3]\, B => 
        HIEFFPLA_NET_0_120349, C => HIEFFPLA_NET_0_120361, Y => 
        HIEFFPLA_NET_0_120362);
    
    HIEFFPLA_INST_0_56662 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_0[3]\, B => 
        HIEFFPLA_NET_0_116797, S => HIEFFPLA_NET_0_117602, Y => 
        HIEFFPLA_NET_0_116821);
    
    HIEFFPLA_INST_0_41709 : MX2
      port map(A => HIEFFPLA_NET_0_119686, B => 
        \U50_PATTERNS/ELINK_RWA[14]\, S => 
        \U50_PATTERNS/SM_BANK_SEL_0[20]\, Y => 
        HIEFFPLA_NET_0_119706);
    
    \U_ELK19_CH/U_ELK1_CMD_TX/SER_OUT_RDEL\ : DFN1C0
      port map(D => \U_ELK19_CH/U_ELK1_CMD_TX/SER_OUT_RI_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_12, Q
         => \U_ELK19_CH/ELK_OUT_R\);
    
    \U50_PATTERNS/ELINK_BLKA[12]/U1\ : DFN1P0
      port map(D => HIEFFPLA_NET_0_119932, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_20, Q => 
        \U50_PATTERNS/ELINK_BLKA[12]\);
    
    HIEFFPLA_INST_0_43826 : MX2
      port map(A => HIEFFPLA_NET_0_119523, B => 
        \U50_PATTERNS/TFC_ADDRA[1]\, S => HIEFFPLA_NET_0_119294, 
        Y => HIEFFPLA_NET_0_119206);
    
    \U50_PATTERNS/ELINK_ADDRA_19[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120009, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_13, Q => 
        \U50_PATTERNS/ELINK_ADDRA_19[6]\);
    
    HIEFFPLA_INST_0_44006 : MX2
      port map(A => \U50_PATTERNS/TFC_STOP_ADDR[3]\, B => 
        \U50_PATTERNS/TFC_STOP_ADDR_T[3]\, S => 
        HIEFFPLA_NET_0_119472, Y => HIEFFPLA_NET_0_119185);
    
    \U_ELK3_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U1\ : IOBI_ID_OD_EB
      port map(DR => \U_ELK3_CH/ELK_OUT_R_i_0\, DF => 
        \U_ELK3_CH/ELK_OUT_F_i_0\, CLR => \GND\, E => 
        \AFLSDF_INV_38\, ICLK => CCC_160M_ADJ, OCLK => 
        CCC_160M_FXD, YIN => 
        \U_ELK3_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\, DOUT => 
        \U_ELK3_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, EOUT => 
        \U_ELK3_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET2\, YR => 
        \U_ELK3_CH/U_DDR_ELK1/ELK_IN_DDR_R\, YF => 
        \U_ELK3_CH/U_DDR_ELK1/ELK_IN_DDR_F\);
    
    HIEFFPLA_INST_0_58552 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_16[2]\, B => 
        HIEFFPLA_NET_0_116687, S => HIEFFPLA_NET_0_117215, Y => 
        HIEFFPLA_NET_0_116506);
    
    HIEFFPLA_INST_0_60738 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_15[3]\, B => 
        HIEFFPLA_NET_0_117186, S => HIEFFPLA_NET_0_117356, Y => 
        HIEFFPLA_NET_0_116227);
    
    \U_ELK11_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]\ : DFN1C0
      port map(D => \U_ELK11_CH/U_SLAVE_1ELK/Q[5]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]_net_1\);
    
    \U_ELK2_CH/ELK_IN_F\ : DFN1C0
      port map(D => \U_ELK2_CH/ELK_IN_DDR_F\, CLK => CCC_160M_ADJ, 
        CLR => DEV_RST_B_c, Q => \U_ELK2_CH/ELK_IN_F_net_1\);
    
    HIEFFPLA_INST_0_63128 : NOR2A
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[5]\, 
        B => HIEFFPLA_NET_0_115920, Y => HIEFFPLA_NET_0_115881);
    
    HIEFFPLA_INST_0_52160 : NAND2B
      port map(A => HIEFFPLA_NET_0_117624, B => 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM[3]_net_1\, Y => 
        HIEFFPLA_NET_0_117619);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_22[4]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116126, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_5, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_22[4]\);
    
    HIEFFPLA_INST_0_63185 : AX1C
      port map(A => HIEFFPLA_NET_0_117338, B => 
        HIEFFPLA_NET_0_117222, C => HIEFFPLA_NET_0_117226, Y => 
        HIEFFPLA_NET_0_115867);
    
    HIEFFPLA_INST_0_60941 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_17[2]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_18[2]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_4[0]\, Y => 
        HIEFFPLA_NET_0_116195);
    
    HIEFFPLA_INST_0_56171 : XA1C
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/MAX_CNT[2]\, 
        B => HIEFFPLA_NET_0_116944, C => HIEFFPLA_NET_0_117112, Y
         => HIEFFPLA_NET_0_116937);
    
    \U_EXEC_MASTER/MPOR_SALT_B_17\ : DFI1P0
      port map(D => HIEFFPLA_NET_0_117781, CLK => CLK_40M_GL, PRE
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_2\, QN => 
        MASTER_SALT_POR_B_i_0_i_17);
    
    HIEFFPLA_INST_0_42235 : AND3A
      port map(A => \U50_PATTERNS/RD_USB_ADBUS[3]\, B => 
        HIEFFPLA_NET_0_119589, C => 
        \U50_PATTERNS/RD_USB_ADBUS[2]\, Y => 
        HIEFFPLA_NET_0_119595);
    
    HIEFFPLA_INST_0_49837 : MX2
      port map(A => 
        \U_ELK4_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]_net_1\, B => 
        \U_ELK4_CH/ELK_TX_DAT[6]\, S => 
        \U_ELK4_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118064);
    
    HIEFFPLA_INST_0_48752 : MX2
      port map(A => HIEFFPLA_NET_0_118260, B => 
        HIEFFPLA_NET_0_118274, S => \BIT_OS_SEL_2[0]\, Y => 
        \U_ELK18_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[2]\);
    
    \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[8]\ : DFN1C0
      port map(D => 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\);
    
    HIEFFPLA_INST_0_46005 : AND3B
      port map(A => HIEFFPLA_NET_0_119426, B => 
        HIEFFPLA_NET_0_119379, C => \U50_PATTERNS/OP_MODE[5]\, Y
         => HIEFFPLA_NET_0_118789);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_7[4]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_115976, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_18, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_7[4]\);
    
    \U50_PATTERNS/ELINKS_STOP_ADDR[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120120, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_14, Q => 
        \U50_PATTERNS/ELINKS_STOP_ADDR[7]\);
    
    HIEFFPLA_INST_0_37077 : XO1
      port map(A => HIEFFPLA_NET_0_120262, B => \TFC_ADDRB[1]\, C
         => \U200A_TFC/GP_PG_SM[10]_net_1\, Y => 
        HIEFFPLA_NET_0_120352);
    
    HIEFFPLA_INST_0_48688 : MX2
      port map(A => \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\, 
        B => \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\, S => 
        \BIT_OS_SEL_0[2]\, Y => HIEFFPLA_NET_0_118266);
    
    HIEFFPLA_INST_0_43300 : MX2
      port map(A => \U50_PATTERNS/SI_CNT[3]\, B => 
        HIEFFPLA_NET_0_119324, S => HIEFFPLA_NET_0_119439, Y => 
        HIEFFPLA_NET_0_119331);
    
    HIEFFPLA_INST_0_38058 : AO1A
      port map(A => \ELKS_STRT_ADDR[4]\, B => 
        HIEFFPLA_NET_0_120219, C => HIEFFPLA_NET_0_120166, Y => 
        HIEFFPLA_NET_0_120163);
    
    HIEFFPLA_INST_0_41530 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_8[0]\, B => 
        HIEFFPLA_NET_0_119578, S => HIEFFPLA_NET_0_119291, Y => 
        HIEFFPLA_NET_0_119727);
    
    HIEFFPLA_INST_0_40234 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_0[0]\, B => 
        HIEFFPLA_NET_0_119578, S => HIEFFPLA_NET_0_119272, Y => 
        HIEFFPLA_NET_0_119871);
    
    HIEFFPLA_INST_0_45578 : AO1A
      port map(A => HIEFFPLA_NET_0_119622, B => 
        \U50_PATTERNS/TFC_STOP_ADDR[2]\, C => 
        HIEFFPLA_NET_0_118779, Y => HIEFFPLA_NET_0_118887);
    
    \U_ELK5_CH/U_SLAVE_1ELK/Q[4]\ : DFN1C0
      port map(D => \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/Q[4]_net_1\);
    
    HIEFFPLA_INST_0_62248 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_31[3]\, B => 
        HIEFFPLA_NET_0_117186, S => HIEFFPLA_NET_0_117319, Y => 
        HIEFFPLA_NET_0_116017);
    
    \U50_PATTERNS/U4C_REGCROSS/SAMP_TWO[4]\ : DFN1C0
      port map(D => \U50_PATTERNS/U4C_REGCROSS/SAMP_ONE[4]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_22_0, Q => 
        \U50_PATTERNS/U4C_REGCROSS/SAMP_TWO[4]_net_1\);
    
    HIEFFPLA_INST_0_51579 : AX1C
      port map(A => HIEFFPLA_NET_0_117746, B => 
        HIEFFPLA_NET_0_117753, C => HIEFFPLA_NET_0_117734, Y => 
        HIEFFPLA_NET_0_117740);
    
    HIEFFPLA_INST_0_51463 : MX2
      port map(A => HIEFFPLA_NET_0_117762, B => 
        \U_EXEC_MASTER/PRESCALE[0]\, S => HIEFFPLA_NET_0_117787, 
        Y => HIEFFPLA_NET_0_117768);
    
    \U200B_ELINKS/GP_PG_SM[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120214, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_29, Q => 
        \U200B_ELINKS/GP_PG_SM[2]_net_1\);
    
    HIEFFPLA_INST_0_45342 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_4[2]\, C => 
        \U50_PATTERNS/SM_BANK_SEL[15]\, Y => 
        HIEFFPLA_NET_0_118935);
    
    HIEFFPLA_INST_0_57122 : AO1A
      port map(A => HIEFFPLA_NET_0_116740, B => 
        HIEFFPLA_NET_0_116774, C => HIEFFPLA_NET_0_116708, Y => 
        HIEFFPLA_NET_0_116735);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_9[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_115963, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_20, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_9[2]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/PHASE_ADJ[0]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[0]_net_1\, CLK
         => CLK_40M_GL, CLR => P_MASTER_POR_B_c, Q => 
        \U_MASTER_DES/PHASE_ADJ_160_L[0]\);
    
    HIEFFPLA_INST_0_42546 : NAND3
      port map(A => \U50_PATTERNS/REG_ADDR[2]\, B => 
        \U50_PATTERNS/REG_ADDR[1]\, C => 
        \U50_PATTERNS/REG_ADDR[0]\, Y => HIEFFPLA_NET_0_119514);
    
    \U_ELK0_SERDAT_SOURCE/SERDAT[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118659, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_10, Q => \ELK0_TX_DAT[1]\);
    
    HIEFFPLA_INST_0_45036 : AND3B
      port map(A => \U50_PATTERNS/REG_STATE[0]_net_1\, B => 
        \U50_PATTERNS/USB_TXE_B\, C => HIEFFPLA_NET_0_119424, Y
         => HIEFFPLA_NET_0_118993);
    
    \U_ELK4_CH/U_ELK1_SERDAT_SOURCE/SERDAT[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118055, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_16, Q => 
        \U_ELK4_CH/ELK_TX_DAT[3]\);
    
    HIEFFPLA_INST_0_52087 : MX2C
      port map(A => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[72]_net_1\, B => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[73]_net_1\, S => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[0]\, Y => 
        HIEFFPLA_NET_0_117639);
    
    HIEFFPLA_INST_0_39263 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_19[5]\, B => 
        HIEFFPLA_NET_0_119518, S => HIEFFPLA_NET_0_119293, Y => 
        HIEFFPLA_NET_0_120010);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_1[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116785, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_4, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_1[3]\);
    
    HIEFFPLA_INST_0_48118 : NAND2B
      port map(A => \OP_MODE_c_2[1]\, B => \PATT_ELK_DAT_16[1]\, 
        Y => HIEFFPLA_NET_0_118372);
    
    \U50_PATTERNS/SM_BANK_SEL[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119303, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_7, Q => 
        \U50_PATTERNS/SM_BANK_SEL[7]\);
    
    HIEFFPLA_INST_0_59447 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_27[1]\, B => 
        HIEFFPLA_NET_0_116677, S => HIEFFPLA_NET_0_117162, Y => 
        HIEFFPLA_NET_0_116393);
    
    HIEFFPLA_INST_0_45959 : NAND3C
      port map(A => HIEFFPLA_NET_0_118947, B => 
        HIEFFPLA_NET_0_118956, C => HIEFFPLA_NET_0_118701, Y => 
        HIEFFPLA_NET_0_118801);
    
    HIEFFPLA_INST_0_45024 : AND3A
      port map(A => \U50_PATTERNS/USB_TXE_B\, B => 
        HIEFFPLA_NET_0_119267, C => 
        \U50_PATTERNS/REG_STATE_0[5]_net_1\, Y => 
        HIEFFPLA_NET_0_118997);
    
    HIEFFPLA_INST_0_54173 : MX2
      port map(A => HIEFFPLA_NET_0_116134, B => 
        HIEFFPLA_NET_0_116242, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_1[3]_net_1\, Y
         => HIEFFPLA_NET_0_117299);
    
    \U_MASTER_DES/U13C_MASTER_DESER/ARB_WRD_40M_FIXED[2]\ : 
        DFN1C0
      port map(D => \U_MASTER_DES/U13C_MASTER_DESER/Q[2]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_26, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_WRD_40M_FIXED[2]_net_1\);
    
    HIEFFPLA_INST_0_40612 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_14[2]\, B => 
        HIEFFPLA_NET_0_119575, S => HIEFFPLA_NET_0_119249, Y => 
        HIEFFPLA_NET_0_119829);
    
    HIEFFPLA_INST_0_57333 : AOI1A
      port map(A => HIEFFPLA_NET_0_116712, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_3[6]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_3[7]\, Y => 
        HIEFFPLA_NET_0_116697);
    
    HIEFFPLA_INST_0_53578 : MX2
      port map(A => HIEFFPLA_NET_0_116317, B => 
        HIEFFPLA_NET_0_116371, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[3]_net_1\, Y
         => HIEFFPLA_NET_0_117387);
    
    HIEFFPLA_INST_0_49041 : MX2
      port map(A => HIEFFPLA_NET_0_118222, B => 
        HIEFFPLA_NET_0_118205, S => \BIT_OS_SEL_2[0]\, Y => 
        \U_ELK19_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[7]\);
    
    \U_ELK19_CH/ELK_IN_R\ : DFN1C0
      port map(D => \U_ELK19_CH/ELK_IN_DDR_R\, CLK => 
        CCC_160M_ADJ, CLR => DEV_RST_B_c, Q => 
        \U_ELK19_CH/ELK_IN_R_net_1\);
    
    HIEFFPLA_INST_0_111269 : AOI1D
      port map(A => HIEFFPLA_NET_0_116740, B => 
        HIEFFPLA_NET_0_116345, C => HIEFFPLA_NET_0_117328, Y => 
        HIEFFPLA_NET_0_115845);
    
    HIEFFPLA_INST_0_54165 : MX2
      port map(A => HIEFFPLA_NET_0_116196, B => 
        HIEFFPLA_NET_0_116081, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_1[3]_net_1\, Y
         => HIEFFPLA_NET_0_117300);
    
    HIEFFPLA_INST_0_111642 : OA1C
      port map(A => HIEFFPLA_NET_0_115837, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/TUNE_CLKPHASE[0]\, C => 
        HIEFFPLA_NET_0_117077, Y => HIEFFPLA_NET_0_115940);
    
    HIEFFPLA_INST_0_111346 : MX2A
      port map(A => HIEFFPLA_NET_0_115841, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_23[3]\, S => 
        HIEFFPLA_NET_0_117214, Y => HIEFFPLA_NET_0_116435);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_12[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116252, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_21, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_12[3]\);
    
    \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[9]\ : DFN1C0
      port map(D => 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\);
    
    \U_ELK2_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]\ : DFN1C0
      port map(D => \U_ELK2_CH/U_SLAVE_1ELK/Q[7]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]_net_1\);
    
    HIEFFPLA_INST_0_42555 : AND3B
      port map(A => \U50_PATTERNS/REG_ADDR[2]\, B => 
        \U50_PATTERNS/REG_ADDR[4]\, C => 
        \U50_PATTERNS/REG_ADDR[8]\, Y => HIEFFPLA_NET_0_119512);
    
    \U_MASTER_DES/U13C_MASTER_DESER/ARB_WRD_40M_FIXED[12]\ : 
        DFN1C0
      port map(D => \U_MASTER_DES/U13C_MASTER_DESER/Q[12]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_28, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_WRD_40M_FIXED[12]_net_1\);
    
    \U50_PATTERNS/ELINK_DINA_2[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119769, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_9, Q => 
        \U50_PATTERNS/ELINK_DINA_2[6]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_14[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116526, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_13, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_14[2]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_23[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116440, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_17_0, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_23[2]\);
    
    \U50_PATTERNS/OP_MODE[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119614, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_15, Q => \U50_PATTERNS/OP_MODE[3]\);
    
    HIEFFPLA_INST_0_43324 : XA1B
      port map(A => \U50_PATTERNS/SI_CNT[1]\, B => 
        \U50_PATTERNS/SI_CNT[0]\, C => HIEFFPLA_NET_0_119329, Y
         => HIEFFPLA_NET_0_119326);
    
    HIEFFPLA_INST_0_48037 : MX2
      port map(A => HIEFFPLA_NET_0_118400, B => 
        HIEFFPLA_NET_0_118396, S => \BIT_OS_SEL_3[0]\, Y => 
        \U_ELK15_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[6]\);
    
    HIEFFPLA_INST_0_43094 : MX2B
      port map(A => HIEFFPLA_NET_0_119441, B => 
        \U50_PATTERNS/REG_STATE[1]_net_1\, S => 
        \U50_PATTERNS/REG_STATE[0]_net_1\, Y => 
        HIEFFPLA_NET_0_119381);
    
    \U_MASTER_DES/U13C_MASTER_DESER/MAX_CNT[8]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_116946, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_16, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/MAX_CNT[8]\);
    
    HIEFFPLA_INST_0_43178 : AND3B
      port map(A => \U50_PATTERNS/REG_STATE_0[4]_net_1\, B => 
        \U50_PATTERNS/REG_STATE[0]_net_1\, C => 
        HIEFFPLA_NET_0_119429, Y => HIEFFPLA_NET_0_119354);
    
    \U50_PATTERNS/ELINK_ADDRA_15[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120042, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_6, Q => 
        \U50_PATTERNS/ELINK_ADDRA_15[5]\);
    
    \U50_PATTERNS/ELINK_ADDRA_12[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120064, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_3, Q => 
        \U50_PATTERNS/ELINK_ADDRA_12[7]\);
    
    HIEFFPLA_INST_0_111419 : OR3B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[2]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[1]_net_1\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[7]_net_1\, Y => 
        HIEFFPLA_NET_0_115838);
    
    \U_ELK7_CH/U_ELK1_CMD_TX/SER_OUT_RDEL\ : DFN1C0
      port map(D => \U_ELK7_CH/U_ELK1_CMD_TX/SER_OUT_RI_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_8, Q
         => \U_ELK7_CH/ELK_OUT_R\);
    
    HIEFFPLA_INST_0_39362 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_2[0]\, B => 
        HIEFFPLA_NET_0_119524, S => HIEFFPLA_NET_0_119278, Y => 
        HIEFFPLA_NET_0_119999);
    
    \U_ELK7_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U0\ : IOPADP_BI
      port map(N2PIN => 
        \U_ELK7_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2_N2P\, D => 
        \U_ELK7_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, E => 
        \U_ELK7_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET2\, PAD => 
        ELK7_DAT_P, Y => 
        \U_ELK7_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\);
    
    HIEFFPLA_INST_0_40954 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_19[0]\, B => 
        HIEFFPLA_NET_0_119578, S => HIEFFPLA_NET_0_119293, Y => 
        HIEFFPLA_NET_0_119791);
    
    HIEFFPLA_INST_0_45805 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/SM_BANK_SEL[19]\, C => 
        \U50_PATTERNS/ELINK_DOUTA_0[0]\, Y => 
        HIEFFPLA_NET_0_118837);
    
    \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[12]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_115931, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_21, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[12]\);
    
    HIEFFPLA_INST_0_56370 : AO1
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[6]_net_1\, B => 
        HIEFFPLA_NET_0_117431, C => HIEFFPLA_NET_0_116860, Y => 
        HIEFFPLA_NET_0_116884);
    
    HIEFFPLA_INST_0_46013 : AND2A
      port map(A => HIEFFPLA_NET_0_119622, B => 
        \U50_PATTERNS/TFC_STOP_ADDR[0]\, Y => 
        HIEFFPLA_NET_0_118787);
    
    HIEFFPLA_INST_0_47341 : MX2
      port map(A => 
        \U_ELK13_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]_net_1\, B => 
        \U_ELK13_CH/ELK_TX_DAT[4]\, S => 
        \U_ELK13_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118515);
    
    HIEFFPLA_INST_0_61295 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_19[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_20[1]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_4[0]\, Y => 
        HIEFFPLA_NET_0_116146);
    
    HIEFFPLA_INST_0_49120 : NAND2B
      port map(A => \OP_MODE_c_5[1]\, B => \PATT_ELK_DAT_1[7]\, Y
         => HIEFFPLA_NET_0_118186);
    
    HIEFFPLA_INST_0_58066 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_0[3]\, B => 
        HIEFFPLA_NET_0_116563, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_1[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116569);
    
    HIEFFPLA_INST_0_50535 : MX2
      port map(A => HIEFFPLA_NET_0_117958, B => 
        HIEFFPLA_NET_0_117935, S => \BIT_OS_SEL[0]\, Y => 
        \U_ELK6_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[7]\);
    
    \U50_PATTERNS/TFC_STOP_ADDR_T[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119178, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_15, Q => 
        \U50_PATTERNS/TFC_STOP_ADDR_T[2]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117043, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_17, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[2]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/Q[0]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[0]_net_1\, CLK => 
        CCC_160M_FXD, CLR => P_MASTER_POR_B_c_34, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/Q[0]_net_1\);
    
    \U_ELK11_CH/U_SLAVE_1ELK/Q[3]\ : DFN1C0
      port map(D => \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/Q[3]_net_1\);
    
    \U_ELK3_CH/U_SLAVE_1ELK/Q[13]\ : DFN1C0
      port map(D => \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[13]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/Q[13]_net_1\);
    
    \U_ELK15_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U3\ : IOBI_ID_OD_EB
      port map(DR => \U_ELK15_CH/ELK_OUT_R\, DF => 
        \U_ELK15_CH/ELK_OUT_F\, CLR => \GND\, E => 
        \AFLSDF_INV_25\, ICLK => CCC_160M_ADJ, OCLK => 
        CCC_160M_FXD, YIN => 
        \U_ELK15_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\, DOUT => 
        OPEN, EOUT => 
        \U_ELK15_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET3\, YR => OPEN, 
        YF => OPEN);
    
    HIEFFPLA_INST_0_60862 : AND2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[4]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_16[4]\, Y => 
        HIEFFPLA_NET_0_116206);
    
    \U_ELK10_CH/U_SLAVE_1ELK/RECD_SER_WORD[7]\ : DFN1C0
      port map(D => \U_ELK10_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[7]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_10[7]\);
    
    HIEFFPLA_INST_0_43341 : MX2
      port map(A => \U50_PATTERNS/SM_BANK_SEL[0]\, B => 
        HIEFFPLA_NET_0_119228, S => HIEFFPLA_NET_0_118691, Y => 
        HIEFFPLA_NET_0_119322);
    
    HIEFFPLA_INST_0_42420 : AND2
      port map(A => HIEFFPLA_NET_0_119473, B => 
        \U50_PATTERNS/RD_XFER_TYPE[0]_net_1\, Y => 
        HIEFFPLA_NET_0_119541);
    
    \U_ELK7_CH/U_SLAVE_1ELK/Q[7]\ : DFN1C0
      port map(D => \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/Q[7]_net_1\);
    
    \U_ELK3_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]\ : DFN1C0
      port map(D => \U_ELK3_CH/U_SLAVE_1ELK/Q[13]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]_net_1\);
    
    \U_ELK12_CH/U_SLAVE_1ELK/Q[4]\ : DFN1C0
      port map(D => \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/Q[4]_net_1\);
    
    \U50_PATTERNS/ELINK_ADDRA_10[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120082, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_22, Q => 
        \U50_PATTERNS/ELINK_ADDRA_10[5]\);
    
    HIEFFPLA_INST_0_52830 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_15[0]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_16[0]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_2[0]\, Y => 
        HIEFFPLA_NET_0_117504);
    
    HIEFFPLA_INST_0_47981 : MX2
      port map(A => HIEFFPLA_NET_0_118408, B => 
        HIEFFPLA_NET_0_118405, S => \BIT_OS_SEL_2[1]\, Y => 
        HIEFFPLA_NET_0_118395);
    
    HIEFFPLA_INST_0_56152 : NAND3
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/MAX_CNT[0]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/MAX_CNT[1]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/MAX_CNT[2]\, Y => 
        HIEFFPLA_NET_0_116942);
    
    HIEFFPLA_INST_0_39155 : MX2
      port map(A => HIEFFPLA_NET_0_119523, B => 
        \U50_PATTERNS/ELINK_ADDRA_18[1]\, S => 
        HIEFFPLA_NET_0_119264, Y => HIEFFPLA_NET_0_120022);
    
    HIEFFPLA_INST_0_54934 : XA1B
      port map(A => HIEFFPLA_NET_0_117222, B => 
        HIEFFPLA_NET_0_117338, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_0[8]_net_1\, Y => 
        HIEFFPLA_NET_0_117167);
    
    HIEFFPLA_INST_0_39839 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_8[5]\, B => 
        HIEFFPLA_NET_0_119518, S => HIEFFPLA_NET_0_119291, Y => 
        HIEFFPLA_NET_0_119946);
    
    AFLSDF_INV_9 : INV
      port map(A => P_USB_MASTER_EN_c_22_0, Y => \AFLSDF_INV_9\);
    
    \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[0]\ : DFN1C0
      port map(D => 
        \U_ELK10_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\);
    
    HIEFFPLA_INST_0_44962 : AO1A
      port map(A => HIEFFPLA_NET_0_119379, B => 
        HIEFFPLA_NET_0_118995, C => HIEFFPLA_NET_0_119001, Y => 
        HIEFFPLA_NET_0_119011);
    
    \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[7]\ : DFN1C0
      port map(D => \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\);
    
    HIEFFPLA_INST_0_46560 : MX2
      port map(A => \U_ELK0_CMD_TX/SER_CMD_WORD_R[0]_net_1\, B
         => \ELK0_TX_DAT[3]\, S => 
        \U_ELK0_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118664);
    
    \U_MASTER_DES/U13C_MASTER_DESER/MAX_CNT[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_116954, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_15, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/MAX_CNT[0]\);
    
    HIEFFPLA_INST_0_62667 : MX2
      port map(A => HIEFFPLA_NET_0_117100, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_9[4]\, S => 
        HIEFFPLA_NET_0_117183, Y => HIEFFPLA_NET_0_115961);
    
    HIEFFPLA_INST_0_57630 : NAND3
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_5[3]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_5[2]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_5[1]\, Y => 
        HIEFFPLA_NET_0_116648);
    
    HIEFFPLA_INST_0_61670 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_25[1]\, B => 
        HIEFFPLA_NET_0_117167, S => HIEFFPLA_NET_0_117117, Y => 
        HIEFFPLA_NET_0_116094);
    
    HIEFFPLA_INST_0_61544 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_7[4]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_23[4]\, S
         => \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[4]_net_1\, 
        Y => HIEFFPLA_NET_0_116112);
    
    HIEFFPLA_INST_0_59346 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_26[3]\, B => 
        HIEFFPLA_NET_0_116399, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_2[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116403);
    
    HIEFFPLA_INST_0_47120 : AND2
      port map(A => CLK_40M_GL, B => 
        \U_ELK12_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0_net_1\, Y => 
        HIEFFPLA_NET_0_118554);
    
    HIEFFPLA_INST_0_46299 : NAND3B
      port map(A => HIEFFPLA_NET_0_118887, B => 
        HIEFFPLA_NET_0_118869, C => HIEFFPLA_NET_0_119427, Y => 
        HIEFFPLA_NET_0_118722);
    
    HIEFFPLA_INST_0_61622 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_24[4]\, B => 
        HIEFFPLA_NET_0_117166, S => HIEFFPLA_NET_0_117074, Y => 
        HIEFFPLA_NET_0_116101);
    
    HIEFFPLA_INST_0_49610 : AND2
      port map(A => CLK_40M_GL, B => 
        \U_ELK3_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0_net_1\, Y => 
        HIEFFPLA_NET_0_118104);
    
    HIEFFPLA_INST_0_161267 : DFN1C0
      port map(D => \U_ELK1_CH/ELK_TX_DAT[1]\, CLK => 
        CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_4, Q => 
        HIEFFPLA_NET_0_161288);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_28[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116386, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_2, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_28[0]\);
    
    HIEFFPLA_INST_0_44480 : MX2
      port map(A => \ELKS_STRT_ADDR[4]\, B => 
        \U50_PATTERNS/U4C_REGCROSS/SAMP_TWO[4]_net_1\, S => 
        HIEFFPLA_NET_0_119114, Y => HIEFFPLA_NET_0_119108);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_27[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116394, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_1, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_27[0]\);
    
    \U_ELK1_CH/U_SLAVE_1ELK/Q[8]\ : DFN1C0
      port map(D => \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/Q[8]_net_1\);
    
    \U50_PATTERNS/CHKSUM[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120141, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_3, Q => \U50_PATTERNS/CHKSUM[2]\);
    
    \U_ELK10_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL\ : DFN1C0
      port map(D => \U_ELK10_CH/ELK_IN_R_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL_net_1\);
    
    HIEFFPLA_INST_0_47563 : MX2
      port map(A => HIEFFPLA_NET_0_118489, B => 
        HIEFFPLA_NET_0_118473, S => \BIT_OS_SEL_5[1]\, Y => 
        HIEFFPLA_NET_0_118475);
    
    \U_ELK8_CH/U_SLAVE_1ELK/RECD_SER_WORD[7]\ : DFN1C0
      port map(D => \U_ELK8_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[7]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_8[7]\);
    
    HIEFFPLA_INST_0_61964 : MX2
      port map(A => HIEFFPLA_NET_0_117131, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_28[2]\, S => 
        HIEFFPLA_NET_0_117146, Y => HIEFFPLA_NET_0_116053);
    
    HIEFFPLA_INST_0_53475 : MX2
      port map(A => HIEFFPLA_NET_0_117421, B => 
        HIEFFPLA_NET_0_117345, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[1]_net_1\, Y
         => HIEFFPLA_NET_0_117402);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_28[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116385, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_2, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_28[1]\);
    
    HIEFFPLA_INST_0_111822 : MX2B
      port map(A => 
        \U_EXEC_MASTER/USB_MASTER_EN/CNT_EN_60M2S_net_1\, B => 
        HIEFFPLA_NET_0_115828, S => HIEFFPLA_NET_0_117753, Y => 
        HIEFFPLA_NET_0_117738);
    
    HIEFFPLA_INST_0_47033 : MX2
      port map(A => HIEFFPLA_NET_0_118588, B => 
        HIEFFPLA_NET_0_118583, S => \BIT_OS_SEL[0]\, Y => 
        \U_ELK11_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[5]\);
    
    HIEFFPLA_INST_0_37405 : MX2
      port map(A => \U200A_TFC/LOC_STOP_ADDR[0]\, B => 
        \TFC_STOP_ADDR[0]\, S => \U200A_TFC/GP_PG_SM_0[10]_net_1\, 
        Y => HIEFFPLA_NET_0_120290);
    
    \U_EXEC_MASTER/MPOR_B\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117787, CLK => CLK_40M_GL, CLR
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i\, Q => 
        P_MASTER_POR_B_c);
    
    HIEFFPLA_INST_0_54865 : XA1B
      port map(A => HIEFFPLA_NET_0_117225, B => 
        HIEFFPLA_NET_0_115866, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_0[8]_net_1\, Y => 
        HIEFFPLA_NET_0_117186);
    
    HIEFFPLA_INST_0_58574 : AOI1D
      port map(A => HIEFFPLA_NET_0_116675, B => 
        HIEFFPLA_NET_0_116589, C => HIEFFPLA_NET_0_117215, Y => 
        HIEFFPLA_NET_0_116503);
    
    HIEFFPLA_INST_0_45350 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_12[4]\, C => 
        \U50_PATTERNS/SM_BANK_SEL[7]\, Y => HIEFFPLA_NET_0_118933);
    
    \U_ELK8_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]\ : DFN1C0
      port map(D => \U_ELK8_CH/U_SLAVE_1ELK/Q[2]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]_net_1\);
    
    HIEFFPLA_INST_0_55941 : MX2
      port map(A => HIEFFPLA_NET_0_117025, B => 
        HIEFFPLA_NET_0_116958, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[4]\, Y => 
        HIEFFPLA_NET_0_116970);
    
    HIEFFPLA_INST_0_48760 : MX2
      port map(A => HIEFFPLA_NET_0_118274, B => 
        HIEFFPLA_NET_0_118269, S => \BIT_OS_SEL_2[0]\, Y => 
        \U_ELK18_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[3]\);
    
    HIEFFPLA_INST_0_48519 : MX2
      port map(A => HIEFFPLA_NET_0_118315, B => 
        HIEFFPLA_NET_0_118313, S => \BIT_OS_SEL_3[0]\, Y => 
        \U_ELK17_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[4]\);
    
    \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[11]\ : DFN1C0
      port map(D => \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\);
    
    HIEFFPLA_INST_0_45898 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/SM_BANK_SEL[13]\, C => 
        \U50_PATTERNS/ELINK_DOUTA_6[3]\, Y => 
        HIEFFPLA_NET_0_118817);
    
    \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[8]\ : DFN1C0
      port map(D => \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\);
    
    HIEFFPLA_INST_0_40084 : AOI1D
      port map(A => HIEFFPLA_NET_0_119389, B => 
        HIEFFPLA_NET_0_119464, C => \U50_PATTERNS/SM_BANK_SEL[9]\, 
        Y => HIEFFPLA_NET_0_119912);
    
    \U_ELK17_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118330, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_14, Q => 
        \U_ELK17_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]_net_1\);
    
    HIEFFPLA_INST_0_63123 : AX1A
      port map(A => HIEFFPLA_NET_0_115905, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[3]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[4]\, Y => 
        HIEFFPLA_NET_0_115882);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_2[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116753, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_5, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_2[2]\);
    
    HIEFFPLA_INST_0_62693 : XNOR3
      port map(A => HIEFFPLA_NET_0_115958, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_CLKPHASE[2]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_SEQCNT[3]\, Y => 
        HIEFFPLA_NET_0_115956);
    
    \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[3]\ : DFN1C0
      port map(D => 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[3]_net_1\);
    
    \U_ELK15_CH/U_ELK1_CMD_TX/SER_OUT_FI\ : DFN1C0
      port map(D => 
        \U_ELK15_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_1, Q => 
        \U_ELK15_CH/U_ELK1_CMD_TX/SER_OUT_FI_net_1\);
    
    \U50_PATTERNS/TFC_STRT_ADDR[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119169, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_13, Q => 
        \U50_PATTERNS/TFC_STRT_ADDR[3]\);
    
    HIEFFPLA_INST_0_41993 : AO1
      port map(A => HIEFFPLA_NET_0_119584, B => 
        HIEFFPLA_NET_0_119630, C => HIEFFPLA_NET_0_119417, Y => 
        HIEFFPLA_NET_0_119636);
    
    \P_TFC_SYNC_DET_pad/U0/U1\ : IOTRI_OB_EB
      port map(D => P_TFC_SYNC_DET_c, E => \VCC\, DOUT => 
        \P_TFC_SYNC_DET_pad/U0/NET1\, EOUT => 
        \P_TFC_SYNC_DET_pad/U0/NET2\);
    
    \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[1]\ : DFN1C0
      port map(D => 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[1]_net_1\);
    
    HIEFFPLA_INST_0_63055 : AND2B
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[9]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[10]\, Y => 
        HIEFFPLA_NET_0_115901);
    
    HIEFFPLA_INST_0_52054 : MX2C
      port map(A => \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[46]\, B
         => \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[47]\, S => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[0]\, Y => 
        HIEFFPLA_NET_0_117645);
    
    HIEFFPLA_INST_0_43368 : MX2
      port map(A => \U50_PATTERNS/SM_BANK_SEL[12]\, B => 
        HIEFFPLA_NET_0_119225, S => HIEFFPLA_NET_0_118691, Y => 
        HIEFFPLA_NET_0_119319);
    
    \U_EXEC_MASTER/SYNC_BRD_RST_BI_2\ : DFI1P0
      port map(D => \U_EXEC_MASTER/DEV_RST_1B_i\, CLK => 
        CCC_160M_FXD, PRE => DEV_RST_B_c, QN => 
        \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_2\);
    
    \U50_PATTERNS/ELINK_ADDRA_1[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120003, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_20, Q => 
        \U50_PATTERNS/ELINK_ADDRA_1[4]\);
    
    \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_S\ : DFN1C0
      port map(D => 
        \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_40M_net_1\, CLK => 
        CLK60MHZ, CLR => P_MASTER_POR_B_c_34_0, Q => 
        \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_S_net_1\);
    
    \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[11]\ : DFN1C0
      port map(D => \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\);
    
    HIEFFPLA_INST_0_43579 : NAND2B
      port map(A => \U50_PATTERNS/SM_BANK_SEL[5]\, B => 
        HIEFFPLA_NET_0_119259, Y => HIEFFPLA_NET_0_119282);
    
    \U50_PATTERNS/U4D_REGCROSS/LOCAL_REG_VAL[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119091, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_3, Q => \ELKS_STOP_ADDR[0]\);
    
    \U_ELK9_CH/U_ELK1_CMD_TX/SER_OUT_FDEL\ : DFN1C0
      port map(D => \U_ELK9_CH/U_ELK1_CMD_TX/SER_OUT_FI_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_16, Q
         => \U_ELK9_CH/ELK_OUT_F\);
    
    \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[13]\ : DFN1C0
      port map(D => 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[13]_net_1\);
    
    \U_ELK17_CH/U_ELK1_SERDAT_SOURCE/SERDAT[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118326, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_11, Q => 
        \U_ELK17_CH/ELK_TX_DAT[2]\);
    
    HIEFFPLA_INST_0_46622 : AND2
      port map(A => CLK_40M_GL, B => 
        \U_ELK10_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0_net_1\, Y => 
        HIEFFPLA_NET_0_118644);
    
    \U_MASTER_DES/U13C_MASTER_DESER/Q[5]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[5]_net_1\, CLK => 
        CCC_160M_FXD, CLR => P_MASTER_POR_B_c_34, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/Q[5]_net_1\);
    
    \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[3]\ : DFN1C0
      port map(D => 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[3]_net_1\);
    
    \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[0]\ : DFN1C0
      port map(D => 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[0]_net_1\);
    
    \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[5]\ : DFN1C0
      port map(D => 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\);
    
    \U50_PATTERNS/ELINK_DINA_16[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119813, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_18, Q => 
        \U50_PATTERNS/ELINK_DINA_16[2]\);
    
    HIEFFPLA_INST_0_50120 : MX2
      port map(A => HIEFFPLA_NET_0_118001, B => 
        HIEFFPLA_NET_0_117999, S => \BIT_OS_SEL_6[1]\, Y => 
        HIEFFPLA_NET_0_118005);
    
    \U200A_TFC/ADDR_POINTER[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120362, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_30, Q => \TFC_ADDRB[3]\);
    
    \U_ELK2_CH/U_ELK1_SERDAT_SOURCE/SERDAT[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118145, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_13, Q => 
        \U_ELK2_CH/ELK_TX_DAT[3]\);
    
    HIEFFPLA_INST_0_53424 : NAND3C
      port map(A => HIEFFPLA_NET_0_116810, B => 
        HIEFFPLA_NET_0_117340, C => HIEFFPLA_NET_0_117406, Y => 
        HIEFFPLA_NET_0_117410);
    
    HIEFFPLA_INST_0_46165 : AO1
      port map(A => HIEFFPLA_NET_0_119254, B => 
        \U50_PATTERNS/ELINK_DOUTA_6[2]\, C => 
        HIEFFPLA_NET_0_118927, Y => HIEFFPLA_NET_0_118752);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_18[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116190, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_8, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_18[0]\);
    
    HIEFFPLA_INST_0_50503 : MX2
      port map(A => HIEFFPLA_NET_0_117956, B => 
        HIEFFPLA_NET_0_117951, S => \BIT_OS_SEL[0]\, Y => 
        \U_ELK6_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[3]\);
    
    HIEFFPLA_INST_0_46104 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/SM_BANK_SEL[16]\, C => 
        \U50_PATTERNS/ELINK_DOUTA_3[0]\, Y => 
        HIEFFPLA_NET_0_118765);
    
    HIEFFPLA_INST_0_51110 : AND2A
      port map(A => \OP_MODE_c_3[1]\, B => \PATT_ELK_DAT_9[5]\, Y
         => HIEFFPLA_NET_0_117828);
    
    \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[12]\ : DFN1C0
      port map(D => \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\);
    
    \U_ELK3_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]\ : DFN1C0
      port map(D => \U_ELK3_CH/U_SLAVE_1ELK/Q[3]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]_net_1\);
    
    HIEFFPLA_INST_0_46150 : AO1
      port map(A => HIEFFPLA_NET_0_119290, B => 
        \U50_PATTERNS/ELINK_DOUTA_17[7]\, C => 
        HIEFFPLA_NET_0_118930, Y => HIEFFPLA_NET_0_118755);
    
    \U_MASTER_DES/U13C_MASTER_DESER/ARB_WRD_40M_FIXED[6]\ : 
        DFN1C0
      port map(D => \U_MASTER_DES/U13C_MASTER_DESER/Q[6]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_26, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_WRD_40M_FIXED[6]_net_1\);
    
    HIEFFPLA_INST_0_52122 : AND2
      port map(A => HIEFFPLA_NET_0_117661, B => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[5]\, Y => 
        HIEFFPLA_NET_0_117632);
    
    HIEFFPLA_INST_0_42733 : XO1
      port map(A => \U50_PATTERNS/REG_STATE[0]_net_1\, B => 
        \U50_PATTERNS/REG_STATE_0[2]_net_1\, C => 
        HIEFFPLA_NET_0_119436, Y => HIEFFPLA_NET_0_119473);
    
    \U50_PATTERNS/OP_MODE[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119611, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_15, Q => \U50_PATTERNS/OP_MODE[6]\);
    
    HIEFFPLA_INST_0_51562 : MX2B
      port map(A => 
        \U_EXEC_MASTER/USB_MASTER_EN/CNT_EN_60M2S_net_1\, B => 
        \U_EXEC_MASTER/USB_MASTER_EN/T_CNT60M[0]_net_1\, S => 
        HIEFFPLA_NET_0_117753, Y => HIEFFPLA_NET_0_117743);
    
    HIEFFPLA_INST_0_42639 : AND3A
      port map(A => \U50_PATTERNS/REG_STATE_0[5]_net_1\, B => 
        \U50_PATTERNS/REG_STATE_0[4]_net_1\, C => 
        \U50_PATTERNS/REG_STATE[0]_net_1\, Y => 
        HIEFFPLA_NET_0_119494);
    
    \U_EXEC_MASTER/MPOR_B_31\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117787, CLK => CLK_40M_GL, CLR
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_0\, Q => 
        P_MASTER_POR_B_c_31);
    
    HIEFFPLA_INST_0_60286 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_8[3]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_24[3]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_1[4]_net_1\, Y
         => HIEFFPLA_NET_0_116286);
    
    HIEFFPLA_INST_0_51429 : XA1A
      port map(A => HIEFFPLA_NET_0_117786, B => 
        \U_EXEC_MASTER/DEL_CNT[2]\, C => 
        \U_EXEC_MASTER/CCC_1_LOCK_STAT_1D_net_1\, Y => 
        HIEFFPLA_NET_0_117776);
    
    HIEFFPLA_INST_0_48373 : NAND2B
      port map(A => \OP_MODE_c_6[1]\, B => \PATT_ELK_DAT_17[7]\, 
        Y => HIEFFPLA_NET_0_118321);
    
    HIEFFPLA_INST_0_61886 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_11[0]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_27[0]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_2[4]_net_1\, Y
         => HIEFFPLA_NET_0_116065);
    
    HIEFFPLA_INST_0_46624 : NAND2B
      port map(A => \OP_MODE_c_3[1]\, B => \PATT_ELK_DAT_10[1]\, 
        Y => HIEFFPLA_NET_0_118642);
    
    HIEFFPLA_INST_0_37057 : AOI1A
      port map(A => \TFC_STRT_ADDR[6]\, B => 
        HIEFFPLA_NET_0_120349, C => HIEFFPLA_NET_0_120355, Y => 
        HIEFFPLA_NET_0_120356);
    
    HIEFFPLA_INST_0_55834 : MX2
      port map(A => HIEFFPLA_NET_0_116989, B => 
        HIEFFPLA_NET_0_117004, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[2]\, Y => 
        HIEFFPLA_NET_0_116984);
    
    HIEFFPLA_INST_0_43582 : AND2B
      port map(A => \U50_PATTERNS/SM_BANK_SEL_0[21]\, B => 
        \U50_PATTERNS/SM_BANK_SEL[8]\, Y => HIEFFPLA_NET_0_119280);
    
    \U50_PATTERNS/U4A_REGCROSS/SYNC_SM[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119146, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_27, Q => 
        \U50_PATTERNS/U4A_REGCROSS/SYNC_SM[0]_net_1\);
    
    \U_ELK7_CH/U_SLAVE_1ELK/RECD_SER_WORD[0]\ : DFN1C0
      port map(D => \U_ELK7_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[0]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_7[0]\);
    
    HIEFFPLA_INST_0_41638 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_9[4]\, B => 
        HIEFFPLA_NET_0_119570, S => HIEFFPLA_NET_0_119292, Y => 
        HIEFFPLA_NET_0_119715);
    
    HIEFFPLA_INST_0_37196 : AND3C
      port map(A => \U200A_TFC/GP_PG_SM[2]_net_1\, B => 
        \U200A_TFC/GP_PG_SM[3]_net_1\, C => 
        \U200A_TFC/GP_PG_SM[0]_net_1\, Y => HIEFFPLA_NET_0_120326);
    
    HIEFFPLA_INST_0_60989 : MX2
      port map(A => HIEFFPLA_NET_0_117181, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_18[2]\, S => 
        HIEFFPLA_NET_0_117134, Y => HIEFFPLA_NET_0_116188);
    
    HIEFFPLA_INST_0_58916 : MX2
      port map(A => HIEFFPLA_NET_0_116687, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_20[2]\, S => 
        HIEFFPLA_NET_0_117203, Y => HIEFFPLA_NET_0_116458);
    
    HIEFFPLA_INST_0_43264 : AND3
      port map(A => HIEFFPLA_NET_0_119354, B => 
        HIEFFPLA_NET_0_119561, C => HIEFFPLA_NET_0_119568, Y => 
        HIEFFPLA_NET_0_119335);
    
    HIEFFPLA_INST_0_56950 : XA1B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_1[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_1[0]\, C => 
        HIEFFPLA_NET_0_117085, Y => HIEFFPLA_NET_0_116767);
    
    HIEFFPLA_INST_0_55176 : NAND3C
      port map(A => HIEFFPLA_NET_0_117378, B => 
        HIEFFPLA_NET_0_116768, C => HIEFFPLA_NET_0_117350, Y => 
        HIEFFPLA_NET_0_117105);
    
    \U_ELK11_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]\ : DFN1C0
      port map(D => \U_ELK11_CH/U_SLAVE_1ELK/Q[0]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]_net_1\);
    
    HIEFFPLA_INST_0_38237 : AND2A
      port map(A => HIEFFPLA_NET_0_119452, B => 
        \U50_PATTERNS/RD_USB_ADBUS[7]\, Y => 
        HIEFFPLA_NET_0_120128);
    
    HIEFFPLA_INST_0_39830 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_8[4]\, B => 
        HIEFFPLA_NET_0_119519, S => HIEFFPLA_NET_0_119291, Y => 
        HIEFFPLA_NET_0_119947);
    
    \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[8]\ : DFN1C0
      port map(D => \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\);
    
    HIEFFPLA_INST_0_48680 : MX2
      port map(A => HIEFFPLA_NET_0_118268, B => 
        HIEFFPLA_NET_0_118265, S => \BIT_OS_SEL_1[1]\, Y => 
        HIEFFPLA_NET_0_118267);
    
    HIEFFPLA_INST_0_48973 : MX2
      port map(A => \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\, 
        B => \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[13]_net_1\, S => 
        \BIT_OS_SEL_0[2]\, Y => HIEFFPLA_NET_0_118216);
    
    \U_ELK13_CH/ELK_IN_F\ : DFN1C0
      port map(D => \U_ELK13_CH/ELK_IN_DDR_F\, CLK => 
        CCC_160M_ADJ, CLR => DEV_RST_B_c, Q => 
        \U_ELK13_CH/ELK_IN_F_net_1\);
    
    HIEFFPLA_INST_0_61982 : MX2
      port map(A => HIEFFPLA_NET_0_117100, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_28[4]\, S => 
        HIEFFPLA_NET_0_117146, Y => HIEFFPLA_NET_0_116051);
    
    HIEFFPLA_INST_0_43151 : AO1D
      port map(A => HIEFFPLA_NET_0_119451, B => 
        \U50_PATTERNS/REG_STATE[5]_net_1\, C => 
        HIEFFPLA_NET_0_119345, Y => HIEFFPLA_NET_0_119360);
    
    HIEFFPLA_INST_0_37846 : AND3A
      port map(A => \U200B_ELINKS/N_232_li\, B => 
        HIEFFPLA_NET_0_120233, C => 
        \U200B_ELINKS/GP_PG_SM[9]_net_1\, Y => 
        HIEFFPLA_NET_0_120192);
    
    \U_TFC_CMD_TX/SER_OUT_RI\ : DFN1C0
      port map(D => \U_TFC_CMD_TX/SER_CMD_WORD_R[3]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_TFC_CMD_TX/SER_OUT_RI_net_1\);
    
    \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_2S_22\ : DFN1C0
      port map(D => 
        \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_1S_0_net_1\, CLK
         => CLK60MHZ, CLR => \U_EXEC_MASTER/P_MASTER_POR_B_c_0\, 
        Q => P_USB_MASTER_EN_c_22);
    
    HIEFFPLA_INST_0_62923 : MX2
      port map(A => HIEFFPLA_NET_0_115892, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[2]\, S => 
        HIEFFPLA_NET_0_117073, Y => HIEFFPLA_NET_0_115928);
    
    \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[10]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117720, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_33, Q => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[10]_net_1\);
    
    HIEFFPLA_INST_0_51833 : AND2B
      port map(A => \U_MASTER_DES/U13A_ADJ_160M/BITCNT[0]\, B => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[2]\, Y => 
        HIEFFPLA_NET_0_117681);
    
    \U50_PATTERNS/ELINKS_STOP_ADDR_T[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120115, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_7, Q => 
        \U50_PATTERNS/ELINKS_STOP_ADDR_T[4]\);
    
    HIEFFPLA_INST_0_47222 : MX2
      port map(A => HIEFFPLA_NET_0_118537, B => 
        HIEFFPLA_NET_0_118533, S => \BIT_OS_SEL_4[1]\, Y => 
        HIEFFPLA_NET_0_118532);
    
    HIEFFPLA_INST_0_43835 : MX2
      port map(A => HIEFFPLA_NET_0_119522, B => 
        \U50_PATTERNS/TFC_ADDRA[2]\, S => HIEFFPLA_NET_0_119294, 
        Y => HIEFFPLA_NET_0_119205);
    
    \U_ELK17_CH/U_SLAVE_1ELK/Q[9]\ : DFN1C0
      port map(D => \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/Q[9]_net_1\);
    
    HIEFFPLA_INST_0_43619 : NAND3C
      port map(A => \U50_PATTERNS/SM_BANK_SEL[7]\, B => 
        \U50_PATTERNS/SM_BANK_SEL[3]\, C => HIEFFPLA_NET_0_119274, 
        Y => HIEFFPLA_NET_0_119266);
    
    HIEFFPLA_INST_0_38394 : MX2
      port map(A => \U50_PATTERNS/ELINKS_STRT_ADDR[3]\, B => 
        \U50_PATTERNS/ELINKS_STRT_ADDR_T[3]\, S => 
        HIEFFPLA_NET_0_119472, Y => HIEFFPLA_NET_0_120108);
    
    \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[9]\ : DFN1C0
      port map(D => \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\);
    
    \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[9]\ : DFN1C0
      port map(D => 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\);
    
    HIEFFPLA_INST_0_41942 : NAND2
      port map(A => HIEFFPLA_NET_0_119389, B => 
        \U50_PATTERNS/SM_BANK_SEL[2]\, Y => HIEFFPLA_NET_0_119652);
    
    \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[10]\ : DFN1C0
      port map(D => 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]_net_1\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\);
    
    \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[34]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117715, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_33, Q => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[34]_net_1\);
    
    \U50_PATTERNS/ELINK_RWA[3]/U1\ : DFN1P0
      port map(D => HIEFFPLA_NET_0_119698, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_6, Q => \U50_PATTERNS/ELINK_RWA[3]\);
    
    \U200B_ELINKS/LOC_STOP_ADDR[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120184, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_7, Q => 
        \U200B_ELINKS/LOC_STOP_ADDR[3]\);
    
    HIEFFPLA_INST_0_53328 : AND3A
      port map(A => \BIT_OS_SEL_1[0]\, B => HIEFFPLA_NET_0_117425, 
        C => \BIT_OS_SEL_1[2]\, Y => HIEFFPLA_NET_0_117428);
    
    HIEFFPLA_INST_0_44512 : MX2B
      port map(A => HIEFFPLA_NET_0_119103, B => 
        HIEFFPLA_NET_0_119114, S => 
        \U50_PATTERNS/U4C_REGCROSS/SYNC_SM[0]_net_1\, Y => 
        HIEFFPLA_NET_0_119104);
    
    HIEFFPLA_INST_0_39389 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_2[3]\, B => 
        HIEFFPLA_NET_0_119520, S => HIEFFPLA_NET_0_119278, Y => 
        HIEFFPLA_NET_0_119996);
    
    \U50_PATTERNS/ELINK_DINA_10[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119860, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_9, Q => 
        \U50_PATTERNS/ELINK_DINA_10[3]\);
    
    HIEFFPLA_INST_0_43910 : MX2
      port map(A => HIEFFPLA_NET_0_119576, B => 
        \U50_PATTERNS/TFC_DINA[1]\, S => HIEFFPLA_NET_0_119294, Y
         => HIEFFPLA_NET_0_119196);
    
    HIEFFPLA_INST_0_40927 : MX2
      port map(A => HIEFFPLA_NET_0_119567, B => 
        \U50_PATTERNS/ELINK_DINA_18[5]\, S => 
        HIEFFPLA_NET_0_119264, Y => HIEFFPLA_NET_0_119794);
    
    HIEFFPLA_INST_0_57984 : NAND2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_7[0]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_7[1]\, Y => 
        HIEFFPLA_NET_0_116584);
    
    \U_TFC_SERDAT_SOURCE/SERDAT[1]\ : DFN1C0
      port map(D => \U_TFC_SERDAT_SOURCE/N_SERDAT[1]\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \TFC_TX_DAT[1]\);
    
    \U50_PATTERNS/CHKSUM[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120142, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_3, Q => \U50_PATTERNS/CHKSUM[1]\);
    
    HIEFFPLA_INST_0_60468 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_11[3]\, B => 
        HIEFFPLA_NET_0_117075, S => HIEFFPLA_NET_0_117348, Y => 
        HIEFFPLA_NET_0_116262);
    
    HIEFFPLA_INST_0_40036 : MX2
      port map(A => HIEFFPLA_NET_0_119890, B => 
        \U50_PATTERNS/ELINK_BLKA[4]\, S => 
        \U50_PATTERNS/SM_BANK_SEL[20]\, Y => 
        HIEFFPLA_NET_0_119921);
    
    \U50_PATTERNS/U4E_REGCROSS/LOCAL_REG_VAL[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119064, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_6, Q => \OP_MODE_c[6]\);
    
    HIEFFPLA_INST_0_57426 : NAND2B
      port map(A => HIEFFPLA_NET_0_116593, B => 
        HIEFFPLA_NET_0_116678, Y => HIEFFPLA_NET_0_116687);
    
    HIEFFPLA_INST_0_37495 : MX2
      port map(A => \U200A_TFC/LOC_STRT_ADDR[7]\, B => 
        \TFC_STRT_ADDR[7]\, S => \U200A_TFC/GP_PG_SM[10]_net_1\, 
        Y => HIEFFPLA_NET_0_120275);
    
    HIEFFPLA_INST_0_60072 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_6[0]\, B => 
        HIEFFPLA_NET_0_116310, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_0[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116314);
    
    HIEFFPLA_INST_0_111418 : AND3A
      port map(A => HIEFFPLA_NET_0_115838, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[0]_net_1\, C => 
        HIEFFPLA_NET_0_117593, Y => HIEFFPLA_NET_0_117584);
    
    \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[5]\ : DFN1C0
      port map(D => \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_17[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116500, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_18, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_17[1]\);
    
    HIEFFPLA_INST_0_60935 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_1[4]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_17[4]\, S
         => \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_3[4]_net_1\, 
        Y => HIEFFPLA_NET_0_116196);
    
    HIEFFPLA_INST_0_57661 : XA1C
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_5[4]\, B => 
        HIEFFPLA_NET_0_116647, C => HIEFFPLA_NET_0_117179, Y => 
        HIEFFPLA_NET_0_116640);
    
    HIEFFPLA_INST_0_38130 : AX1C
      port map(A => \ELKS_ADDRB[6]\, B => HIEFFPLA_NET_0_120144, 
        C => \ELKS_ADDRB[7]\, Y => HIEFFPLA_NET_0_120147);
    
    \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[2]\ : DFN1C0
      port map(D => 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[2]_net_1\);
    
    HIEFFPLA_INST_0_41665 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_9[7]\, B => 
        HIEFFPLA_NET_0_119560, S => HIEFFPLA_NET_0_119292, Y => 
        HIEFFPLA_NET_0_119712);
    
    HIEFFPLA_INST_0_59546 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_12[2]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_28[2]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[4]_net_1\, Y
         => HIEFFPLA_NET_0_116380);
    
    HIEFFPLA_INST_0_57830 : XA1C
      port map(A => HIEFFPLA_NET_0_116617, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_6[4]\, C => 
        HIEFFPLA_NET_0_117179, Y => HIEFFPLA_NET_0_116611);
    
    \U50_PATTERNS/ELINK_ADDRA_15[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120041, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_6, Q => 
        \U50_PATTERNS/ELINK_ADDRA_15[6]\);
    
    \U_ELK13_CH/U_SLAVE_1ELK/Q[4]\ : DFN1C0
      port map(D => \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/Q[4]_net_1\);
    
    HIEFFPLA_INST_0_59148 : AO1B
      port map(A => HIEFFPLA_NET_0_117254, B => 
        HIEFFPLA_NET_0_116425, C => HIEFFPLA_NET_0_117263, Y => 
        HIEFFPLA_NET_0_116429);
    
    HIEFFPLA_INST_0_51719 : NAND2B
      port map(A => 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM[4]_net_1\, B => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[72]_net_1\, Y => 
        HIEFFPLA_NET_0_117707);
    
    \U_MASTER_DES/U13C_MASTER_DESER/Q[2]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[2]_net_1\, CLK => 
        CCC_160M_FXD, CLR => P_MASTER_POR_B_c_34, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/Q[2]_net_1\);
    
    \U_ELK19_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118242, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_4, Q => 
        \U_ELK19_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]_net_1\);
    
    HIEFFPLA_INST_0_40143 : AOI1C
      port map(A => \U50_PATTERNS/ELINK_BLKA[3]\, B => 
        HIEFFPLA_NET_0_119645, C => HIEFFPLA_NET_0_119891, Y => 
        HIEFFPLA_NET_0_119892);
    
    HIEFFPLA_INST_0_62021 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_29[0]\, B => 
        HIEFFPLA_NET_0_117096, S => HIEFFPLA_NET_0_117072, Y => 
        HIEFFPLA_NET_0_116045);
    
    \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[8]\ : DFN1C0
      port map(D => \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\);
    
    HIEFFPLA_INST_0_48362 : MX2
      port map(A => 
        \U_ELK17_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]_net_1\, B => 
        \U_ELK17_CH/ELK_TX_DAT[7]\, S => 
        \U_ELK17_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118330);
    
    \U50_PATTERNS/REG_STATE[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119468, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_22_0, Q => 
        \U50_PATTERNS/REG_STATE[1]_net_1\);
    
    HIEFFPLA_INST_0_62137 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_2[4]\, 
        B => HIEFFPLA_NET_0_117166, S => HIEFFPLA_NET_0_117176, Y
         => HIEFFPLA_NET_0_116031);
    
    \U_ELK4_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]\ : DFN1C0
      port map(D => \U_ELK4_CH/U_SLAVE_1ELK/Q[1]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]_net_1\);
    
    \U50_PATTERNS/ELINK_DINA_10[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119856, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_9, Q => 
        \U50_PATTERNS/ELINK_DINA_10[7]\);
    
    HIEFFPLA_INST_0_44338 : XOR2
      port map(A => \U50_PATTERNS/U4A_REGCROSS/DELCNT[0]_net_1\, 
        B => \U50_PATTERNS/U4A_REGCROSS/DELCNT[1]_net_1\, Y => 
        HIEFFPLA_NET_0_119136);
    
    HIEFFPLA_INST_0_48854 : MX2
      port map(A => 
        \U_ELK19_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]_net_1\, B => 
        \U_ELK19_CH/ELK_TX_DAT[5]\, S => 
        \U_ELK19_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118241);
    
    \U_ELK9_CH/U_SLAVE_1ELK/Q[6]\ : DFN1C0
      port map(D => \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/Q[6]_net_1\);
    
    HIEFFPLA_INST_0_49320 : MX2
      port map(A => \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\, 
        B => \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[14]_net_1\, S => 
        \BIT_OS_SEL_1[2]\, Y => HIEFFPLA_NET_0_118158);
    
    \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[6]\ : DFN1C0
      port map(D => \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\);
    
    \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[11]\ : DFN1C0
      port map(D => \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\);
    
    HIEFFPLA_INST_0_43137 : AOI1A
      port map(A => HIEFFPLA_NET_0_119387, B => 
        HIEFFPLA_NET_0_119360, C => HIEFFPLA_NET_0_119362, Y => 
        HIEFFPLA_NET_0_119363);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_10[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116272, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_18, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_10[3]\);
    
    \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[7]\ : DFN1C0
      port map(D => \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\);
    
    HIEFFPLA_INST_0_46959 : MX2
      port map(A => HIEFFPLA_NET_0_118590, B => 
        HIEFFPLA_NET_0_118587, S => \BIT_OS_SEL_4[1]\, Y => 
        HIEFFPLA_NET_0_118579);
    
    HIEFFPLA_INST_0_45468 : AO1
      port map(A => HIEFFPLA_NET_0_119250, B => 
        \U50_PATTERNS/ELINK_DOUTA_5[5]\, C => 
        HIEFFPLA_NET_0_118815, Y => HIEFFPLA_NET_0_118908);
    
    \U_ELK19_CH/U_SLAVE_1ELK/Q[6]\ : DFN1C0
      port map(D => \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/Q[6]_net_1\);
    
    \U_ELK3_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U0\ : IOPADP_BI
      port map(N2PIN => 
        \U_ELK3_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2_N2P\, D => 
        \U_ELK3_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, E => 
        \U_ELK3_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET2\, PAD => 
        ELK3_DAT_P, Y => 
        \U_ELK3_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\);
    
    \U50_PATTERNS/U4A_REGCROSS/SAMP_TWO[0]\ : DFN1C0
      port map(D => \U50_PATTERNS/U4A_REGCROSS/SAMP_ONE[0]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_21, Q => 
        \U50_PATTERNS/U4A_REGCROSS/SAMP_TWO[0]_net_1\);
    
    \U200B_ELINKS/RX_SER_WORD_1DEL[7]\ : DFN1C0
      port map(D => \ELK_RX_SER_WORD_0[7]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_23, Q => 
        \U200B_ELINKS/RX_SER_WORD_1DEL[7]_net_1\);
    
    \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[6]\ : DFN1C0
      port map(D => \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\);
    
    \U_ELK5_CH/ELK_IN_R\ : DFN1C0
      port map(D => \U_ELK5_CH/ELK_IN_DDR_R\, CLK => CCC_160M_ADJ, 
        CLR => DEV_RST_B_c, Q => \U_ELK5_CH/ELK_IN_R_net_1\);
    
    \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[8]\ : DFN1C0
      port map(D => \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\);
    
    HIEFFPLA_INST_0_59168 : AO1C
      port map(A => HIEFFPLA_NET_0_117208, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_24[1]\, C => 
        HIEFFPLA_NET_0_117264, Y => HIEFFPLA_NET_0_116425);
    
    HIEFFPLA_INST_0_46668 : MX2
      port map(A => HIEFFPLA_NET_0_118631, B => 
        HIEFFPLA_NET_0_118626, S => \BIT_OS_SEL_5[1]\, Y => 
        HIEFFPLA_NET_0_118630);
    
    \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[13]\ : DFN1C0
      port map(D => \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[13]_net_1\);
    
    HIEFFPLA_INST_0_52716 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_25[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_26[1]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_3[0]\, Y => 
        HIEFFPLA_NET_0_117523);
    
    \U200A_TFC/RX_SER_WORD_1DEL[6]\ : DFN1C0
      port map(D => \TFC_RX_SER_WORD[6]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_31, Q => 
        \U200A_TFC/RX_SER_WORD_1DEL[6]_net_1\);
    
    HIEFFPLA_INST_0_44546 : XOR2
      port map(A => \U50_PATTERNS/U4C_REGCROSS/DELCNT[0]_net_1\, 
        B => \U50_PATTERNS/U4C_REGCROSS/DELCNT[1]_net_1\, Y => 
        HIEFFPLA_NET_0_119094);
    
    \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[10]\ : DFN1C0
      port map(D => 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]_net_1\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\);
    
    HIEFFPLA_INST_0_50784 : MX2
      port map(A => HIEFFPLA_NET_0_117913, B => 
        HIEFFPLA_NET_0_117890, S => \BIT_OS_SEL[0]\, Y => 
        \U_ELK7_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[7]\);
    
    \U200A_TFC/GP_PG_SM[4]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120317, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_28, Q => 
        \U200A_TFC/GP_PG_SM[4]_net_1\);
    
    HIEFFPLA_INST_0_52920 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_23[3]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_24[3]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_2[0]\, Y => 
        HIEFFPLA_NET_0_117489);
    
    HIEFFPLA_INST_0_40882 : MX2
      port map(A => HIEFFPLA_NET_0_119578, B => 
        \U50_PATTERNS/ELINK_DINA_18[0]\, S => 
        HIEFFPLA_NET_0_119264, Y => HIEFFPLA_NET_0_119799);
    
    HIEFFPLA_INST_0_62838 : MX2
      port map(A => HIEFFPLA_NET_0_115878, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/TUNE_CLKPHASE[4]\, S => 
        HIEFFPLA_NET_0_117102, Y => HIEFFPLA_NET_0_115938);
    
    HIEFFPLA_INST_0_62538 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_7[3]\, 
        B => HIEFFPLA_NET_0_117075, S => HIEFFPLA_NET_0_117174, Y
         => HIEFFPLA_NET_0_115977);
    
    \U_ELK13_CH/U_ELK1_SERDAT_SOURCE/SERDAT[4]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118504, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_4, Q => 
        \U_ELK13_CH/ELK_TX_DAT[4]\);
    
    \U50_PATTERNS/CHKSUM[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120137, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_4, Q => \U50_PATTERNS/CHKSUM[6]\);
    
    \U200B_ELINKS/RX_SER_WORD_2DEL[0]\ : DFN1C0
      port map(D => \U200B_ELINKS/RX_SER_WORD_1DEL[0]_net_1\, CLK
         => CLK_40M_GL, CLR => P_MASTER_POR_B_c_25, Q => 
        \U200B_ELINKS/RX_SER_WORD_2DEL[0]_net_1\);
    
    HIEFFPLA_INST_0_47626 : NAND2B
      port map(A => \OP_MODE_c_2[1]\, B => \PATT_ELK_DAT_14[7]\, 
        Y => HIEFFPLA_NET_0_118456);
    
    HIEFFPLA_INST_0_46619 : MX2
      port map(A => 
        \U_ELK10_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]_net_1\, B => 
        \U_ELK10_CH/ELK_TX_DAT[7]\, S => 
        \U_ELK10_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118645);
    
    HIEFFPLA_INST_0_54237 : MX2
      port map(A => HIEFFPLA_NET_0_116566, B => 
        HIEFFPLA_NET_0_116288, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_1[3]_net_1\, Y
         => HIEFFPLA_NET_0_117291);
    
    HIEFFPLA_INST_0_44248 : MX2
      port map(A => \TFC_STRT_ADDR[1]\, B => 
        \U50_PATTERNS/U4A_REGCROSS/SAMP_TWO[1]_net_1\, S => 
        HIEFFPLA_NET_0_119156, Y => HIEFFPLA_NET_0_119153);
    
    HIEFFPLA_INST_0_61817 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_10[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_26[1]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_4[4]_net_1\, Y
         => HIEFFPLA_NET_0_116074);
    
    HIEFFPLA_INST_0_38354 : MX2
      port map(A => \U50_PATTERNS/ELINKS_STOP_ADDR_T[6]\, B => 
        \U50_PATTERNS/RD_USB_ADBUS[6]\, S => 
        HIEFFPLA_NET_0_119413, Y => HIEFFPLA_NET_0_120113);
    
    \U_ELK11_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]\ : DFN1C0
      port map(D => \U_ELK11_CH/U_SLAVE_1ELK/Q[7]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]_net_1\);
    
    HIEFFPLA_INST_0_38306 : MX2
      port map(A => \U50_PATTERNS/ELINKS_STOP_ADDR_T[0]\, B => 
        \U50_PATTERNS/RD_USB_ADBUS[0]\, S => 
        HIEFFPLA_NET_0_119413, Y => HIEFFPLA_NET_0_120119);
    
    HIEFFPLA_INST_0_44142 : MX2
      port map(A => \U50_PATTERNS/TFC_STRT_ADDR[4]\, B => 
        \U50_PATTERNS/TFC_STRT_ADDR_T[4]\, S => 
        HIEFFPLA_NET_0_119472, Y => HIEFFPLA_NET_0_119168);
    
    \U50_PATTERNS/CHKSUM[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120136, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_4, Q => \U50_PATTERNS/CHKSUM[7]\);
    
    HIEFFPLA_INST_0_46837 : MX2
      port map(A => 
        \U_ELK11_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]_net_1\, B => 
        \U_ELK11_CH/ELK_TX_DAT[2]\, S => 
        \U_ELK11_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118606);
    
    \U_ELK9_CH/U_SLAVE_1ELK/RECD_SER_WORD[7]\ : DFN1C0
      port map(D => \U_ELK9_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[7]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_9[7]\);
    
    \U_ELK3_CH/U_ELK1_SERDAT_SOURCE/SERDAT[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118102, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_15, Q => 
        \U_ELK3_CH/ELK_TX_DAT[1]\);
    
    HIEFFPLA_INST_0_61550 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_23[0]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_24[0]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[0]\, Y => 
        HIEFFPLA_NET_0_116111);
    
    HIEFFPLA_INST_0_42928 : NAND2A
      port map(A => \U50_PATTERNS/REG_STATE[5]_net_1\, B => 
        \U50_PATTERNS/REG_STATE[4]_net_1\, Y => 
        HIEFFPLA_NET_0_119422);
    
    HIEFFPLA_INST_0_56899 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_1[8]\, B => 
        HIEFFPLA_NET_0_116759, S => HIEFFPLA_NET_0_117600, Y => 
        HIEFFPLA_NET_0_116780);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_18[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116492, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_19, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_18[3]\);
    
    \U50_PATTERNS/SM_BANK_SEL_0[21]/U1\ : DFN1P0
      port map(D => HIEFFPLA_NET_0_119299, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_2_0, Q => 
        \U50_PATTERNS/SM_BANK_SEL_0[21]\);
    
    HIEFFPLA_INST_0_38849 : MX2
      port map(A => HIEFFPLA_NET_0_119516, B => 
        \U50_PATTERNS/ELINK_ADDRA_13[7]\, S => 
        HIEFFPLA_NET_0_119285, Y => HIEFFPLA_NET_0_120056);
    
    \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[6]\ : DFN1C0
      port map(D => \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\);
    
    \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[11]\ : DFN1C0
      port map(D => \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\);
    
    HIEFFPLA_INST_0_39893 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_9[3]\, B => 
        HIEFFPLA_NET_0_119520, S => HIEFFPLA_NET_0_119292, Y => 
        HIEFFPLA_NET_0_119940);
    
    \U50_PATTERNS/ELINK_DINA_4[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119752, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_13, Q => 
        \U50_PATTERNS/ELINK_DINA_4[7]\);
    
    HIEFFPLA_INST_0_58013 : AND3B
      port map(A => HIEFFPLA_NET_0_116574, B => 
        HIEFFPLA_NET_0_117179, C => HIEFFPLA_NET_0_116585, Y => 
        HIEFFPLA_NET_0_116578);
    
    HIEFFPLA_INST_0_48346 : AND2
      port map(A => \U_ELK17_CH/ELK_TX_DAT[1]\, B => 
        \U_ELK17_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118333);
    
    HIEFFPLA_INST_0_61793 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_26[3]\, B => 
        HIEFFPLA_NET_0_117075, S => HIEFFPLA_NET_0_117138, Y => 
        HIEFFPLA_NET_0_116077);
    
    HIEFFPLA_INST_0_39677 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_6[3]\, B => 
        HIEFFPLA_NET_0_119520, S => HIEFFPLA_NET_0_119258, Y => 
        HIEFFPLA_NET_0_119964);
    
    HIEFFPLA_INST_0_37033 : AOI1A
      port map(A => HIEFFPLA_NET_0_120351, B => 
        HIEFFPLA_NET_0_120325, C => HIEFFPLA_NET_0_120363, Y => 
        HIEFFPLA_NET_0_120364);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_21[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116455, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_14, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_21[1]\);
    
    HIEFFPLA_INST_0_42010 : AOI1C
      port map(A => \U50_PATTERNS/ELK_N_ACTIVE_net_1\, B => 
        \U50_PATTERNS/SM_BANK_SEL[20]\, C => 
        \U50_PATTERNS/SM_BANK_SEL_0[21]\, Y => 
        HIEFFPLA_NET_0_119632);
    
    HIEFFPLA_INST_0_52252 : AO1
      port map(A => HIEFFPLA_NET_0_117590, B => 
        HIEFFPLA_NET_0_117596, C => HIEFFPLA_NET_0_117179, Y => 
        HIEFFPLA_NET_0_117600);
    
    HIEFFPLA_INST_0_49563 : MX2
      port map(A => \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[0]_net_1\, B
         => \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\, S => 
        \BIT_OS_SEL_7[2]\, Y => HIEFFPLA_NET_0_118114);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_9[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_115962, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_20, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_9[3]\);
    
    \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[5]\ : DFN1C0
      port map(D => \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\);
    
    HIEFFPLA_INST_0_58509 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_16[0]\, B => 
        HIEFFPLA_NET_0_116508, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_1[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116512);
    
    HIEFFPLA_INST_0_54405 : MX2
      port map(A => HIEFFPLA_NET_0_116209, B => 
        HIEFFPLA_NET_0_116099, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_2[3]_net_1\, Y
         => HIEFFPLA_NET_0_117270);
    
    HIEFFPLA_INST_0_44988 : AND3B
      port map(A => HIEFFPLA_NET_0_119451, B => 
        \U50_PATTERNS/USB_TXE_B\, C => 
        \U50_PATTERNS/REG_STATE[0]_net_1\, Y => 
        HIEFFPLA_NET_0_119006);
    
    \U50_PATTERNS/ELINK_ADDRA_4[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119977, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_2_0, Q => 
        \U50_PATTERNS/ELINK_ADDRA_4[6]\);
    
    HIEFFPLA_INST_0_50945 : MX2
      port map(A => HIEFFPLA_NET_0_117861, B => 
        HIEFFPLA_NET_0_117857, S => \BIT_OS_SEL_3[1]\, Y => 
        HIEFFPLA_NET_0_117859);
    
    \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[10]\ : DFN1C0
      port map(D => 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]_net_1\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\);
    
    HIEFFPLA_INST_0_60606 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_13[4]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_14[4]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_3[0]\, Y => 
        HIEFFPLA_NET_0_116245);
    
    HIEFFPLA_INST_0_42077 : AO1A
      port map(A => HIEFFPLA_NET_0_119622, B => 
        \U50_PATTERNS/TFC_STOP_ADDR[3]\, C => 
        HIEFFPLA_NET_0_118670, Y => HIEFFPLA_NET_0_119620);
    
    \U_ELK18_CH/U_SLAVE_1ELK/Q[7]\ : DFN1C0
      port map(D => \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/Q[7]_net_1\);
    
    HIEFFPLA_INST_0_48736 : MX2
      port map(A => HIEFFPLA_NET_0_118251, B => 
        HIEFFPLA_NET_0_118264, S => \BIT_OS_SEL_2[0]\, Y => 
        \U_ELK18_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[0]\);
    
    \U_ELK18_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118290, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_3, Q => 
        \U_ELK18_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]_net_1\);
    
    HIEFFPLA_INST_0_60203 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_7[3]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_23[3]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_4[4]_net_1\, Y
         => HIEFFPLA_NET_0_116296);
    
    HIEFFPLA_INST_0_46396 : AO1
      port map(A => HIEFFPLA_NET_0_119244, B => 
        \U50_PATTERNS/ELINK_DOUTA_2[4]\, C => 
        HIEFFPLA_NET_0_118841, Y => HIEFFPLA_NET_0_118699);
    
    \U_ELK8_CH/U_SLAVE_1ELK/Q[6]\ : DFN1C0
      port map(D => \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/Q[6]_net_1\);
    
    HIEFFPLA_INST_0_48423 : MX2
      port map(A => HIEFFPLA_NET_0_118314, B => 
        HIEFFPLA_NET_0_118311, S => \BIT_OS_SEL_1[1]\, Y => 
        HIEFFPLA_NET_0_118313);
    
    HIEFFPLA_INST_0_38370 : MX2
      port map(A => \U50_PATTERNS/ELINKS_STRT_ADDR[0]\, B => 
        \U50_PATTERNS/ELINKS_STRT_ADDR_T[0]\, S => 
        HIEFFPLA_NET_0_119472, Y => HIEFFPLA_NET_0_120111);
    
    \U_EXEC_MASTER/USB_MASTER_EN/T_CNT60M[5]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117738, CLK => CLK60MHZ, CLR
         => P_MASTER_POR_B_c_28, Q => 
        \U_EXEC_MASTER/USB_MASTER_EN/T_CNT60M[5]_net_1\);
    
    \U50_PATTERNS/U4A_REGCROSS/SAMP_ONE[4]\ : DFN1C0
      port map(D => \U50_PATTERNS/TFC_STRT_ADDR[4]\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_32_0, Q => 
        \U50_PATTERNS/U4A_REGCROSS/SAMP_ONE[4]_net_1\);
    
    \U200A_TFC/ADDR_POINTER[5]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120358, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_30, Q => \TFC_ADDRB[5]\);
    
    HIEFFPLA_INST_0_112149 : AOI1A
      port map(A => HIEFFPLA_NET_0_120190, B => 
        HIEFFPLA_NET_0_120231, C => 
        \U200B_ELINKS/GP_PG_SM[10]_net_1\, Y => 
        HIEFFPLA_NET_0_115819);
    
    \U50_PATTERNS/OP_MODE[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119613, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_15, Q => \U50_PATTERNS/OP_MODE[4]\);
    
    HIEFFPLA_INST_0_58431 : MX2
      port map(A => HIEFFPLA_NET_0_116687, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_14[2]\, S => 
        HIEFFPLA_NET_0_117219, Y => HIEFFPLA_NET_0_116522);
    
    HIEFFPLA_INST_0_53738 : MX2
      port map(A => HIEFFPLA_NET_0_117379, B => 
        HIEFFPLA_NET_0_117293, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[2]_net_1\, Y
         => HIEFFPLA_NET_0_117362);
    
    \U_ELK19_CH/U_SLAVE_1ELK/Q[4]\ : DFN1C0
      port map(D => \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/Q[4]_net_1\);
    
    HIEFFPLA_INST_0_47864 : MX2
      port map(A => 
        \U_ELK15_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]_net_1\, B => 
        \U_ELK15_CH/ELK_TX_DAT[7]\, S => 
        \U_ELK15_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118420);
    
    HIEFFPLA_INST_0_42230 : NAND3C
      port map(A => \U50_PATTERNS/RD_USB_ADBUS[6]\, B => 
        HIEFFPLA_NET_0_119020, C => 
        \U50_PATTERNS/RD_USB_ADBUS[5]\, Y => 
        HIEFFPLA_NET_0_119598);
    
    \U_ELK9_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]\ : DFN1C0
      port map(D => \U_ELK9_CH/U_SLAVE_1ELK/Q[10]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]_net_1\);
    
    \U_DDR_TFC/BIBUF_LVDS_0/U0/U3\ : IOBI_ID_OD_EB
      port map(DR => TFC_OUT_R, DF => TFC_OUT_F, CLR => \GND\, E
         => DCB_SALT_SEL_c, ICLK => CCC_160M_ADJ, OCLK => 
        CCC_160M_FXD, YIN => \U_DDR_TFC/BIBUF_LVDS_0/U0/NET4\, 
        DOUT => OPEN, EOUT => \U_DDR_TFC/BIBUF_LVDS_0/U0/NET3\, 
        YR => OPEN, YF => OPEN);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_12[4]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116251, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_21, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_12[4]\);
    
    HIEFFPLA_INST_0_53632 : MX2
      port map(A => HIEFFPLA_NET_0_116686, B => 
        HIEFFPLA_NET_0_116649, S => HIEFFPLA_NET_0_117325, Y => 
        HIEFFPLA_NET_0_117380);
    
    \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_SEL_5[2]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_BIT_OS_VAL[2]\, CLK
         => CLK_40M_GL, CLR => P_MASTER_POR_B_c_27_0, Q => 
        \BIT_OS_SEL_5[2]\);
    
    HIEFFPLA_INST_0_47123 : NAND2B
      port map(A => \OP_MODE_c_3[1]\, B => \PATT_ELK_DAT_12[2]\, 
        Y => HIEFFPLA_NET_0_118551);
    
    HIEFFPLA_INST_0_52045 : MX2
      port map(A => HIEFFPLA_NET_0_117638, B => 
        HIEFFPLA_NET_0_117637, S => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[1]\, Y => 
        HIEFFPLA_NET_0_117647);
    
    HIEFFPLA_INST_0_50365 : NAND2B
      port map(A => \OP_MODE_c_1[1]\, B => \PATT_ELK_DAT_6[7]\, Y
         => HIEFFPLA_NET_0_117961);
    
    HIEFFPLA_INST_0_52151 : AND3B
      port map(A => \U_MASTER_DES/U13A_ADJ_160M/BITCNT[7]\, B => 
        HIEFFPLA_NET_0_117687, C => 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM[2]_net_1\, Y => 
        HIEFFPLA_NET_0_117624);
    
    \U_ELK17_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]\ : DFN1C0
      port map(D => \U_ELK17_CH/U_SLAVE_1ELK/Q[11]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]_net_1\);
    
    HIEFFPLA_INST_0_49812 : MX2
      port map(A => \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[0]_net_1\, B
         => \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\, S => 
        \BIT_OS_SEL_7[2]\, Y => HIEFFPLA_NET_0_118069);
    
    HIEFFPLA_INST_0_43187 : AOI1C
      port map(A => \U50_PATTERNS/REG_STATE[3]_net_1\, B => 
        \U50_PATTERNS/REG_STATE_0[2]_net_1\, C => 
        HIEFFPLA_NET_0_119380, Y => HIEFFPLA_NET_0_119352);
    
    HIEFFPLA_INST_0_46623 : AND2A
      port map(A => \OP_MODE_c_3[1]\, B => \PATT_ELK_DAT_10[0]\, 
        Y => HIEFFPLA_NET_0_118643);
    
    \U50_PATTERNS/TFC_STRT_ADDR_T[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119160, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_4, Q => 
        \U50_PATTERNS/TFC_STRT_ADDR_T[4]\);
    
    HIEFFPLA_INST_0_40008 : MX2
      port map(A => HIEFFPLA_NET_0_119898, B => 
        \U50_PATTERNS/ELINK_BLKA[19]\, S => 
        \U50_PATTERNS/SM_BANK_SEL[20]\, Y => 
        HIEFFPLA_NET_0_119925);
    
    \U50_PATTERNS/TFC_STRT_ADDR[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119170, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_13, Q => 
        \U50_PATTERNS/TFC_STRT_ADDR[2]\);
    
    \U_ELK12_CH/U_ELK1_SERDAT_SOURCE/SERDAT[4]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118549, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_2, Q => 
        \U_ELK12_CH/ELK_TX_DAT[4]\);
    
    HIEFFPLA_INST_0_56487 : AO1
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[7]_net_1\, B => 
        HIEFFPLA_NET_0_117428, C => HIEFFPLA_NET_0_116837, Y => 
        HIEFFPLA_NET_0_116853);
    
    HIEFFPLA_INST_0_45597 : AO1A
      port map(A => HIEFFPLA_NET_0_119475, B => 
        \U50_PATTERNS/ELINKS_STOP_ADDR[6]\, C => 
        HIEFFPLA_NET_0_118775, Y => HIEFFPLA_NET_0_118883);
    
    HIEFFPLA_INST_0_45507 : AND3A
      port map(A => HIEFFPLA_NET_0_119437, B => 
        \U50_PATTERNS/WR_XFER_TYPE[5]_net_1\, C => 
        HIEFFPLA_NET_0_119367, Y => HIEFFPLA_NET_0_118900);
    
    HIEFFPLA_INST_0_56167 : XA1B
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/MAX_CNT[1]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/MAX_CNT[0]\, C => 
        HIEFFPLA_NET_0_117112, Y => HIEFFPLA_NET_0_116938);
    
    AFLSDF_INV_13 : INV
      port map(A => DCB_SALT_SEL_c, Y => \AFLSDF_INV_13\);
    
    HIEFFPLA_INST_0_60250 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_8[2]\, B => 
        HIEFFPLA_NET_0_116687, S => HIEFFPLA_NET_0_117160, Y => 
        HIEFFPLA_NET_0_116291);
    
    \U_ELK3_CH/U_ELK1_SERDAT_SOURCE/SERDAT[4]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118099, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_15, Q => 
        \U_ELK3_CH/ELK_TX_DAT[4]\);
    
    HIEFFPLA_INST_0_38137 : AND2
      port map(A => \ELKS_ADDRB[1]\, B => HIEFFPLA_NET_0_120150, 
        Y => HIEFFPLA_NET_0_120145);
    
    \U_EXEC_MASTER/MPOR_B_12\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117787, CLK => CLK_40M_GL, CLR
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_1\, Q => 
        P_MASTER_POR_B_c_12);
    
    \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[4]\ : DFN1C0
      port map(D => 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\);
    
    \U_ELK18_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U3\ : IOBI_ID_OD_EB
      port map(DR => \U_ELK18_CH/ELK_OUT_R\, DF => 
        \U_ELK18_CH/ELK_OUT_F\, CLR => \GND\, E => 
        \AFLSDF_INV_31\, ICLK => CCC_160M_ADJ, OCLK => 
        CCC_160M_FXD, YIN => 
        \U_ELK18_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\, DOUT => 
        OPEN, EOUT => 
        \U_ELK18_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET3\, YR => OPEN, 
        YF => OPEN);
    
    HIEFFPLA_INST_0_56051 : AND3A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_0[8]_net_1\, B => 
        HIEFFPLA_NET_0_115872, C => HIEFFPLA_NET_0_117027, Y => 
        HIEFFPLA_NET_0_116956);
    
    HIEFFPLA_INST_0_52218 : MX2
      port map(A => ALIGN_ACTIVE, B => \OP_MODE_c[5]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_0[8]_net_1\, Y => 
        HIEFFPLA_NET_0_117609);
    
    \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[6]\ : DFN1C0
      port map(D => \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\);
    
    \U_ELK3_CH/U_SLAVE_1ELK/Q[12]\ : DFN1C0
      port map(D => \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/Q[12]_net_1\);
    
    \U_ELK18_CH/U_SLAVE_1ELK/Q[12]\ : DFN1C0
      port map(D => \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/Q[12]_net_1\);
    
    \U50_PATTERNS/ELINK_DINA_7[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119729, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_17, Q => 
        \U50_PATTERNS/ELINK_DINA_7[6]\);
    
    HIEFFPLA_INST_0_46081 : AND3A
      port map(A => HIEFFPLA_NET_0_119376, B => 
        \U50_PATTERNS/TFC_STRT_ADDR[4]\, C => 
        HIEFFPLA_NET_0_119431, Y => HIEFFPLA_NET_0_118771);
    
    HIEFFPLA_INST_0_42335 : AND3A
      port map(A => \U50_PATTERNS/RD_USB_ADBUS[2]\, B => 
        HIEFFPLA_NET_0_119564, C => 
        \U50_PATTERNS/RD_USB_ADBUS[3]\, Y => 
        HIEFFPLA_NET_0_119568);
    
    HIEFFPLA_INST_0_61451 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_6[1]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_22[1]\, S
         => \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_5[4]_net_1\, 
        Y => HIEFFPLA_NET_0_116125);
    
    HIEFFPLA_INST_0_52230 : AND2A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[1]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[2]_net_1\, Y => 
        HIEFFPLA_NET_0_117605);
    
    \U_ELK19_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118245, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_7, Q => 
        \U_ELK19_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]_net_1\);
    
    \U50_PATTERNS/REG_ADDR[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119528, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_10, Q => \U50_PATTERNS/REG_ADDR[5]\);
    
    \U200A_TFC/RX_SER_WORD_3DEL[3]\ : DFN1P0
      port map(D => \AFLSDF_INV_54\, CLK => CLK_40M_GL, PRE => 
        P_MASTER_POR_B_c_24, Q => 
        \U200A_TFC/RX_SER_WORD_3DEL_i_0[3]\);
    
    \U200A_TFC/LOC_STRT_ADDR[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120280, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_4, Q => \U200A_TFC/LOC_STRT_ADDR[2]\);
    
    \U_ELK12_CH/U_SLAVE_1ELK/RECD_SER_WORD[7]\ : DFN1C0
      port map(D => \U_ELK12_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[7]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_12[7]\);
    
    HIEFFPLA_INST_0_43210 : NAND3C
      port map(A => HIEFFPLA_NET_0_119341, B => 
        HIEFFPLA_NET_0_119337, C => HIEFFPLA_NET_0_119339, Y => 
        HIEFFPLA_NET_0_119347);
    
    \U50_PATTERNS/ELINK_ADDRA_0[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120090, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_18, Q => 
        \U50_PATTERNS/ELINK_ADDRA_0[5]\);
    
    \U_ELK4_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]\ : DFN1C0
      port map(D => \U_ELK4_CH/U_SLAVE_1ELK/Q[6]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]_net_1\);
    
    HIEFFPLA_INST_0_57696 : AOI1A
      port map(A => HIEFFPLA_NET_0_116645, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_5[6]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_5[7]\, Y => 
        HIEFFPLA_NET_0_116633);
    
    HIEFFPLA_INST_0_48621 : AND2A
      port map(A => \OP_MODE_c_2[1]\, B => \PATT_ELK_DAT_18[6]\, 
        Y => HIEFFPLA_NET_0_118277);
    
    \U_MASTER_DES/U13C_MASTER_DESER/ARB_WRD_40M_FIXED[3]\ : 
        DFN1C0
      port map(D => \U_MASTER_DES/U13C_MASTER_DESER/Q[3]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_26, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_WRD_40M_FIXED[3]_net_1\);
    
    \U50_PATTERNS/ELINK_DINA_6[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119740, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_16, Q => 
        \U50_PATTERNS/ELINK_DINA_6[3]\);
    
    \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[10]\ : DFN1C0
      port map(D => \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\);
    
    HIEFFPLA_INST_0_43624 : NAND3C
      port map(A => \U50_PATTERNS/SM_BANK_SEL[8]\, B => 
        \U50_PATTERNS/SM_BANK_SEL[0]\, C => HIEFFPLA_NET_0_119234, 
        Y => HIEFFPLA_NET_0_119265);
    
    HIEFFPLA_INST_0_45195 : NAND3C
      port map(A => HIEFFPLA_NET_0_118959, B => 
        HIEFFPLA_NET_0_118755, C => HIEFFPLA_NET_0_118967, Y => 
        HIEFFPLA_NET_0_118968);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_24[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116104, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_8, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_24[1]\);
    
    HIEFFPLA_INST_0_62824 : AOI1B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[8]_net_1\, B => 
        \OP_MODE_c[5]\, C => HIEFFPLA_NET_0_115936, Y => 
        HIEFFPLA_NET_0_115941);
    
    \U50_PATTERNS/U4C_REGCROSS/SAMP_TWO[0]\ : DFN1C0
      port map(D => \U50_PATTERNS/U4C_REGCROSS/SAMP_ONE[0]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_22_0, Q => 
        \U50_PATTERNS/U4C_REGCROSS/SAMP_TWO[0]_net_1\);
    
    HIEFFPLA_INST_0_50752 : MX2
      port map(A => HIEFFPLA_NET_0_117911, B => 
        HIEFFPLA_NET_0_117906, S => \BIT_OS_SEL_5[0]\, Y => 
        \U_ELK7_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[3]\);
    
    \U200B_ELINKS/LOC_DIR_MODE/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120189, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_2, Q => \U200B_ELINKS/N_232_li\);
    
    HIEFFPLA_INST_0_57349 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_4[1]\, B => 
        HIEFFPLA_NET_0_116670, S => HIEFFPLA_NET_0_117122, Y => 
        HIEFFPLA_NET_0_116695);
    
    HIEFFPLA_INST_0_50128 : MX2
      port map(A => HIEFFPLA_NET_0_117994, B => 
        HIEFFPLA_NET_0_117992, S => \BIT_OS_SEL_6[1]\, Y => 
        HIEFFPLA_NET_0_118004);
    
    HIEFFPLA_INST_0_42149 : MX2
      port map(A => \U50_PATTERNS/OP_MODE[7]\, B => 
        \U50_PATTERNS/OP_MODE_T[7]\, S => HIEFFPLA_NET_0_119472, 
        Y => HIEFFPLA_NET_0_119610);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_4[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116695, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_9, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_4[1]\);
    
    HIEFFPLA_INST_0_60768 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_31[0]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_15[0]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[4]_net_1\, Y
         => HIEFFPLA_NET_0_116223);
    
    HIEFFPLA_INST_0_39065 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_16[7]\, B => 
        HIEFFPLA_NET_0_119516, S => HIEFFPLA_NET_0_119257, Y => 
        HIEFFPLA_NET_0_120032);
    
    \U_ELK6_CH/U_SLAVE_1ELK/RECD_SER_WORD[3]\ : DFN1C0
      port map(D => \U_ELK6_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[3]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_6[3]\);
    
    \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[7]\ : DFN1C0
      port map(D => \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\);
    
    HIEFFPLA_INST_0_51512 : AND3
      port map(A => \U_EXEC_MASTER/CCC_1_LOCK_STAT_1D_net_1\, B
         => HIEFFPLA_NET_0_117764, C => HIEFFPLA_NET_0_117757, Y
         => HIEFFPLA_NET_0_117758);
    
    HIEFFPLA_INST_0_62580 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_7[4]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_8[4]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[0]\, Y => 
        HIEFFPLA_NET_0_115971);
    
    HIEFFPLA_INST_0_58873 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_20[2]\, B => 
        HIEFFPLA_NET_0_116458, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_1[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116465);
    
    HIEFFPLA_INST_0_46541 : MX2
      port map(A => \U_ELK0_CMD_TX/SER_CMD_WORD_F[0]_net_1\, B
         => \ELK0_TX_DAT[2]\, S => 
        \U_ELK0_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118668);
    
    HIEFFPLA_INST_0_44592 : MX2
      port map(A => \ELKS_STOP_ADDR[5]\, B => 
        \U50_PATTERNS/U4D_REGCROSS/SAMP_TWO[5]_net_1\, S => 
        HIEFFPLA_NET_0_119093, Y => HIEFFPLA_NET_0_119086);
    
    \U_ELK14_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]\ : DFN1C0
      port map(D => \U_ELK14_CH/U_SLAVE_1ELK/Q[13]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]_net_1\);
    
    \U_ELK5_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL\ : DFN1C0
      port map(D => 
        \U_ELK5_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL_net_1\);
    
    HIEFFPLA_INST_0_43769 : AND3B
      port map(A => HIEFFPLA_NET_0_119208, B => 
        HIEFFPLA_NET_0_119559, C => HIEFFPLA_NET_0_119562, Y => 
        HIEFFPLA_NET_0_119218);
    
    HIEFFPLA_INST_0_53440 : MX2
      port map(A => HIEFFPLA_NET_0_116461, B => 
        HIEFFPLA_NET_0_116380, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[3]_net_1\, Y
         => HIEFFPLA_NET_0_117408);
    
    HIEFFPLA_INST_0_44818 : AND3
      port map(A => HIEFFPLA_NET_0_119039, B => 
        HIEFFPLA_NET_0_119561, C => HIEFFPLA_NET_0_119568, Y => 
        HIEFFPLA_NET_0_119042);
    
    HIEFFPLA_INST_0_43594 : NAND2B
      port map(A => \U50_PATTERNS/SM_BANK_SEL[15]\, B => 
        \U50_PATTERNS/SM_BANK_SEL[16]\, Y => 
        HIEFFPLA_NET_0_119273);
    
    HIEFFPLA_INST_0_49831 : MX2
      port map(A => 
        \U_ELK4_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]_net_1\, B => 
        \U_ELK4_CH/ELK_TX_DAT[4]\, S => 
        \U_ELK4_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118065);
    
    HIEFFPLA_INST_0_57119 : AND3
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_2[3]\, B => 
        HIEFFPLA_NET_0_116746, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_2[4]\, Y => 
        HIEFFPLA_NET_0_116736);
    
    \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[6]\ : DFN1C0
      port map(D => 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\);
    
    \U_ELK18_CH/U_SLAVE_1ELK/Q[1]\ : DFN1C0
      port map(D => \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/Q[1]_net_1\);
    
    \U50_PATTERNS/TFC_STOP_ADDR[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119188, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_8, Q => 
        \U50_PATTERNS/TFC_STOP_ADDR[0]\);
    
    HIEFFPLA_INST_0_37161 : XO1
      port map(A => HIEFFPLA_NET_0_120256, B => \TFC_ADDRB[6]\, C
         => \U200A_TFC/GP_PG_SM[10]_net_1\, Y => 
        HIEFFPLA_NET_0_120337);
    
    \U_ELK19_CH/U_SLAVE_1ELK/RECD_SER_WORD[7]\ : DFN1C0
      port map(D => \U_ELK19_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[7]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_19[7]\);
    
    \U50_PATTERNS/SM_BANK_SEL[10]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119321, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_1_0, Q => 
        \U50_PATTERNS/SM_BANK_SEL[10]\);
    
    HIEFFPLA_INST_0_57925 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_7[6]\, B => 
        HIEFFPLA_NET_0_116578, S => HIEFFPLA_NET_0_117113, Y => 
        HIEFFPLA_NET_0_116597);
    
    HIEFFPLA_INST_0_43661 : AND2A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/SM_BANK_SEL[14]\, Y => 
        HIEFFPLA_NET_0_119250);
    
    HIEFFPLA_INST_0_46987 : MX2
      port map(A => \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[2]_net_1\, 
        B => \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\, S => 
        \BIT_OS_SEL_4[2]\, Y => HIEFFPLA_NET_0_118575);
    
    HIEFFPLA_INST_0_38840 : MX2
      port map(A => HIEFFPLA_NET_0_119517, B => 
        \U50_PATTERNS/ELINK_ADDRA_13[6]\, S => 
        HIEFFPLA_NET_0_119285, Y => HIEFFPLA_NET_0_120057);
    
    HIEFFPLA_INST_0_53322 : NAND3B
      port map(A => \BIT_OS_SEL[0]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_SEL[3]_net_1\, C
         => \BIT_OS_SEL_1[1]\, Y => HIEFFPLA_NET_0_117430);
    
    HIEFFPLA_INST_0_43315 : NAND2A
      port map(A => HIEFFPLA_NET_0_119330, B => 
        \U50_PATTERNS/SI_CNT[3]\, Y => HIEFFPLA_NET_0_119328);
    
    HIEFFPLA_INST_0_48101 : MX2
      port map(A => 
        \U_ELK16_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]_net_1\, B => 
        \U_ELK16_CH/ELK_TX_DAT[3]\, S => 
        \U_ELK16_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118377);
    
    HIEFFPLA_INST_0_53947 : NAND3
      port map(A => HIEFFPLA_NET_0_117235, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[0]_net_1\, C
         => \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_2[3]_net_1\, 
        Y => HIEFFPLA_NET_0_117329);
    
    \U_ELK6_CH/U_SLAVE_1ELK/Q[10]\ : DFN1C0
      port map(D => \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/Q[10]_net_1\);
    
    \U50_PATTERNS/ELINK_DINA_13[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119834, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_14, Q => 
        \U50_PATTERNS/ELINK_DINA_13[5]\);
    
    \U50_PATTERNS/ELINK_ADDRA_8[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119948, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_8, Q => 
        \U50_PATTERNS/ELINK_ADDRA_8[3]\);
    
    HIEFFPLA_INST_0_52606 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_5[0]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_6[0]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_1[0]\, Y => 
        HIEFFPLA_NET_0_117540);
    
    HIEFFPLA_INST_0_48045 : MX2
      port map(A => HIEFFPLA_NET_0_118396, B => 
        HIEFFPLA_NET_0_118385, S => \BIT_OS_SEL_3[0]\, Y => 
        \U_ELK15_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[7]\);
    
    \U_ELK15_CH/U_ELK1_SERDAT_SOURCE/SERDAT[4]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118414, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_8, Q => 
        \U_ELK15_CH/ELK_TX_DAT[4]\);
    
    HIEFFPLA_INST_0_50302 : MX2
      port map(A => HIEFFPLA_NET_0_117993, B => 
        HIEFFPLA_NET_0_117978, S => \BIT_OS_SEL[1]\, Y => 
        HIEFFPLA_NET_0_117980);
    
    HIEFFPLA_INST_0_44637 : XO1
      port map(A => \ELKS_STOP_ADDR[5]\, B => 
        \U50_PATTERNS/U4D_REGCROSS/SAMP_TWO[5]_net_1\, C => 
        HIEFFPLA_NET_0_119078, Y => HIEFFPLA_NET_0_119079);
    
    HIEFFPLA_INST_0_52710 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_25[0]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_26[0]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_3[0]\, Y => 
        HIEFFPLA_NET_0_117524);
    
    \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[5]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117056, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_27, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[5]_net_1\);
    
    HIEFFPLA_INST_0_57287 : XA1B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_3[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_3[0]\, C => 
        HIEFFPLA_NET_0_117179, Y => HIEFFPLA_NET_0_116707);
    
    \U50_PATTERNS/U112_PATT_ELINK_BLK/DPRT_512X9_SRAM_R0C0\ : 
        RAM4K9
      generic map(MEMORYFILE => "DPRT_512X9_SRAM_R0C0.mem")

      port map(ADDRA11 => AFLSDF_GND, ADDRA10 => AFLSDF_GND, 
        ADDRA9 => AFLSDF_GND, ADDRA8 => \GND\, ADDRA7 => 
        \U50_PATTERNS/ELINK_ADDRA_12[7]\, ADDRA6 => 
        \U50_PATTERNS/ELINK_ADDRA_12[6]\, ADDRA5 => 
        \U50_PATTERNS/ELINK_ADDRA_12[5]\, ADDRA4 => 
        \U50_PATTERNS/ELINK_ADDRA_12[4]\, ADDRA3 => 
        \U50_PATTERNS/ELINK_ADDRA_12[3]\, ADDRA2 => 
        \U50_PATTERNS/ELINK_ADDRA_12[2]\, ADDRA1 => 
        \U50_PATTERNS/ELINK_ADDRA_12[1]\, ADDRA0 => 
        \U50_PATTERNS/ELINK_ADDRA_12[0]\, ADDRB11 => AFLSDF_GND, 
        ADDRB10 => AFLSDF_GND, ADDRB9 => AFLSDF_GND, ADDRB8 => 
        \GND\, ADDRB7 => \ELKS_ADDRB[7]\, ADDRB6 => 
        \ELKS_ADDRB_0[6]\, ADDRB5 => \ELKS_ADDRB[5]\, ADDRB4 => 
        \ELKS_ADDRB_0[4]\, ADDRB3 => \ELKS_ADDRB[3]\, ADDRB2 => 
        \ELKS_ADDRB_0[2]\, ADDRB1 => \ELKS_ADDRB[1]\, ADDRB0 => 
        \ELKS_ADDRB[0]\, DINA8 => \GND\, DINA7 => 
        \U50_PATTERNS/ELINK_DINA_12[7]\, DINA6 => 
        \U50_PATTERNS/ELINK_DINA_12[6]\, DINA5 => 
        \U50_PATTERNS/ELINK_DINA_12[5]\, DINA4 => 
        \U50_PATTERNS/ELINK_DINA_12[4]\, DINA3 => 
        \U50_PATTERNS/ELINK_DINA_12[3]\, DINA2 => 
        \U50_PATTERNS/ELINK_DINA_12[2]\, DINA1 => 
        \U50_PATTERNS/ELINK_DINA_12[1]\, DINA0 => 
        \U50_PATTERNS/ELINK_DINA_12[0]\, DINB8 => \GND\, DINB7
         => \ELK_RX_SER_WORD_12[7]\, DINB6 => 
        \ELK_RX_SER_WORD_12[6]\, DINB5 => \ELK_RX_SER_WORD_12[5]\, 
        DINB4 => \ELK_RX_SER_WORD_12[4]\, DINB3 => 
        \ELK_RX_SER_WORD_12[3]\, DINB2 => \ELK_RX_SER_WORD_12[2]\, 
        DINB1 => \ELK_RX_SER_WORD_12[1]\, DINB0 => 
        \ELK_RX_SER_WORD_12[0]\, WIDTHA0 => \VCC\, WIDTHA1 => 
        \VCC\, WIDTHB0 => \VCC\, WIDTHB1 => \VCC\, PIPEA => \VCC\, 
        PIPEB => \VCC\, WMODEA => \GND\, WMODEB => \GND\, BLKA
         => \U50_PATTERNS/ELINK_BLKA[12]\, BLKB => 
        ELKS_RAM_BLKB_EN, WENA => \U50_PATTERNS/ELINK_RWA[12]\, 
        WENB => ELKS_RWB, CLKA => CLK60MHZ, CLKB => CLK_40M_GL, 
        RESET => P_USB_MASTER_EN_c_0, DOUTA8 => OPEN, DOUTA7 => 
        \U50_PATTERNS/ELINK_DOUTA_12[7]\, DOUTA6 => 
        \U50_PATTERNS/ELINK_DOUTA_12[6]\, DOUTA5 => 
        \U50_PATTERNS/ELINK_DOUTA_12[5]\, DOUTA4 => 
        \U50_PATTERNS/ELINK_DOUTA_12[4]\, DOUTA3 => 
        \U50_PATTERNS/ELINK_DOUTA_12[3]\, DOUTA2 => 
        \U50_PATTERNS/ELINK_DOUTA_12[2]\, DOUTA1 => 
        \U50_PATTERNS/ELINK_DOUTA_12[1]\, DOUTA0 => 
        \U50_PATTERNS/ELINK_DOUTA_12[0]\, DOUTB8 => OPEN, DOUTB7
         => \PATT_ELK_DAT_12[7]\, DOUTB6 => \PATT_ELK_DAT_12[6]\, 
        DOUTB5 => \PATT_ELK_DAT_12[5]\, DOUTB4 => 
        \PATT_ELK_DAT_12[4]\, DOUTB3 => \PATT_ELK_DAT_12[3]\, 
        DOUTB2 => \PATT_ELK_DAT_12[2]\, DOUTB1 => 
        \PATT_ELK_DAT_12[1]\, DOUTB0 => \PATT_ELK_DAT_12[0]\);
    
    \U50_PATTERNS/ELINK_ADDRA_8[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119945, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_8, Q => 
        \U50_PATTERNS/ELINK_ADDRA_8[6]\);
    
    HIEFFPLA_INST_0_54285 : MX2
      port map(A => HIEFFPLA_NET_0_116207, B => 
        HIEFFPLA_NET_0_116097, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_2[3]_net_1\, Y
         => HIEFFPLA_NET_0_117285);
    
    HIEFFPLA_INST_0_50971 : MX2
      port map(A => \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\, B
         => \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[13]_net_1\, S => 
        \BIT_OS_SEL_4[2]\, Y => HIEFFPLA_NET_0_117855);
    
    AFLSDF_INV_16 : INV
      port map(A => DCB_SALT_SEL_c, Y => \AFLSDF_INV_16\);
    
    HIEFFPLA_INST_0_47160 : MX2
      port map(A => \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\, 
        B => \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\, S => 
        \BIT_OS_SEL_3[2]\, Y => HIEFFPLA_NET_0_118541);
    
    \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117717, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_31, Q => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[2]_net_1\);
    
    HIEFFPLA_INST_0_57135 : XA1B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_2[2]\, B => 
        HIEFFPLA_NET_0_116738, C => HIEFFPLA_NET_0_117179, Y => 
        HIEFFPLA_NET_0_116733);
    
    HIEFFPLA_INST_0_56789 : XA1C
      port map(A => HIEFFPLA_NET_0_116809, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_0[4]\, C => 
        HIEFFPLA_NET_0_117179, Y => HIEFFPLA_NET_0_116796);
    
    HIEFFPLA_INST_0_52246 : AO1
      port map(A => HIEFFPLA_NET_0_117589, B => 
        HIEFFPLA_NET_0_117597, C => HIEFFPLA_NET_0_117179, Y => 
        HIEFFPLA_NET_0_117601);
    
    HIEFFPLA_INST_0_44296 : MX2
      port map(A => \TFC_STRT_ADDR[7]\, B => 
        \U50_PATTERNS/U4A_REGCROSS/SAMP_TWO[7]_net_1\, S => 
        HIEFFPLA_NET_0_119156, Y => HIEFFPLA_NET_0_119147);
    
    \U50_PATTERNS/ELINK_ADDRA_18[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120022, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_12, Q => 
        \U50_PATTERNS/ELINK_ADDRA_18[1]\);
    
    HIEFFPLA_INST_0_50607 : AND2A
      port map(A => \OP_MODE_c_4[1]\, B => \PATT_ELK_DAT_7[0]\, Y
         => HIEFFPLA_NET_0_117923);
    
    HIEFFPLA_INST_0_112589 : AO18
      port map(A => HIEFFPLA_NET_0_115814, B => 
        HIEFFPLA_NET_0_116978, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_SEQCNT[3]\, Y => 
        HIEFFPLA_NET_0_115835);
    
    HIEFFPLA_INST_0_39191 : MX2
      port map(A => HIEFFPLA_NET_0_119518, B => 
        \U50_PATTERNS/ELINK_ADDRA_18[5]\, S => 
        HIEFFPLA_NET_0_119264, Y => HIEFFPLA_NET_0_120018);
    
    \U50_PATTERNS/TFC_STRT_ADDR[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119165, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_13, Q => 
        \U50_PATTERNS/TFC_STRT_ADDR[7]\);
    
    \U50_PATTERNS/ELINK_ADDRA_15[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120040, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_6, Q => 
        \U50_PATTERNS/ELINK_ADDRA_15[7]\);
    
    \U_ELK16_CH/U_SLAVE_1ELK/RECD_SER_WORD[3]\ : DFN1C0
      port map(D => \U_ELK16_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[3]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_16[3]\);
    
    \U_ELK5_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]\ : DFN1C0
      port map(D => \U_ELK5_CH/U_SLAVE_1ELK/Q[5]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]_net_1\);
    
    HIEFFPLA_INST_0_45935 : AND3A
      port map(A => HIEFFPLA_NET_0_119376, B => 
        \U50_PATTERNS/TFC_STRT_ADDR[5]\, C => 
        HIEFFPLA_NET_0_119431, Y => HIEFFPLA_NET_0_118807);
    
    HIEFFPLA_INST_0_61526 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_7[2]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_23[2]\, S
         => \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[4]_net_1\, 
        Y => HIEFFPLA_NET_0_116115);
    
    \U_ELK1_CH/U_ELK1_SERDAT_SOURCE/SERDAT[7]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118186, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_11, Q => 
        \U_ELK1_CH/ELK_TX_DAT[7]\);
    
    AFLSDF_INV_25 : INV
      port map(A => DCB_SALT_SEL_c, Y => \AFLSDF_INV_25\);
    
    \U_ELK7_CH/U_SLAVE_1ELK/RECD_SER_WORD[3]\ : DFN1C0
      port map(D => \U_ELK7_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[3]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_7[3]\);
    
    \U_TFC_SERDAT_SOURCE/SERDAT[3]\ : DFN1C0
      port map(D => \U_TFC_SERDAT_SOURCE/N_SERDAT[3]\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \TFC_TX_DAT[3]\);
    
    HIEFFPLA_INST_0_45411 : NAND2A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_4[5]\, Y => 
        HIEFFPLA_NET_0_118918);
    
    \U_EXEC_MASTER/MPOR_SALT_B_14\ : DFI1P0
      port map(D => HIEFFPLA_NET_0_117781, CLK => CLK_40M_GL, PRE
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_2\, QN => 
        MASTER_SALT_POR_B_i_0_i_14);
    
    \U_ELK8_CH/U_ELK1_SERDAT_SOURCE/SERDAT[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117875, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_5, Q => 
        \U_ELK8_CH/ELK_TX_DAT[3]\);
    
    HIEFFPLA_INST_0_46210 : AO1
      port map(A => HIEFFPLA_NET_0_119246, B => 
        \U50_PATTERNS/ELINK_DOUTA_3[2]\, C => 
        HIEFFPLA_NET_0_118911, Y => HIEFFPLA_NET_0_118742);
    
    \U_ELK2_CH/U_SLAVE_1ELK/Q[4]\ : DFN1C0
      port map(D => \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/Q[4]_net_1\);
    
    HIEFFPLA_INST_0_57960 : NAND2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_7[3]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_7[2]\, Y => 
        HIEFFPLA_NET_0_116591);
    
    HIEFFPLA_INST_0_44686 : MX2
      port map(A => \OP_MODE[4]\, B => 
        \U50_PATTERNS/U4E_REGCROSS/SAMP_TWO[4]_net_1\, S => 
        HIEFFPLA_NET_0_119072, Y => HIEFFPLA_NET_0_119066);
    
    HIEFFPLA_INST_0_38102 : AND2B
      port map(A => \U200B_ELINKS/GP_PG_SM[10]_net_1\, B => 
        \U200B_ELINKS/GP_PG_SM[1]_net_1\, Y => 
        HIEFFPLA_NET_0_120152);
    
    \U_ELK9_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2\ : IOPADN_BI
      port map(DB => \U_ELK9_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, 
        E => \U_ELK9_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET3\, PAD => 
        ELK9_DAT_N, N2POUT => 
        \U_ELK9_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2_N2P\);
    
    \U50_PATTERNS/ELINK_DINA_5[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119748, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_14, Q => 
        \U50_PATTERNS/ELINK_DINA_5[3]\);
    
    HIEFFPLA_INST_0_57297 : AOI1A
      port map(A => HIEFFPLA_NET_0_116713, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_3[0]\, C => 
        HIEFFPLA_NET_0_116704, Y => HIEFFPLA_NET_0_116705);
    
    \U50_PATTERNS/U4A_REGCROSS/LOCAL_REG_VAL[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119149, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_17, Q => \TFC_STRT_ADDR[5]\);
    
    HIEFFPLA_INST_0_55721 : AO1
      port map(A => HIEFFPLA_NET_0_117087, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_3[0]\, C => 
        HIEFFPLA_NET_0_116997, Y => HIEFFPLA_NET_0_116999);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_30[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116027, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_8, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_30[3]\);
    
    \U_ELK9_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U3\ : IOBI_ID_OD_EB
      port map(DR => \U_ELK9_CH/ELK_OUT_R\, DF => 
        \U_ELK9_CH/ELK_OUT_F\, CLR => \GND\, E => \AFLSDF_INV_51\, 
        ICLK => CCC_160M_ADJ, OCLK => CCC_160M_FXD, YIN => 
        \U_ELK9_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\, DOUT => OPEN, 
        EOUT => \U_ELK9_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET3\, YR
         => OPEN, YF => OPEN);
    
    HIEFFPLA_INST_0_111798 : XA1A
      port map(A => HIEFFPLA_NET_0_115831, B => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[4]\, C => 
        HIEFFPLA_NET_0_117674, Y => HIEFFPLA_NET_0_117678);
    
    HIEFFPLA_INST_0_55936 : NAND3A
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[1]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[2]\, C
         => \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[4]\, Y => 
        HIEFFPLA_NET_0_116971);
    
    HIEFFPLA_INST_0_47407 : MX2
      port map(A => \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\, 
        B => \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\, S => 
        \BIT_OS_SEL_3[2]\, Y => HIEFFPLA_NET_0_118496);
    
    HIEFFPLA_INST_0_37240 : AO1
      port map(A => HIEFFPLA_NET_0_120326, B => 
        HIEFFPLA_NET_0_120306, C => HIEFFPLA_NET_0_120298, Y => 
        HIEFFPLA_NET_0_120317);
    
    \U_ELK5_CH/U_SLAVE_1ELK/Q[14]\ : DFN1C0
      port map(D => \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[14]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/Q[14]_net_1\);
    
    HIEFFPLA_INST_0_63161 : AX1C
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[0]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[1]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[2]\, Y => 
        HIEFFPLA_NET_0_115871);
    
    HIEFFPLA_INST_0_60510 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_11[4]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_12[4]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_4[0]\, Y => 
        HIEFFPLA_NET_0_116256);
    
    HIEFFPLA_INST_0_40432 : MX2
      port map(A => HIEFFPLA_NET_0_119566, B => 
        \U50_PATTERNS/ELINK_DINA_11[6]\, S => 
        HIEFFPLA_NET_0_119280, Y => HIEFFPLA_NET_0_119849);
    
    \U_ELK5_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]\ : DFN1C0
      port map(D => \U_ELK5_CH/U_SLAVE_1ELK/Q[11]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]_net_1\);
    
    HIEFFPLA_INST_0_44433 : XOR2
      port map(A => \TFC_STOP_ADDR[3]\, B => 
        \U50_PATTERNS/U4B_REGCROSS/SAMP_TWO[3]_net_1\, Y => 
        HIEFFPLA_NET_0_119119);
    
    HIEFFPLA_INST_0_42019 : AO1
      port map(A => HIEFFPLA_NET_0_119552, B => 
        HIEFFPLA_NET_0_119555, C => 
        \U50_PATTERNS/ELK_N_ACTIVE_net_1\, Y => 
        HIEFFPLA_NET_0_119630);
    
    \U_ELK10_CH/U_SLAVE_1ELK/Q[11]\ : DFN1C0
      port map(D => \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/Q[11]_net_1\);
    
    \U_ELK17_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2\ : IOPADN_BI
      port map(DB => \U_ELK17_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, 
        E => \U_ELK17_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET3\, PAD
         => ELK17_DAT_N, N2POUT => 
        \U_ELK17_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2_N2P\);
    
    \U_ELK10_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]\ : DFN1C0
      port map(D => \U_ELK10_CH/U_SLAVE_1ELK/Q[2]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]_net_1\);
    
    HIEFFPLA_INST_0_57817 : AND3B
      port map(A => HIEFFPLA_NET_0_117179, B => 
        HIEFFPLA_NET_0_116606, C => HIEFFPLA_NET_0_116623, Y => 
        HIEFFPLA_NET_0_116614);
    
    \U50_PATTERNS/ELINK_DINA_10[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119857, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_9, Q => 
        \U50_PATTERNS/ELINK_DINA_10[6]\);
    
    HIEFFPLA_INST_0_47718 : MX2
      port map(A => HIEFFPLA_NET_0_118445, B => 
        HIEFFPLA_NET_0_118441, S => \BIT_OS_SEL_2[1]\, Y => 
        HIEFFPLA_NET_0_118442);
    
    HIEFFPLA_INST_0_58091 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_0[2]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_16[2]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_1[4]_net_1\, Y
         => HIEFFPLA_NET_0_116565);
    
    \U50_PATTERNS/ELINK_DINA_14[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119826, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_16, Q => 
        \U50_PATTERNS/ELINK_DINA_14[5]\);
    
    HIEFFPLA_INST_0_53584 : AND3A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[0]_net_1\, B
         => \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[2]_net_1\, C
         => \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[1]_net_1\, 
        Y => HIEFFPLA_NET_0_117386);
    
    \U50_PATTERNS/ELINK_ADDRA_9[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119942, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_10, Q => 
        \U50_PATTERNS/ELINK_ADDRA_9[1]\);
    
    \U200A_TFC/RX_SER_WORD_3DEL[0]\ : DFN1C0
      port map(D => \U200A_TFC/RX_SER_WORD_2DEL[0]_net_1\, CLK
         => CLK_40M_GL, CLR => P_MASTER_POR_B_c_24, Q => 
        \U200A_TFC/RX_SER_WORD_3DEL[0]_net_1\);
    
    \U_ELK14_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL\ : DFN1C0
      port map(D => 
        \U_ELK14_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL_net_1\);
    
    \U_ELK10_CH/U_ELK1_SERDAT_SOURCE/SERDAT[7]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118636, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_17, Q => 
        \U_ELK10_CH/ELK_TX_DAT[7]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/ALIGN_ACTIVE/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117609, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_9, Q => ALIGN_ACTIVE);
    
    HIEFFPLA_INST_0_40351 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_10[5]\, B => 
        HIEFFPLA_NET_0_119567, S => HIEFFPLA_NET_0_119239, Y => 
        HIEFFPLA_NET_0_119858);
    
    \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[6]\ : DFN1C0
      port map(D => \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\);
    
    \U_ELK5_CH/U_SLAVE_1ELK/Q[9]\ : DFN1C0
      port map(D => \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/Q[9]_net_1\);
    
    HIEFFPLA_INST_0_55181 : NAND2B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[8]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[0]_net_1\, Y => 
        HIEFFPLA_NET_0_117102);
    
    HIEFFPLA_INST_0_50565 : MX2
      port map(A => \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\, 
        B => \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[14]_net_1\, S => 
        \BIT_OS_SEL_7[2]\, Y => HIEFFPLA_NET_0_117933);
    
    HIEFFPLA_INST_0_38858 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_14[0]\, B => 
        HIEFFPLA_NET_0_119524, S => HIEFFPLA_NET_0_119249, Y => 
        HIEFFPLA_NET_0_120055);
    
    \U50_PATTERNS/WR_USB_ADBUS[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118983, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_15, Q => 
        \U50_PATTERNS/WR_USB_ADBUS[2]\);
    
    HIEFFPLA_INST_0_42864 : NAND3B
      port map(A => \U50_PATTERNS/REG_STATE[3]_net_1\, B => 
        HIEFFPLA_NET_0_119435, C => 
        \U50_PATTERNS/REG_STATE[0]_net_1\, Y => 
        HIEFFPLA_NET_0_119444);
    
    HIEFFPLA_INST_0_57683 : XA1C
      port map(A => HIEFFPLA_NET_0_116651, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_5[8]\, C => 
        HIEFFPLA_NET_0_117179, Y => HIEFFPLA_NET_0_116636);
    
    HIEFFPLA_INST_0_54349 : MX2
      port map(A => HIEFFPLA_NET_0_116155, B => 
        HIEFFPLA_NET_0_116047, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_2[3]_net_1\, Y
         => HIEFFPLA_NET_0_117277);
    
    HIEFFPLA_INST_0_47230 : MX2
      port map(A => \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[1]_net_1\, 
        B => \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\, S => 
        \BIT_OS_SEL_3[2]\, Y => HIEFFPLA_NET_0_118531);
    
    \U_ELK4_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]\ : DFN1C0
      port map(D => \U_ELK4_CH/U_SLAVE_1ELK/Q[8]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]_net_1\);
    
    HIEFFPLA_INST_0_61034 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_2[4]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_18[4]\, S
         => \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_4[4]_net_1\, 
        Y => HIEFFPLA_NET_0_116182);
    
    HIEFFPLA_INST_0_52146 : AOI1D
      port map(A => HIEFFPLA_NET_0_117683, B => 
        HIEFFPLA_NET_0_117688, C => 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM[0]_net_1\, Y => 
        HIEFFPLA_NET_0_117625);
    
    HIEFFPLA_INST_0_46035 : AND3
      port map(A => \U50_PATTERNS/TFC_DOUTA[0]\, B => 
        HIEFFPLA_NET_0_118997, C => HIEFFPLA_NET_0_119365, Y => 
        HIEFFPLA_NET_0_118781);
    
    HIEFFPLA_INST_0_41947 : AO1A
      port map(A => \U50_PATTERNS/SM_BANK_SEL[8]\, B => 
        HIEFFPLA_NET_0_119240, C => \U50_PATTERNS/ELINK_RWA[19]\, 
        Y => HIEFFPLA_NET_0_119650);
    
    HIEFFPLA_INST_0_52686 : MX2
      port map(A => HIEFFPLA_NET_0_117479, B => 
        HIEFFPLA_NET_0_117475, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[4]\, Y => 
        HIEFFPLA_NET_0_117527);
    
    \U_ELK6_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117973, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_6, Q => 
        \U_ELK6_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]_net_1\);
    
    \U_ELK3_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]\ : DFN1C0
      port map(D => \U_ELK3_CH/U_SLAVE_1ELK/Q[8]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]_net_1\);
    
    HIEFFPLA_INST_0_57835 : XA1C
      port map(A => HIEFFPLA_NET_0_116622, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_6[5]\, C => 
        HIEFFPLA_NET_0_117179, Y => HIEFFPLA_NET_0_116610);
    
    HIEFFPLA_INST_0_40138 : AOI1C
      port map(A => \U50_PATTERNS/ELINK_BLKA[2]\, B => 
        HIEFFPLA_NET_0_119646, C => HIEFFPLA_NET_0_119893, Y => 
        HIEFFPLA_NET_0_119894);
    
    HIEFFPLA_INST_0_111665 : AOI1B
      port map(A => HIEFFPLA_NET_0_115833, B => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[0]\, C => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[5]\, Y => 
        HIEFFPLA_NET_0_117667);
    
    HIEFFPLA_INST_0_49071 : MX2
      port map(A => \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\, 
        B => \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[14]_net_1\, S => 
        \BIT_OS_SEL_1[2]\, Y => HIEFFPLA_NET_0_118203);
    
    \U_ELK17_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL\ : DFN1C0
      port map(D => \U_ELK17_CH/ELK_IN_R_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL_net_1\);
    
    \U_ELK7_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]\ : DFN1C0
      port map(D => \U_ELK7_CH/U_SLAVE_1ELK/Q[6]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]_net_1\);
    
    \U_ELK16_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]\ : DFN1C0
      port map(D => \U_ELK16_CH/U_SLAVE_1ELK/Q[0]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]_net_1\);
    
    \U50_PATTERNS/TFC_ADDRA[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119200, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_10, Q => 
        \U50_PATTERNS/TFC_ADDRA[7]\);
    
    HIEFFPLA_INST_0_48327 : AND2
      port map(A => \U_ELK17_CH/ELK_TX_DAT[0]\, B => 
        \U_ELK17_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118337);
    
    \U_ELK16_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]\ : DFN1C0
      port map(D => \U_ELK16_CH/U_SLAVE_1ELK/Q[4]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]_net_1\);
    
    \U50_PATTERNS/ELINK_DINA_0[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119866, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_5, Q => 
        \U50_PATTERNS/ELINK_DINA_0[5]\);
    
    \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[10]\ : DFN1C0
      port map(D => \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\);
    
    \U_ELK17_CH/U_SLAVE_1ELK/Q[13]\ : DFN1C0
      port map(D => \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[13]_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/Q[13]_net_1\);
    
    HIEFFPLA_INST_0_57479 : NAND3C
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_4[4]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_4[8]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_4[5]\, Y => 
        HIEFFPLA_NET_0_116674);
    
    HIEFFPLA_INST_0_45548 : AO1A
      port map(A => HIEFFPLA_NET_0_119475, B => 
        \U50_PATTERNS/ELINKS_STOP_ADDR[5]\, C => 
        HIEFFPLA_NET_0_118807, Y => HIEFFPLA_NET_0_118892);
    
    HIEFFPLA_INST_0_37637 : AND3B
      port map(A => \U200B_ELINKS/LOC_STRT_ADDR[1]\, B => 
        HIEFFPLA_NET_0_120190, C => HIEFFPLA_NET_0_120234, Y => 
        HIEFFPLA_NET_0_120242);
    
    HIEFFPLA_INST_0_49844 : MX2
      port map(A => 
        \U_ELK4_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]_net_1\, B => 
        \U_ELK4_CH/ELK_TX_DAT[3]\, S => 
        \U_ELK4_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118062);
    
    \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_SEL_6[1]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_BIT_OS_VAL[1]\, CLK
         => CLK_40M_GL, CLR => P_MASTER_POR_B_c_27_0, Q => 
        \BIT_OS_SEL_6[1]\);
    
    \U_ELK11_CH/U_ELK1_CMD_TX/START_RISE\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118599, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_10, Q => 
        \U_ELK11_CH/U_ELK1_CMD_TX/START_RISE_net_1\);
    
    \U50_PATTERNS/U4E_REGCROSS/SAMP_TWO[6]\ : DFN1C0
      port map(D => \U50_PATTERNS/U4E_REGCROSS/SAMP_ONE[6]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_24, Q => 
        \U50_PATTERNS/U4E_REGCROSS/SAMP_TWO[6]_net_1\);
    
    HIEFFPLA_INST_0_40576 : MX2
      port map(A => HIEFFPLA_NET_0_119566, B => 
        \U50_PATTERNS/ELINK_DINA_13[6]\, S => 
        HIEFFPLA_NET_0_119285, Y => HIEFFPLA_NET_0_119833);
    
    \U_ELK6_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL\ : DFN1C0
      port map(D => \U_ELK6_CH/ELK_IN_R_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL_net_1\);
    
    \U50_PATTERNS/ELINK_BLKA[8]/U1\ : DFN1P0
      port map(D => HIEFFPLA_NET_0_119917, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_19, Q => 
        \U50_PATTERNS/ELINK_BLKA[8]\);
    
    \U_ELK1_CH/U_SLAVE_1ELK/Q[13]\ : DFN1C0
      port map(D => \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[13]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/Q[13]_net_1\);
    
    HIEFFPLA_INST_0_61829 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_10[3]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_26[3]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_4[4]_net_1\, Y
         => HIEFFPLA_NET_0_116072);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_7[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116300, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_3, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_7[3]\);
    
    HIEFFPLA_INST_0_47335 : MX2
      port map(A => 
        \U_ELK13_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]_net_1\, B => 
        \U_ELK13_CH/ELK_TX_DAT[2]\, S => 
        \U_ELK13_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118516);
    
    HIEFFPLA_INST_0_45765 : AO1
      port map(A => HIEFFPLA_NET_0_119288, B => 
        \U50_PATTERNS/ELINK_DOUTA_16[4]\, C => 
        HIEFFPLA_NET_0_118767, Y => HIEFFPLA_NET_0_118849);
    
    \U_ELK19_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL\ : DFN1C0
      port map(D => 
        \U_ELK19_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL_net_1\);
    
    HIEFFPLA_INST_0_48350 : MX2
      port map(A => 
        \U_ELK17_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]_net_1\, B => 
        \U_ELK17_CH/ELK_TX_DAT[3]\, S => 
        \U_ELK17_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118332);
    
    HIEFFPLA_INST_0_54566 : NAND2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[4]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[2]_net_1\, Y => 
        HIEFFPLA_NET_0_117247);
    
    HIEFFPLA_INST_0_52848 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_15[3]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_16[3]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_2[0]\, Y => 
        HIEFFPLA_NET_0_117501);
    
    TFC_SYNC_DET : DFN1C0
      port map(D => HIEFFPLA_NET_0_116906, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_23, Q => P_TFC_SYNC_DET_c);
    
    HIEFFPLA_INST_0_60342 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_9[3]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_25[3]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[4]_net_1\, Y
         => HIEFFPLA_NET_0_116278);
    
    HIEFFPLA_INST_0_54003 : NAND3C
      port map(A => HIEFFPLA_NET_0_117344, B => 
        HIEFFPLA_NET_0_117067, C => HIEFFPLA_NET_0_117389, Y => 
        HIEFFPLA_NET_0_117321);
    
    \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[10]\ : DFN1C0
      port map(D => \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\);
    
    \U_ELK5_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118020, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_6, Q => 
        \U_ELK5_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]_net_1\);
    
    \U_ELK1_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]\ : DFN1C0
      port map(D => \U_ELK1_CH/U_SLAVE_1ELK/Q[10]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]_net_1\);
    
    HIEFFPLA_INST_0_55045 : AO1A
      port map(A => HIEFFPLA_NET_0_117204, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[6]_net_1\, C => 
        HIEFFPLA_NET_0_117182, Y => HIEFFPLA_NET_0_117134);
    
    HIEFFPLA_INST_0_49864 : AND2A
      port map(A => \OP_MODE_c_1[1]\, B => \PATT_ELK_DAT_4[4]\, Y
         => HIEFFPLA_NET_0_118054);
    
    HIEFFPLA_INST_0_38984 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_15[6]\, B => 
        HIEFFPLA_NET_0_119517, S => HIEFFPLA_NET_0_119297, Y => 
        HIEFFPLA_NET_0_120041);
    
    HIEFFPLA_INST_0_60411 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_9[0]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_10[0]\, S
         => \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_1[0]\, Y
         => HIEFFPLA_NET_0_116270);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_1[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116475, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_17, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_1[0]\);
    
    \U50_PATTERNS/OP_MODE_T[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119604, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_17, Q => 
        \U50_PATTERNS/OP_MODE_T[5]\);
    
    \U_ELK2_CH/U_SLAVE_1ELK/Q[10]\ : DFN1C0
      port map(D => \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/Q[10]_net_1\);
    
    HIEFFPLA_INST_0_55778 : MX2
      port map(A => HIEFFPLA_NET_0_116148, B => 
        HIEFFPLA_NET_0_116062, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[3]\, Y => 
        HIEFFPLA_NET_0_116991);
    
    \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM[4]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117622, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_22, Q => 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM[4]_net_1\);
    
    \U_ELK11_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U3\ : IOBI_ID_OD_EB
      port map(DR => \U_ELK11_CH/ELK_OUT_R\, DF => 
        \U_ELK11_CH/ELK_OUT_F\, CLR => \GND\, E => 
        \AFLSDF_INV_17\, ICLK => CCC_160M_ADJ, OCLK => 
        CCC_160M_FXD, YIN => 
        \U_ELK11_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\, DOUT => 
        OPEN, EOUT => 
        \U_ELK11_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET3\, YR => OPEN, 
        YF => OPEN);
    
    HIEFFPLA_INST_0_41807 : MX2
      port map(A => HIEFFPLA_NET_0_119667, B => 
        \U50_PATTERNS/ELINK_RWA[9]\, S => 
        \U50_PATTERNS/SM_BANK_SEL_0[20]\, Y => 
        HIEFFPLA_NET_0_119692);
    
    HIEFFPLA_INST_0_39344 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_1[6]\, B => 
        HIEFFPLA_NET_0_119517, S => HIEFFPLA_NET_0_119243, Y => 
        HIEFFPLA_NET_0_120001);
    
    \U_ELK14_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]\ : DFN1C0
      port map(D => \U_ELK14_CH/U_SLAVE_1ELK/Q[3]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]_net_1\);
    
    \U_ELK13_CH/U_SLAVE_1ELK/Q[3]\ : DFN1C0
      port map(D => \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/Q[3]_net_1\);
    
    HIEFFPLA_INST_0_59162 : AO1A
      port map(A => HIEFFPLA_NET_0_117243, B => 
        HIEFFPLA_NET_0_116649, C => HIEFFPLA_NET_0_116589, Y => 
        HIEFFPLA_NET_0_116426);
    
    HIEFFPLA_INST_0_44762 : MX2B
      port map(A => HIEFFPLA_NET_0_119054, B => 
        HIEFFPLA_NET_0_119072, S => 
        \U50_PATTERNS/U4E_REGCROSS/SYNC_SM[0]_net_1\, Y => 
        HIEFFPLA_NET_0_119055);
    
    \U50_PATTERNS/ELINK_DINA_9[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119712, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_20, Q => 
        \U50_PATTERNS/ELINK_DINA_9[7]\);
    
    HIEFFPLA_INST_0_37276 : NAND3
      port map(A => HIEFFPLA_NET_0_120293, B => 
        \U200A_TFC/GP_PG_SM[2]_net_1\, C => \OP_MODE_c[2]\, Y => 
        HIEFFPLA_NET_0_120309);
    
    \U_EXEC_MASTER/MPOR_B_24\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117787, CLK => CLK_40M_GL, CLR
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_0\, Q => 
        P_MASTER_POR_B_c_24);
    
    \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[12]\ : DFN1C0
      port map(D => \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_2[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116033, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_10, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_2[2]\);
    
    \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_2S_15\ : DFN1C0
      port map(D => 
        \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_1S_0_net_1\, CLK
         => CLK60MHZ, CLR => \U_EXEC_MASTER/P_MASTER_POR_B_c_0\, 
        Q => P_USB_MASTER_EN_c_15);
    
    \U50_PATTERNS/ELINK_RWA[2]/U1\ : DFN1P0
      port map(D => HIEFFPLA_NET_0_119699, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_6, Q => \U50_PATTERNS/ELINK_RWA[2]\);
    
    \U_ELK7_CH/U_SLAVE_1ELK/Q[2]\ : DFN1C0
      port map(D => \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/Q[2]_net_1\);
    
    HIEFFPLA_INST_0_111911 : XA1B
      port map(A => \U50_PATTERNS/WR_XFER_TYPE[1]_net_1\, B => 
        \U50_PATTERNS/WR_XFER_TYPE[0]_net_1\, C => 
        HIEFFPLA_NET_0_118692, Y => HIEFFPLA_NET_0_115823);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_26[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116077, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_12, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_26[3]\);
    
    HIEFFPLA_INST_0_59376 : AO1C
      port map(A => HIEFFPLA_NET_0_117337, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_26[2]\, C => 
        HIEFFPLA_NET_0_117404, Y => HIEFFPLA_NET_0_116400);
    
    HIEFFPLA_INST_0_40603 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_14[1]\, B => 
        HIEFFPLA_NET_0_119576, S => HIEFFPLA_NET_0_119249, Y => 
        HIEFFPLA_NET_0_119830);
    
    \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[5]\ : DFN1C0
      port map(D => \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\);
    
    HIEFFPLA_INST_0_53864 : AND3A
      port map(A => HIEFFPLA_NET_0_117325, B => 
        HIEFFPLA_NET_0_116686, C => HIEFFPLA_NET_0_117334, Y => 
        HIEFFPLA_NET_0_117340);
    
    HIEFFPLA_INST_0_44548 : AND2A
      port map(A => \U50_PATTERNS/U4D_REGCROSS/DELCNT[0]_net_1\, 
        B => \U50_PATTERNS/U4D_REGCROSS/SYNC_SM[0]_net_1\, Y => 
        HIEFFPLA_NET_0_119092);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_12[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116546, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_10, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_12[2]\);
    
    HIEFFPLA_INST_0_56586 : AND3
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[12]_net_1\, B
         => HIEFFPLA_NET_0_117426, C => HIEFFPLA_NET_0_117425, Y
         => HIEFFPLA_NET_0_116833);
    
    \U_ELK9_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]\ : DFN1C0
      port map(D => \U_ELK9_CH/U_SLAVE_1ELK/Q[13]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]_net_1\);
    
    HIEFFPLA_INST_0_52287 : AND3A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[6]_net_1\, B => 
        HIEFFPLA_NET_0_117605, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[4]_net_1\, Y => 
        HIEFFPLA_NET_0_117590);
    
    HIEFFPLA_INST_0_53110 : MX2
      port map(A => HIEFFPLA_NET_0_117548, B => 
        HIEFFPLA_NET_0_117544, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[3]\, Y => 
        HIEFFPLA_NET_0_117464);
    
    HIEFFPLA_INST_0_55033 : AO1C
      port map(A => HIEFFPLA_NET_0_117396, B => 
        HIEFFPLA_NET_0_117164, C => HIEFFPLA_NET_0_117180, Y => 
        HIEFFPLA_NET_0_117137);
    
    HIEFFPLA_INST_0_42525 : NAND3A
      port map(A => HIEFFPLA_NET_0_119514, B => 
        \U50_PATTERNS/REG_ADDR[4]\, C => 
        \U50_PATTERNS/REG_ADDR[3]\, Y => HIEFFPLA_NET_0_119521);
    
    \U50_PATTERNS/SM_BANK_SEL[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119306, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_7, Q => 
        \U50_PATTERNS/SM_BANK_SEL[4]\);
    
    HIEFFPLA_INST_0_54985 : AO1C
      port map(A => HIEFFPLA_NET_0_117202, B => 
        HIEFFPLA_NET_0_117164, C => HIEFFPLA_NET_0_117180, Y => 
        HIEFFPLA_NET_0_117148);
    
    \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[6]\ : DFN1C0
      port map(D => 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\);
    
    \U_ELK10_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL\ : DFN1C0
      port map(D => \U_ELK10_CH/ELK_IN_F_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL_net_1\);
    
    \U_TFC_CMD_TX/SER_CMD_WORD_R[0]\ : DFN1C0
      port map(D => \U_TFC_CMD_TX/N_SER_CMD_WORD_R[0]\, CLK => 
        CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_TFC_CMD_TX/SER_CMD_WORD_R[0]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/Q[9]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[9]_net_1\, CLK => 
        CCC_160M_FXD, CLR => P_MASTER_POR_B_c_34, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/Q[9]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_8[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_115970, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_19, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_8[0]\);
    
    HIEFFPLA_INST_0_57313 : XA1C
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_3[6]\, B => 
        HIEFFPLA_NET_0_116712, C => HIEFFPLA_NET_0_117179, Y => 
        HIEFFPLA_NET_0_116701);
    
    HIEFFPLA_INST_0_57114 : NAND3C
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_2[5]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_2[4]\, C => 
        HIEFFPLA_NET_0_116741, Y => HIEFFPLA_NET_0_116739);
    
    \U_EXEC_MASTER/MPOR_SALT_B_1\ : DFI1P0
      port map(D => HIEFFPLA_NET_0_117781, CLK => CLK_40M_GL, PRE
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i\, QN => 
        MASTER_SALT_POR_B_i_0_i_1);
    
    HIEFFPLA_INST_0_62787 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/TUNE_CLKPHASE[2]\, B => 
        HIEFFPLA_NET_0_115956, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[1]_net_1\, Y => 
        HIEFFPLA_NET_0_115947);
    
    \U50_PATTERNS/SM_BANK_SEL[20]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119310, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_1_0, Q => 
        \U50_PATTERNS/SM_BANK_SEL[20]\);
    
    HIEFFPLA_INST_0_62191 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_14[4]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_30[4]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[4]_net_1\, Y => 
        HIEFFPLA_NET_0_116025);
    
    HIEFFPLA_INST_0_44913 : AND3C
      port map(A => \U50_PATTERNS/REG_STATE[1]_net_1\, B => 
        \U50_PATTERNS/REG_STATE[0]_net_1\, C => 
        \U50_PATTERNS/USB_RXF_B\, Y => HIEFFPLA_NET_0_119022);
    
    HIEFFPLA_INST_0_53417 : AND2
      port map(A => HIEFFPLA_NET_0_116649, B => 
        HIEFFPLA_NET_0_117337, Y => HIEFFPLA_NET_0_117411);
    
    HIEFFPLA_INST_0_42916 : NOR3A
      port map(A => HIEFFPLA_NET_0_119328, B => 
        HIEFFPLA_NET_0_119380, C => 
        \U50_PATTERNS/REG_STATE[3]_net_1\, Y => 
        HIEFFPLA_NET_0_119425);
    
    \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[9]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_WRD_40M_FIXED[9]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_27_1, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[9]_net_1\);
    
    \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[4]\ : DFN1C0
      port map(D => 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\);
    
    \U_ELK3_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118106, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_12, Q => 
        \U_ELK3_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]_net_1\);
    
    \U_ELK2_CH/U_SLAVE_1ELK/Q[1]\ : DFN1C0
      port map(D => \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/Q[1]_net_1\);
    
    \U50_PATTERNS/ELINK_ADDRA_7[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119959, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_5, Q => 
        \U50_PATTERNS/ELINK_ADDRA_7[0]\);
    
    \P_CCC_160M_FXD_pad/U0/U0\ : IOPAD_TRI_U
      port map(D => \P_CCC_160M_FXD_pad/U0/NET1\, E => 
        \P_CCC_160M_FXD_pad/U0/NET2\, PAD => P_CCC_160M_FXD);
    
    HIEFFPLA_INST_0_46194 : NAND3C
      port map(A => HIEFFPLA_NET_0_118913, B => 
        HIEFFPLA_NET_0_118916, C => HIEFFPLA_NET_0_118922, Y => 
        HIEFFPLA_NET_0_118745);
    
    HIEFFPLA_INST_0_48595 : AND2
      port map(A => \U_ELK18_CH/ELK_TX_DAT[1]\, B => 
        \U_ELK18_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118288);
    
    HIEFFPLA_INST_0_43587 : AND2A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/SM_BANK_SEL[8]\, Y => HIEFFPLA_NET_0_119277);
    
    HIEFFPLA_INST_0_56755 : NAND2B
      port map(A => HIEFFPLA_NET_0_116774, B => 
        HIEFFPLA_NET_0_116813, Y => HIEFFPLA_NET_0_116806);
    
    \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[9]\ : DFN1C0
      port map(D => \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\);
    
    HIEFFPLA_INST_0_50846 : MX2
      port map(A => 
        \U_ELK8_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]_net_1\, B => 
        \U_ELK8_CH/ELK_TX_DAT[5]\, S => 
        \U_ELK8_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_117881);
    
    HIEFFPLA_INST_0_42542 : AND3B
      port map(A => \U50_PATTERNS/REG_ADDR[1]\, B => 
        \U50_PATTERNS/REG_ADDR[0]\, C => HIEFFPLA_NET_0_119512, Y
         => HIEFFPLA_NET_0_119515);
    
    HIEFFPLA_INST_0_49140 : MX2
      port map(A => HIEFFPLA_NET_0_118180, B => 
        HIEFFPLA_NET_0_118178, S => \BIT_OS_SEL_0[1]\, Y => 
        HIEFFPLA_NET_0_118183);
    
    \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[1]\ : DFN1C0
      port map(D => 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[1]_net_1\);
    
    HIEFFPLA_INST_0_47360 : MX2
      port map(A => 
        \U_ELK13_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]_net_1\, B => 
        \U_ELK13_CH/ELK_TX_DAT[5]\, S => 
        \U_ELK13_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118511);
    
    \U_ELK3_CH/U_SLAVE_1ELK/RECD_SER_WORD[5]\ : DFN1C0
      port map(D => \U_ELK3_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[5]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_3[5]\);
    
    \U50_PATTERNS/ELINK_RWA[14]/U1\ : DFN1P0
      port map(D => HIEFFPLA_NET_0_119706, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_12, Q => 
        \U50_PATTERNS/ELINK_RWA[14]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[6]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_WRD_40M_FIXED[6]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_27, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[6]_net_1\);
    
    HIEFFPLA_INST_0_42407 : AO1A
      port map(A => HIEFFPLA_NET_0_119019, B => 
        \U50_PATTERNS/RD_USB_ADBUS[5]\, C => 
        HIEFFPLA_NET_0_119536, Y => HIEFFPLA_NET_0_119544);
    
    \U50_PATTERNS/ELINK_DINA_10[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119861, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_9, Q => 
        \U50_PATTERNS/ELINK_DINA_10[2]\);
    
    HIEFFPLA_INST_0_48841 : MX2
      port map(A => 
        \U_ELK19_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]_net_1\, B => 
        \U_ELK19_CH/ELK_TX_DAT[6]\, S => 
        \U_ELK19_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118244);
    
    \U_ELK1_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118197, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_4, Q => 
        \U_ELK1_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]_net_1\);
    
    HIEFFPLA_INST_0_46583 : NAND2B
      port map(A => \OP_MODE_c_4[1]\, B => \PATT_ELK_DAT_0[7]\, Y
         => HIEFFPLA_NET_0_118653);
    
    \U_ELK17_CH/U_ELK1_SERDAT_SOURCE/SERDAT[5]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118323, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_11, Q => 
        \U_ELK17_CH/ELK_TX_DAT[5]\);
    
    \U50_PATTERNS/U4C_REGCROSS/SAMP_ONE[0]\ : DFN1C0
      port map(D => \U50_PATTERNS/ELINKS_STRT_ADDR[0]\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_33, Q => 
        \U50_PATTERNS/U4C_REGCROSS/SAMP_ONE[0]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_SEL_1[2]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_BIT_OS_VAL[2]\, CLK
         => CLK_40M_GL, CLR => P_MASTER_POR_B_c_27_1, Q => 
        \BIT_OS_SEL_1[2]\);
    
    \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[5]\ : DFN1C0
      port map(D => 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\);
    
    HIEFFPLA_INST_0_42968 : AO1
      port map(A => \U50_PATTERNS/REG_STATE[3]_net_1\, B => 
        HIEFFPLA_NET_0_119380, C => HIEFFPLA_NET_0_119022, Y => 
        HIEFFPLA_NET_0_119414);
    
    HIEFFPLA_INST_0_38570 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_10[0]\, B => 
        HIEFFPLA_NET_0_119524, S => HIEFFPLA_NET_0_119239, Y => 
        HIEFFPLA_NET_0_120087);
    
    HIEFFPLA_INST_0_112354 : MX2A
      port map(A => HIEFFPLA_NET_0_115815, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_13[1]\, S => 
        HIEFFPLA_NET_0_117396, Y => HIEFFPLA_NET_0_116536);
    
    \U50_PATTERNS/U4D_REGCROSS/SAMP_TWO[4]\ : DFN1C0
      port map(D => \U50_PATTERNS/U4D_REGCROSS/SAMP_ONE[4]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_30, Q => 
        \U50_PATTERNS/U4D_REGCROSS/SAMP_TWO[4]_net_1\);
    
    \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[12]\ : DFN1C0
      port map(D => 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[12]_net_1\);
    
    HIEFFPLA_INST_0_55246 : XA1C
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[5]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[0]_net_1\, C => 
        HIEFFPLA_NET_0_117102, Y => HIEFFPLA_NET_0_117077);
    
    \U_MASTER_DES/U13C_MASTER_DESER/RECD_SER_WORD[6]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_116898, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_30, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/RECD_SER_WORD[6]_net_1\);
    
    \U_ELK6_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117971, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_6, Q => 
        \U_ELK6_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]_net_1\);
    
    \U50_PATTERNS/U4A_REGCROSS/SAMP_TWO[7]\ : DFN1C0
      port map(D => \U50_PATTERNS/U4A_REGCROSS/SAMP_ONE[7]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_22, Q => 
        \U50_PATTERNS/U4A_REGCROSS/SAMP_TWO[7]_net_1\);
    
    HIEFFPLA_INST_0_49160 : MX2
      port map(A => \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[3]_net_1\, B
         => \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\, S => 
        \BIT_OS_SEL[2]\, Y => HIEFFPLA_NET_0_118180);
    
    HIEFFPLA_INST_0_38732 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_12[2]\, B => 
        HIEFFPLA_NET_0_119522, S => HIEFFPLA_NET_0_119295, Y => 
        HIEFFPLA_NET_0_120069);
    
    \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[2]\ : DFN1C0
      port map(D => \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_7[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_115980, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_17_0, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_7[0]\);
    
    \U_ELK13_CH/U_SLAVE_1ELK/Q[14]\ : DFN1C0
      port map(D => \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[14]_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/Q[14]_net_1\);
    
    HIEFFPLA_INST_0_41969 : AND3C
      port map(A => HIEFFPLA_NET_0_119237, B => 
        HIEFFPLA_NET_0_119270, C => 
        \U50_PATTERNS/SM_BANK_SEL[11]\, Y => 
        HIEFFPLA_NET_0_119642);
    
    HIEFFPLA_INST_0_60756 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_15[3]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_16[3]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[0]\, Y => 
        HIEFFPLA_NET_0_116225);
    
    \U200A_TFC/RX_SER_WORD_3DEL[4]\ : DFN1C0
      port map(D => \U200A_TFC/RX_SER_WORD_2DEL[4]_net_1\, CLK
         => CLK_40M_GL, CLR => P_MASTER_POR_B_c_24, Q => 
        \U200A_TFC/RX_SER_WORD_3DEL[4]_net_1\);
    
    HIEFFPLA_INST_0_42246 : AND3B
      port map(A => \U50_PATTERNS/RD_USB_ADBUS[0]\, B => 
        HIEFFPLA_NET_0_119208, C => 
        \U50_PATTERNS/RD_USB_ADBUS[1]\, Y => 
        HIEFFPLA_NET_0_119592);
    
    HIEFFPLA_INST_0_60624 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_13[2]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_29[2]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_2[4]_net_1\, Y
         => HIEFFPLA_NET_0_116242);
    
    HIEFFPLA_INST_0_38282 : MX2
      port map(A => \U50_PATTERNS/ELINKS_STOP_ADDR[5]\, B => 
        \U50_PATTERNS/ELINKS_STOP_ADDR_T[5]\, S => 
        HIEFFPLA_NET_0_119472, Y => HIEFFPLA_NET_0_120122);
    
    \U_ELK19_CH/U_SLAVE_1ELK/Q[11]\ : DFN1C0
      port map(D => \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/Q[11]_net_1\);
    
    HIEFFPLA_INST_0_43638 : NAND3C
      port map(A => \U50_PATTERNS/SM_BANK_SEL[8]\, B => 
        \U50_PATTERNS/SM_BANK_SEL[0]\, C => HIEFFPLA_NET_0_119269, 
        Y => HIEFFPLA_NET_0_119259);
    
    HIEFFPLA_INST_0_51523 : AO1A
      port map(A => 
        \U_EXEC_MASTER/USB_MASTER_EN/TERMCNT_FG40M2S_net_1\, B
         => \U_EXEC_MASTER/USB_MASTER_EN/TEST_SM[1]_net_1\, C => 
        \U_EXEC_MASTER/USB_MASTER_EN/TEST_SM[3]_net_1\, Y => 
        HIEFFPLA_NET_0_117754);
    
    HIEFFPLA_INST_0_60965 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_1[1]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_17[1]\, S
         => \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_3[4]_net_1\, 
        Y => HIEFFPLA_NET_0_116191);
    
    \U50_PATTERNS/ELINKS_STOP_ADDR_T[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120114, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_7, Q => 
        \U50_PATTERNS/ELINKS_STOP_ADDR_T[5]\);
    
    HIEFFPLA_INST_0_54692 : MX2
      port map(A => HIEFFPLA_NET_0_117376, B => 
        HIEFFPLA_NET_0_117253, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[0]_net_1\, Y => 
        HIEFFPLA_NET_0_117222);
    
    \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[7]\ : DFN1C0
      port map(D => \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\);
    
    HIEFFPLA_INST_0_47057 : MX2
      port map(A => HIEFFPLA_NET_0_118564, B => 
        HIEFFPLA_NET_0_118575, S => \BIT_OS_SEL_4[1]\, Y => 
        HIEFFPLA_NET_0_118566);
    
    HIEFFPLA_INST_0_46092 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_9[2]\, C => 
        \U50_PATTERNS/SM_BANK_SEL[10]\, Y => 
        HIEFFPLA_NET_0_118768);
    
    \U50_PATTERNS/U4B_REGCROSS/DELCNT[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119115, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_30, Q => 
        \U50_PATTERNS/U4B_REGCROSS/DELCNT[1]_net_1\);
    
    HIEFFPLA_INST_0_61178 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_1[2]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_2[2]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_1[0]\, Y => 
        HIEFFPLA_NET_0_116163);
    
    HIEFFPLA_INST_0_58648 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_18[2]\, B => 
        HIEFFPLA_NET_0_116489, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_2[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116493);
    
    HIEFFPLA_INST_0_44337 : XOR2
      port map(A => \TFC_STRT_ADDR[7]\, B => 
        \U50_PATTERNS/U4A_REGCROSS/SAMP_TWO[7]_net_1\, Y => 
        HIEFFPLA_NET_0_119137);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_4[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116326, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_21, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_4[3]\);
    
    HIEFFPLA_INST_0_48128 : MX2
      port map(A => \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[1]_net_1\, 
        B => \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\, S => 
        \BIT_OS_SEL_1[2]\, Y => HIEFFPLA_NET_0_118365);
    
    HIEFFPLA_INST_0_47086 : MX2
      port map(A => 
        \U_ELK12_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]_net_1\, B => 
        \U_ELK12_CH/ELK_TX_DAT[2]\, S => 
        \U_ELK12_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118561);
    
    HIEFFPLA_INST_0_49057 : MX2
      port map(A => HIEFFPLA_NET_0_118218, B => 
        HIEFFPLA_NET_0_118203, S => \BIT_OS_SEL_1[1]\, Y => 
        HIEFFPLA_NET_0_118205);
    
    \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[13]\ : DFN1C0
      port map(D => \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[13]_net_1\);
    
    \U_ELK18_CH/U_ELK1_SERDAT_SOURCE/SERDAT[7]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118276, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_13, Q => 
        \U_ELK18_CH/ELK_TX_DAT[7]\);
    
    HIEFFPLA_INST_0_57241 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_3[7]\, B => 
        HIEFFPLA_NET_0_116700, S => HIEFFPLA_NET_0_117120, Y => 
        HIEFFPLA_NET_0_116718);
    
    HIEFFPLA_INST_0_53316 : AND3A
      port map(A => \BIT_OS_SEL_1[0]\, B => HIEFFPLA_NET_0_117423, 
        C => \BIT_OS_SEL_1[1]\, Y => HIEFFPLA_NET_0_117431);
    
    \U50_PATTERNS/U4E_REGCROSS/LOCAL_REG_VAL[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119067, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_6, Q => 
        \U50_PATTERNS/U4E_REGCROSS/LOCAL_REG_VAL[3]\);
    
    HIEFFPLA_INST_0_51542 : AO1
      port map(A => 
        \U_EXEC_MASTER/USB_MASTER_EN/TEST_SM[3]_net_1\, B => 
        \U_EXEC_MASTER/USB_MASTER_EN/TERMCNT_FG40M2S_net_1\, C
         => \U_EXEC_MASTER/USB_MASTER_EN/TEST_SM[4]_net_1\, Y => 
        HIEFFPLA_NET_0_117749);
    
    \U_ELK6_CH/U_ELK1_CMD_TX/START_RISE\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117969, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_12, Q => 
        \U_ELK6_CH/U_ELK1_CMD_TX/START_RISE_net_1\);
    
    HIEFFPLA_INST_0_42397 : AO1A
      port map(A => HIEFFPLA_NET_0_119019, B => 
        \U50_PATTERNS/RD_USB_ADBUS[3]\, C => 
        HIEFFPLA_NET_0_119538, Y => HIEFFPLA_NET_0_119546);
    
    HIEFFPLA_INST_0_55368 : AND3
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[0]\, 
        B => \U_MASTER_DES/CCC_RX_CLK_LOCK\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[1]\, Y => 
        HIEFFPLA_NET_0_117048);
    
    \U200B_ELINKS/LOC_STOP_ADDR[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120183, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_7, Q => 
        \U200B_ELINKS/LOC_STOP_ADDR[4]\);
    
    HIEFFPLA_INST_0_62066 : MX2
      port map(A => HIEFFPLA_NET_0_116137, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_29[1]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_2[3]\, Y => 
        HIEFFPLA_NET_0_116040);
    
    HIEFFPLA_INST_0_45570 : AO1A
      port map(A => HIEFFPLA_NET_0_119428, B => 
        \U50_PATTERNS/ELINKS_STRT_ADDR[1]\, C => 
        HIEFFPLA_NET_0_118793, Y => HIEFFPLA_NET_0_118888);
    
    HIEFFPLA_INST_0_48829 : MX2
      port map(A => 
        \U_ELK19_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]_net_1\, B => 
        \U_ELK19_CH/ELK_TX_DAT[2]\, S => 
        \U_ELK19_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118246);
    
    HIEFFPLA_INST_0_60116 : MX2
      port map(A => HIEFFPLA_NET_0_116687, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_6[2]\, S => 
        HIEFFPLA_NET_0_117211, Y => HIEFFPLA_NET_0_116308);
    
    HIEFFPLA_INST_0_111274 : MX2A
      port map(A => HIEFFPLA_NET_0_115844, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_2[3]\, S => 
        HIEFFPLA_NET_0_117206, Y => HIEFFPLA_NET_0_116357);
    
    HIEFFPLA_INST_0_57962 : NAND3A
      port map(A => HIEFFPLA_NET_0_116592, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_7[4]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_7[3]\, Y => 
        HIEFFPLA_NET_0_116590);
    
    HIEFFPLA_INST_0_52024 : MX2C
      port map(A => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[40]_net_1\, B => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[41]_net_1\, S => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[0]\, Y => 
        HIEFFPLA_NET_0_117650);
    
    \U_ELK2_CH/U_ELK1_CMD_TX/SER_OUT_RDEL\ : DFN1C0
      port map(D => \U_ELK2_CH/U_ELK1_CMD_TX/SER_OUT_RI_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_8, Q
         => \U_ELK2_CH/ELK_OUT_R\);
    
    HIEFFPLA_INST_0_51112 : NAND2B
      port map(A => \OP_MODE_c_3[1]\, B => \PATT_ELK_DAT_9[7]\, Y
         => HIEFFPLA_NET_0_117826);
    
    \U_ELK15_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]\ : DFN1C0
      port map(D => \U_ELK15_CH/U_SLAVE_1ELK/Q[6]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]_net_1\);
    
    \U_ELK13_CH/U_SLAVE_1ELK/Q[0]\ : DFN1C0
      port map(D => \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/Q[0]_net_1\);
    
    \U_ELK4_CH/U_SLAVE_1ELK/Q[8]\ : DFN1C0
      port map(D => \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/Q[8]_net_1\);
    
    \U_ELK2_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118155, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_12, Q => 
        \U_ELK2_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]_net_1\);
    
    HIEFFPLA_INST_0_45336 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/SM_BANK_SEL[8]\, C => 
        \U50_PATTERNS/ELINK_DOUTA_11[0]\, Y => 
        HIEFFPLA_NET_0_118937);
    
    HIEFFPLA_INST_0_56626 : AND3
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[14]_net_1\, B
         => HIEFFPLA_NET_0_117424, C => HIEFFPLA_NET_0_117427, Y
         => HIEFFPLA_NET_0_116825);
    
    HIEFFPLA_INST_0_49116 : NAND2B
      port map(A => \OP_MODE_c_5[1]\, B => \PATT_ELK_DAT_1[3]\, Y
         => HIEFFPLA_NET_0_118190);
    
    \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[7]\ : DFN1C0
      port map(D => \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\);
    
    HIEFFPLA_INST_0_56561 : AND3
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[7]_net_1\, B => 
        HIEFFPLA_NET_0_117426, C => HIEFFPLA_NET_0_117425, Y => 
        HIEFFPLA_NET_0_116838);
    
    HIEFFPLA_INST_0_44979 : NAND3C
      port map(A => HIEFFPLA_NET_0_119452, B => 
        HIEFFPLA_NET_0_119389, C => HIEFFPLA_NET_0_119000, Y => 
        HIEFFPLA_NET_0_119007);
    
    HIEFFPLA_INST_0_54594 : NAND3
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[4]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[2]_net_1\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[1]_net_1\, Y => 
        HIEFFPLA_NET_0_117237);
    
    \U_ELK8_CH/U_ELK1_CMD_TX/SER_OUT_FI\ : DFN1C0
      port map(D => 
        \U_ELK8_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_3, Q => 
        \U_ELK8_CH/U_ELK1_CMD_TX/SER_OUT_FI_net_1\);
    
    HIEFFPLA_INST_0_37204 : NAND2B
      port map(A => HIEFFPLA_NET_0_120293, B => 
        HIEFFPLA_NET_0_120334, Y => HIEFFPLA_NET_0_120325);
    
    \U_ELK8_CH/U_ELK1_CMD_TX/SER_OUT_RDEL\ : DFN1C0
      port map(D => \U_ELK8_CH/U_ELK1_CMD_TX/SER_OUT_RI_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_2, Q
         => \U_ELK8_CH/ELK_OUT_R\);
    
    HIEFFPLA_INST_0_50591 : MX2
      port map(A => 
        \U_ELK7_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]_net_1\, B => 
        \U_ELK7_CH/ELK_TX_DAT[3]\, S => 
        \U_ELK7_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_117927);
    
    HIEFFPLA_INST_0_38206 : MX2
      port map(A => \U50_PATTERNS/CHKSUM[6]\, B => 
        HIEFFPLA_NET_0_120129, S => HIEFFPLA_NET_0_119470, Y => 
        HIEFFPLA_NET_0_120137);
    
    HIEFFPLA_INST_0_59918 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_3[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_19[1]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_5[4]_net_1\, Y
         => HIEFFPLA_NET_0_116334);
    
    \U_MASTER_DES/U13B_CCC/Core\ : DYNCCC
      generic map(VCOFREQUENCY => 160.0)

      port map(CLKA => CLK_40M_BUF_RECD, EXTFB => \GND\, 
        POWERDOWN => \VCC\, GLA => CCC_160M_ADJ, LOCK => 
        \U_MASTER_DES/CCC_RX_CLK_LOCK\, CLKB => \GND\, GLB => 
        OPEN, YB => OPEN, CLKC => \GND\, GLC => OPEN, YC => OPEN, 
        SDIN => \U_MASTER_DES/AUX_SDIN\, SCLK => \AFLSDF_INV_52\, 
        SSHIFT => \U_MASTER_DES/AUX_SSHIFT\, SUPDATE => 
        \U_MASTER_DES/AUX_SUPDATE\, MODE => 
        \U_MASTER_DES/AUX_MODE\, SDOUT => OPEN, OADIV0 => \GND\, 
        OADIV1 => \GND\, OADIV2 => \GND\, OADIV3 => \GND\, OADIV4
         => \GND\, OAMUX0 => \GND\, OAMUX1 => \GND\, OAMUX2 => 
        \VCC\, DLYGLA0 => \GND\, DLYGLA1 => \GND\, DLYGLA2 => 
        \GND\, DLYGLA3 => \GND\, DLYGLA4 => \GND\, OBDIV0 => 
        \GND\, OBDIV1 => \GND\, OBDIV2 => \GND\, OBDIV3 => \GND\, 
        OBDIV4 => \GND\, OBMUX0 => \GND\, OBMUX1 => \GND\, OBMUX2
         => \VCC\, DLYYB0 => \GND\, DLYYB1 => \GND\, DLYYB2 => 
        \GND\, DLYYB3 => \GND\, DLYYB4 => \GND\, DLYGLB0 => \GND\, 
        DLYGLB1 => \GND\, DLYGLB2 => \GND\, DLYGLB3 => \GND\, 
        DLYGLB4 => \GND\, OCDIV0 => \GND\, OCDIV1 => \GND\, 
        OCDIV2 => \GND\, OCDIV3 => \GND\, OCDIV4 => \GND\, OCMUX0
         => \GND\, OCMUX1 => \GND\, OCMUX2 => \VCC\, DLYYC0 => 
        \GND\, DLYYC1 => \GND\, DLYYC2 => \GND\, DLYYC3 => \GND\, 
        DLYYC4 => \GND\, DLYGLC0 => \GND\, DLYGLC1 => \GND\, 
        DLYGLC2 => \GND\, DLYGLC3 => \GND\, DLYGLC4 => \GND\, 
        FINDIV0 => \VCC\, FINDIV1 => \VCC\, FINDIV2 => \VCC\, 
        FINDIV3 => \GND\, FINDIV4 => \GND\, FINDIV5 => \GND\, 
        FINDIV6 => \GND\, FBDIV0 => \VCC\, FBDIV1 => \VCC\, 
        FBDIV2 => \VCC\, FBDIV3 => \VCC\, FBDIV4 => \VCC\, FBDIV5
         => \GND\, FBDIV6 => \GND\, FBDLY0 => \VCC\, FBDLY1 => 
        \VCC\, FBDLY2 => \VCC\, FBDLY3 => \GND\, FBDLY4 => \VCC\, 
        FBSEL0 => \GND\, FBSEL1 => \VCC\, XDLYSEL => \GND\, 
        VCOSEL0 => \GND\, VCOSEL1 => \GND\, VCOSEL2 => \VCC\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_24[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116103, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_8, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_24[2]\);
    
    \U200A_TFC/LOC_STOP_ADDR[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120286, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_1, Q => \U200A_TFC/LOC_STOP_ADDR[4]\);
    
    HIEFFPLA_INST_0_53848 : NAND2B
      port map(A => HIEFFPLA_NET_0_117371, B => 
        HIEFFPLA_NET_0_117407, Y => HIEFFPLA_NET_0_117343);
    
    HIEFFPLA_INST_0_60923 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_1[3]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_17[3]\, S
         => \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_3[4]_net_1\, 
        Y => HIEFFPLA_NET_0_116198);
    
    HIEFFPLA_INST_0_59992 : MX2
      port map(A => HIEFFPLA_NET_0_116687, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_4[2]\, S => 
        HIEFFPLA_NET_0_117202, Y => HIEFFPLA_NET_0_116324);
    
    \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[1]\ : DFN1C0
      port map(D => 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[1]_net_1\);
    
    HIEFFPLA_INST_0_56325 : AO1
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[4]_net_1\, B => 
        HIEFFPLA_NET_0_117429, C => HIEFFPLA_NET_0_116869, Y => 
        HIEFFPLA_NET_0_116893);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_29[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116044, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_16_0, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_29[1]\);
    
    HIEFFPLA_INST_0_44272 : MX2
      port map(A => \TFC_STRT_ADDR[4]\, B => 
        \U50_PATTERNS/U4A_REGCROSS/SAMP_TWO[4]_net_1\, S => 
        HIEFFPLA_NET_0_119156, Y => HIEFFPLA_NET_0_119150);
    
    \U_EXEC_MASTER/MPOR_B_31_0\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117787, CLK => CLK_40M_GL, CLR
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_0\, Q => 
        P_MASTER_POR_B_c_31_0);
    
    \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[6]\\\\/U0/U0\ : 
        IOPAD_BI_U
      port map(D => 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[6]\\\\/U0/NET1\, 
        E => 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[6]\\\\/U0/NET2\, 
        Y => 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[6]\\\\/U0/NET3\, 
        PAD => BIDIR_USB_ADBUS(6));
    
    HIEFFPLA_INST_0_57437 : AND3
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_4[3]\, B => 
        HIEFFPLA_NET_0_116683, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_4[4]\, Y => 
        HIEFFPLA_NET_0_116684);
    
    \U_ELK14_CH/U_SLAVE_1ELK/Q[12]\ : DFN1C0
      port map(D => \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/Q[12]_net_1\);
    
    \U50_PATTERNS/ELINK_DINA_15[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119823, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_16, Q => 
        \U50_PATTERNS/ELINK_DINA_15[0]\);
    
    HIEFFPLA_INST_0_58795 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_1[0]\, B => 
        HIEFFPLA_NET_0_116680, S => HIEFFPLA_NET_0_117158, Y => 
        HIEFFPLA_NET_0_116475);
    
    HIEFFPLA_INST_0_58425 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_14[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_30[1]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_3[4]_net_1\, Y
         => HIEFFPLA_NET_0_116523);
    
    HIEFFPLA_INST_0_46917 : MX2
      port map(A => \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\, 
        B => \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\, S => 
        \BIT_OS_SEL_4[2]\, Y => HIEFFPLA_NET_0_118585);
    
    HIEFFPLA_INST_0_50613 : AND2A
      port map(A => \OP_MODE_c_4[1]\, B => \PATT_ELK_DAT_7[6]\, Y
         => HIEFFPLA_NET_0_117917);
    
    HIEFFPLA_INST_0_46862 : MX2
      port map(A => 
        \U_ELK11_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]_net_1\, B => 
        \U_ELK11_CH/ELK_TX_DAT[5]\, S => 
        \U_ELK11_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118601);
    
    HIEFFPLA_INST_0_46776 : MX2
      port map(A => HIEFFPLA_NET_0_118622, B => 
        HIEFFPLA_NET_0_118634, S => \BIT_OS_SEL_0[0]\, Y => 
        \U_ELK10_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[4]\);
    
    HIEFFPLA_INST_0_37027 : AOI1A
      port map(A => HIEFFPLA_NET_0_120352, B => 
        HIEFFPLA_NET_0_120325, C => HIEFFPLA_NET_0_120365, Y => 
        HIEFFPLA_NET_0_120366);
    
    \U50_PATTERNS/ELINK_ADDRA_17[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120031, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_10, Q => 
        \U50_PATTERNS/ELINK_ADDRA_17[0]\);
    
    \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[4]\ : DFN1C0
      port map(D => 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\);
    
    \U_ELK12_CH/U_SLAVE_1ELK/Q[7]\ : DFN1C0
      port map(D => \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/Q[7]_net_1\);
    
    HIEFFPLA_INST_0_56413 : AND3
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[3]_net_1\, B => 
        HIEFFPLA_NET_0_117427, C => HIEFFPLA_NET_0_117423, Y => 
        HIEFFPLA_NET_0_116872);
    
    HIEFFPLA_INST_0_49242 : MX2
      port map(A => HIEFFPLA_NET_0_118172, B => 
        HIEFFPLA_NET_0_118185, S => \BIT_OS_SEL_1[0]\, Y => 
        \U_ELK1_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[1]\);
    
    HIEFFPLA_INST_0_42374 : AND3C
      port map(A => \U50_PATTERNS/RD_XFER_TYPE[4]_net_1\, B => 
        \U50_PATTERNS/RD_XFER_TYPE[7]_net_1\, C => 
        HIEFFPLA_NET_0_119551, Y => HIEFFPLA_NET_0_119552);
    
    HIEFFPLA_INST_0_61955 : MX2
      port map(A => HIEFFPLA_NET_0_117114, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_28[1]\, S => 
        HIEFFPLA_NET_0_117146, Y => HIEFFPLA_NET_0_116054);
    
    HIEFFPLA_INST_0_49772 : MX2
      port map(A => HIEFFPLA_NET_0_118082, B => 
        HIEFFPLA_NET_0_118093, S => \BIT_OS_SEL_1[0]\, Y => 
        \U_ELK3_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[5]\);
    
    AFLSDF_INV_65 : INV
      port map(A => \U200A_TFC/RX_SER_WORD_2DEL[1]_net_1\, Y => 
        \AFLSDF_INV_65\);
    
    \U_ELK1_CH/U_SLAVE_1ELK/RECD_SER_WORD[5]\ : DFN1C0
      port map(D => \U_ELK1_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[5]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_1[5]\);
    
    \U_ELK1_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]\ : DFN1C0
      port map(D => \U_ELK1_CH/U_SLAVE_1ELK/Q[7]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]_net_1\);
    
    \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[4]\ : DFN1C0
      port map(D => \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\);
    
    HIEFFPLA_INST_0_56719 : AND3A
      port map(A => HIEFFPLA_NET_0_116687, B => 
        HIEFFPLA_NET_0_116804, C => HIEFFPLA_NET_0_116776, Y => 
        HIEFFPLA_NET_0_116815);
    
    HIEFFPLA_INST_0_46328 : AO1
      port map(A => HIEFFPLA_NET_0_119250, B => 
        \U50_PATTERNS/ELINK_DOUTA_5[0]\, C => 
        HIEFFPLA_NET_0_118715, Y => HIEFFPLA_NET_0_118716);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_23[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116117, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_6, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_23[3]\);
    
    HIEFFPLA_INST_0_45728 : NAND2A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_18[4]\, Y => 
        HIEFFPLA_NET_0_118857);
    
    HIEFFPLA_INST_0_44496 : MX2
      port map(A => \ELKS_STRT_ADDR[6]\, B => 
        \U50_PATTERNS/U4C_REGCROSS/SAMP_TWO[6]_net_1\, S => 
        HIEFFPLA_NET_0_119114, Y => HIEFFPLA_NET_0_119106);
    
    AFLSDF_INV_43 : INV
      port map(A => DCB_SALT_SEL_c, Y => \AFLSDF_INV_43\);
    
    \U50_PATTERNS/ELINK_ADDRA_9[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119941, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_10, Q => 
        \U50_PATTERNS/ELINK_ADDRA_9[2]\);
    
    HIEFFPLA_INST_0_43688 : AND3C
      port map(A => HIEFFPLA_NET_0_119269, B => 
        HIEFFPLA_NET_0_119234, C => HIEFFPLA_NET_0_119261, Y => 
        HIEFFPLA_NET_0_119240);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_7[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116301, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_3, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_7[2]\);
    
    \U_ELK19_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118244, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_7, Q => 
        \U_ELK19_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]_net_1\);
    
    HIEFFPLA_INST_0_62905 : MX2
      port map(A => HIEFFPLA_NET_0_115894, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[13]\, S => 
        HIEFFPLA_NET_0_117073, Y => HIEFFPLA_NET_0_115930);
    
    \U50_PATTERNS/U4E_REGCROSS/LOCAL_REG_VAL_4[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119058, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_1, Q => \OP_MODE_c_4[1]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_14[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116234, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_2, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_14[1]\);
    
    \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[5]\ : DFN1C0
      port map(D => \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\);
    
    \U_ELK10_CH/U_ELK1_CMD_TX/SER_OUT_FI\ : DFN1C0
      port map(D => 
        \U_ELK10_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_11, Q
         => \U_ELK10_CH/U_ELK1_CMD_TX/SER_OUT_FI_net_1\);
    
    \U50_PATTERNS/ELINK_DINA_19[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119787, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_1, Q => 
        \U50_PATTERNS/ELINK_DINA_19[4]\);
    
    HIEFFPLA_INST_0_43090 : AND3
      port map(A => HIEFFPLA_NET_0_119370, B => 
        \U50_PATTERNS/REG_STATE[5]_net_1\, C => 
        HIEFFPLA_NET_0_119434, Y => HIEFFPLA_NET_0_119382);
    
    AFLSDF_INV_21 : INV
      port map(A => DCB_SALT_SEL_c, Y => \AFLSDF_INV_21\);
    
    \U50_PATTERNS/ELINK_ADDRA_14[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120054, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_5, Q => 
        \U50_PATTERNS/ELINK_ADDRA_14[1]\);
    
    HIEFFPLA_INST_0_60762 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_15[4]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_16[4]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[0]\, Y => 
        HIEFFPLA_NET_0_116224);
    
    HIEFFPLA_INST_0_37660 : AND2A
      port map(A => \ELKS_STRT_ADDR[3]\, B => 
        HIEFFPLA_NET_0_120219, Y => HIEFFPLA_NET_0_120238);
    
    HIEFFPLA_INST_0_49132 : MX2
      port map(A => HIEFFPLA_NET_0_118174, B => 
        HIEFFPLA_NET_0_118171, S => \BIT_OS_SEL_0[1]\, Y => 
        HIEFFPLA_NET_0_118184);
    
    \U_ELK3_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]\ : DFN1C0
      port map(D => \U_ELK3_CH/U_SLAVE_1ELK/Q[6]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]_net_1\);
    
    \U_ELK12_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118557, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_12, Q => 
        \U_ELK12_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]_net_1\);
    
    \U60_TS_RD_BUF/\\\\TRIBUFF_F_24U[0]\\\\/U0/U0\ : IOPAD_TRI_U
      port map(D => 
        \U60_TS_RD_BUF/\\\\TRIBUFF_F_24U[0]\\\\/U0/NET1\, E => 
        \U60_TS_RD_BUF/\\\\TRIBUFF_F_24U[0]\\\\/U0/NET2\, PAD => 
        USB_RD_B);
    
    HIEFFPLA_INST_0_59438 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_27[0]\, B => 
        HIEFFPLA_NET_0_116680, S => HIEFFPLA_NET_0_117162, Y => 
        HIEFFPLA_NET_0_116394);
    
    HIEFFPLA_INST_0_50977 : MX2
      port map(A => HIEFFPLA_NET_0_117846, B => 
        HIEFFPLA_NET_0_117870, S => \BIT_OS_SEL_5[0]\, Y => 
        \U_ELK8_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[0]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/BEST_CLKPHASE[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117448, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_10, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_CLKPHASE[4]\);
    
    HIEFFPLA_INST_0_39848 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_8[6]\, B => 
        HIEFFPLA_NET_0_119517, S => HIEFFPLA_NET_0_119291, Y => 
        HIEFFPLA_NET_0_119945);
    
    HIEFFPLA_INST_0_56907 : NAND3
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_1[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_1[2]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_1[3]\, Y => 
        HIEFFPLA_NET_0_116779);
    
    HIEFFPLA_INST_0_56681 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_0[5]\, B => 
        HIEFFPLA_NET_0_116795, S => HIEFFPLA_NET_0_117602, Y => 
        HIEFFPLA_NET_0_116819);
    
    HIEFFPLA_INST_0_43871 : MX2
      port map(A => HIEFFPLA_NET_0_119517, B => 
        \U50_PATTERNS/TFC_ADDRA[6]\, S => HIEFFPLA_NET_0_119294, 
        Y => HIEFFPLA_NET_0_119201);
    
    \U50_PATTERNS/TFC_ADDRA[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119203, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_9, Q => \U50_PATTERNS/TFC_ADDRA[4]\);
    
    HIEFFPLA_INST_0_48479 : MX2
      port map(A => HIEFFPLA_NET_0_118311, B => 
        HIEFFPLA_NET_0_118307, S => \BIT_OS_SEL_1[1]\, Y => 
        HIEFFPLA_NET_0_118305);
    
    \U50_PATTERNS/U4D_REGCROSS/SAMP_ONE[7]\ : DFN1C0
      port map(D => \U50_PATTERNS/ELINKS_STOP_ADDR[7]\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_25, Q => 
        \U50_PATTERNS/U4D_REGCROSS/SAMP_ONE[7]_net_1\);
    
    HIEFFPLA_INST_0_55119 : AOI1C
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[6]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[8]_net_1\, C => 
        HIEFFPLA_NET_0_116620, Y => HIEFFPLA_NET_0_117118);
    
    HIEFFPLA_INST_0_44432 : XO1
      port map(A => \TFC_STOP_ADDR[4]\, B => 
        \U50_PATTERNS/U4B_REGCROSS/SAMP_TWO[4]_net_1\, C => 
        HIEFFPLA_NET_0_119117, Y => HIEFFPLA_NET_0_119120);
    
    \U_ELK18_CH/ELK_IN_R\ : DFN1C0
      port map(D => \U_ELK18_CH/ELK_IN_DDR_R\, CLK => 
        CCC_160M_ADJ, CLR => DEV_RST_B_c, Q => 
        \U_ELK18_CH/ELK_IN_R_net_1\);
    
    HIEFFPLA_INST_0_56227 : NAND2
      port map(A => HIEFFPLA_NET_0_116928, B => 
        HIEFFPLA_NET_0_116927, Y => HIEFFPLA_NET_0_116925);
    
    \U50_PATTERNS/OP_MODE[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119617, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_15, Q => \U50_PATTERNS/OP_MODE[0]\);
    
    HIEFFPLA_INST_0_111248 : MX2A
      port map(A => HIEFFPLA_NET_0_115846, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_6[3]\, S => 
        HIEFFPLA_NET_0_117211, Y => HIEFFPLA_NET_0_116307);
    
    \U_GEN_REF_CLK/GEN_40M_REFCNT[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117727, CLK => Y, CLR => 
        DEV_RST_B_c, Q => \U_GEN_REF_CLK/GEN_40M_REFCNT[1]_net_1\);
    
    HIEFFPLA_INST_0_41892 : AOI1C
      port map(A => \U50_PATTERNS/ELINK_RWA[6]\, B => 
        HIEFFPLA_NET_0_119641, C => HIEFFPLA_NET_0_119671, Y => 
        HIEFFPLA_NET_0_119672);
    
    \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_2S_6\ : DFN1C0
      port map(D => 
        \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_1S_net_1\, CLK
         => CLK60MHZ, CLR => P_MASTER_POR_B_c_0_0, Q => 
        P_USB_MASTER_EN_c_6);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_21[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116142, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_3, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_21[3]\);
    
    HIEFFPLA_INST_0_42360 : NAND2A
      port map(A => HIEFFPLA_NET_0_119579, B => 
        HIEFFPLA_NET_0_119583, Y => HIEFFPLA_NET_0_119556);
    
    HIEFFPLA_INST_0_43072 : AO1A
      port map(A => HIEFFPLA_NET_0_119633, B => 
        HIEFFPLA_NET_0_119584, C => HIEFFPLA_NET_0_119386, Y => 
        HIEFFPLA_NET_0_119387);
    
    HIEFFPLA_INST_0_42243 : AND3B
      port map(A => \U50_PATTERNS/RD_USB_ADBUS[1]\, B => 
        HIEFFPLA_NET_0_119208, C => 
        \U50_PATTERNS/RD_USB_ADBUS[0]\, Y => 
        HIEFFPLA_NET_0_119593);
    
    \U_ELK17_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118336, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_17, Q => 
        \U_ELK17_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]_net_1\);
    
    \U_ELK4_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118061, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_17, Q => 
        \U_ELK4_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]_net_1\);
    
    HIEFFPLA_INST_0_46876 : AND2A
      port map(A => \OP_MODE_c[1]\, B => \PATT_ELK_DAT_11[4]\, Y
         => HIEFFPLA_NET_0_118594);
    
    \U_ELK2_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118157, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_12, Q => 
        \U_ELK2_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]_net_1\);
    
    \U_ELK17_CH/U_ELK1_SERDAT_SOURCE/SERDAT[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118327, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_11, Q => 
        \U_ELK17_CH/ELK_TX_DAT[1]\);
    
    HIEFFPLA_INST_0_43542 : MX2
      port map(A => \U50_PATTERNS/SM_BANK_SEL_0[21]\, B => 
        HIEFFPLA_NET_0_119018, S => HIEFFPLA_NET_0_118691, Y => 
        HIEFFPLA_NET_0_119299);
    
    \U_ELK1_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]\ : DFN1C0
      port map(D => \U_ELK1_CH/U_SLAVE_1ELK/Q[13]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]_net_1\);
    
    HIEFFPLA_INST_0_41853 : AOI1D
      port map(A => \U50_PATTERNS/ELINK_RWA[17]\, B => 
        HIEFFPLA_NET_0_119233, C => HIEFFPLA_NET_0_119652, Y => 
        HIEFFPLA_NET_0_119682);
    
    \U50_PATTERNS/ELINK_DINA_3[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119761, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_11, Q => 
        \U50_PATTERNS/ELINK_DINA_3[6]\);
    
    HIEFFPLA_INST_0_49595 : MX2
      port map(A => 
        \U_ELK3_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]_net_1\, B => 
        \U_ELK3_CH/ELK_TX_DAT[3]\, S => 
        \U_ELK3_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118107);
    
    \U50_PATTERNS/U4E_REGCROSS/DELCNT[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119071, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_25, Q => 
        \U50_PATTERNS/U4E_REGCROSS/DELCNT[0]_net_1\);
    
    HIEFFPLA_INST_0_62322 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_3[0]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_4[0]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_4[0]\, Y => 
        HIEFFPLA_NET_0_116004);
    
    HIEFFPLA_INST_0_51009 : MX2
      port map(A => HIEFFPLA_NET_0_117860, B => 
        HIEFFPLA_NET_0_117859, S => \BIT_OS_SEL_5[0]\, Y => 
        \U_ELK8_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[4]\);
    
    HIEFFPLA_INST_0_43569 : NAND2B
      port map(A => \U50_PATTERNS/SM_BANK_SEL[14]\, B => 
        \U50_PATTERNS/SM_BANK_SEL[11]\, Y => 
        HIEFFPLA_NET_0_119287);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_8[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116293, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_5, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_8[0]\);
    
    \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[8]\ : DFN1C0
      port map(D => \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\);
    
    HIEFFPLA_INST_0_62101 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_2[0]\, 
        B => HIEFFPLA_NET_0_117190, S => HIEFFPLA_NET_0_117176, Y
         => HIEFFPLA_NET_0_116035);
    
    HIEFFPLA_INST_0_41521 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_7[7]\, B => 
        HIEFFPLA_NET_0_119560, S => HIEFFPLA_NET_0_119289, Y => 
        HIEFFPLA_NET_0_119728);
    
    \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117058, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_27, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[3]_net_1\);
    
    HIEFFPLA_INST_0_63072 : XA1C
      port map(A => HIEFFPLA_NET_0_115912, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[12]\, C => 
        HIEFFPLA_NET_0_117078, Y => HIEFFPLA_NET_0_115895);
    
    HIEFFPLA_INST_0_48634 : MX2
      port map(A => HIEFFPLA_NET_0_118271, B => 
        HIEFFPLA_NET_0_118268, S => \BIT_OS_SEL_0[1]\, Y => 
        HIEFFPLA_NET_0_118274);
    
    HIEFFPLA_INST_0_48186 : MX2
      port map(A => HIEFFPLA_NET_0_118365, B => 
        HIEFFPLA_NET_0_118363, S => \BIT_OS_SEL_1[1]\, Y => 
        HIEFFPLA_NET_0_118356);
    
    \U_ELK7_CH/U_SLAVE_1ELK/Q[10]\ : DFN1C0
      port map(D => \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/Q[10]_net_1\);
    
    \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[13]\ : DFN1C0
      port map(D => \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\, 
        CLK => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[13]_net_1\);
    
    \U_ELK16_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118380, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_14, Q => 
        \U_ELK16_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]_net_1\);
    
    HIEFFPLA_INST_0_59265 : AO1B
      port map(A => HIEFFPLA_NET_0_117394, B => 
        HIEFFPLA_NET_0_116345, C => HIEFFPLA_NET_0_117366, Y => 
        HIEFFPLA_NET_0_116412);
    
    HIEFFPLA_INST_0_42848 : AND3B
      port map(A => \U50_PATTERNS/REG_STATE[1]_net_1\, B => 
        \U50_PATTERNS/REG_STATE[5]_net_1\, C => 
        \U50_PATTERNS/REG_STATE[0]_net_1\, Y => 
        HIEFFPLA_NET_0_119448);
    
    HIEFFPLA_INST_0_47387 : MX2
      port map(A => \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[3]_net_1\, 
        B => \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\, S => 
        \BIT_OS_SEL_3[2]\, Y => HIEFFPLA_NET_0_118499);
    
    \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[0]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_WRD_40M_FIXED[0]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_27, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[0]_net_1\);
    
    HIEFFPLA_INST_0_37177 : AO1C
      port map(A => \U200A_TFC/GP_PG_SM[0]_net_1\, B => 
        HIEFFPLA_NET_0_120291, C => \OP_MODE_c[2]\, Y => 
        HIEFFPLA_NET_0_120332);
    
    \U_MASTER_DES/U13A_ADJ_160M/BITCNT[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117693, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_14, Q => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[5]\);
    
    HIEFFPLA_INST_0_38092 : MX2
      port map(A => HIEFFPLA_NET_0_120153, B => ELKS_RAM_BLKB_EN, 
        S => HIEFFPLA_NET_0_120152, Y => HIEFFPLA_NET_0_120154);
    
    AFLSDF_INV_46 : INV
      port map(A => DCB_SALT_SEL_c, Y => \AFLSDF_INV_46\);
    
    HIEFFPLA_INST_0_37257 : AOI1D
      port map(A => HIEFFPLA_NET_0_120296, B => 
        HIEFFPLA_NET_0_120304, C => HIEFFPLA_NET_0_120330, Y => 
        HIEFFPLA_NET_0_120312);
    
    HIEFFPLA_INST_0_113035 : AO18
      port map(A => HIEFFPLA_NET_0_115813, B => 
        \U200B_ELINKS/LOC_STOP_ADDR[3]\, C => \ELKS_ADDRB[3]\, Y
         => HIEFFPLA_NET_0_115821);
    
    HIEFFPLA_INST_0_54071 : MX2
      port map(A => HIEFFPLA_NET_0_117417, B => 
        HIEFFPLA_NET_0_117256, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[1]_net_1\, Y
         => HIEFFPLA_NET_0_117312);
    
    HIEFFPLA_INST_0_48925 : MX2
      port map(A => HIEFFPLA_NET_0_118215, B => 
        HIEFFPLA_NET_0_118226, S => \BIT_OS_SEL_0[1]\, Y => 
        HIEFFPLA_NET_0_118223);
    
    HIEFFPLA_INST_0_40837 : MX2
      port map(A => HIEFFPLA_NET_0_119574, B => 
        \U50_PATTERNS/ELINK_DINA_17[3]\, S => 
        HIEFFPLA_NET_0_119260, Y => HIEFFPLA_NET_0_119804);
    
    \U_EXEC_MASTER/MPOR_B_19\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117787, CLK => CLK_40M_GL, CLR
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_1\, Q => 
        P_MASTER_POR_B_c_19);
    
    \U_ELK15_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]\ : DFN1C0
      port map(D => \U_ELK15_CH/U_SLAVE_1ELK/Q[8]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]_net_1\);
    
    HIEFFPLA_INST_0_41431 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_6[5]\, B => 
        HIEFFPLA_NET_0_119567, S => HIEFFPLA_NET_0_119258, Y => 
        HIEFFPLA_NET_0_119738);
    
    HIEFFPLA_INST_0_61223 : MX2
      port map(A => HIEFFPLA_NET_0_117186, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_20[3]\, S => 
        HIEFFPLA_NET_0_117141, Y => HIEFFPLA_NET_0_116157);
    
    HIEFFPLA_INST_0_62173 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_30[3]\, B => 
        HIEFFPLA_NET_0_117186, S => HIEFFPLA_NET_0_117330, Y => 
        HIEFFPLA_NET_0_116027);
    
    HIEFFPLA_INST_0_50359 : NAND2B
      port map(A => \OP_MODE_c_0[1]\, B => \PATT_ELK_DAT_6[1]\, Y
         => HIEFFPLA_NET_0_117967);
    
    \U_ELK16_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]\ : DFN1C0
      port map(D => \U_ELK16_CH/U_SLAVE_1ELK/Q[13]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]_net_1\);
    
    \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[1]\ : DFN1C0
      port map(D => 
        \U_ELK12_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\);
    
    HIEFFPLA_INST_0_58243 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_12[2]\, B => 
        HIEFFPLA_NET_0_116544, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_0[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116546);
    
    HIEFFPLA_INST_0_43246 : AOI1B
      port map(A => \U50_PATTERNS/REG_STATE_0[4]_net_1\, B => 
        HIEFFPLA_NET_0_119366, C => 
        \U50_PATTERNS/REG_STATE_0[5]_net_1\, Y => 
        HIEFFPLA_NET_0_119339);
    
    \U_EXEC_MASTER/USB_MASTER_EN/CNT_EN_60M0S\ : DFN1C0
      port map(D => 
        \U_EXEC_MASTER/USB_MASTER_EN/CNT_EN_40M_net_1\, CLK => 
        CLK60MHZ, CLR => P_MASTER_POR_B_c_23, Q => 
        \U_EXEC_MASTER/USB_MASTER_EN/CNT_EN_60M0S_net_1\);
    
    HIEFFPLA_INST_0_59041 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_6[0]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_22[0]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_2[4]_net_1\, Y
         => HIEFFPLA_NET_0_116443);
    
    \U_ELK1_CH/U_SLAVE_1ELK/Q[12]\ : DFN1C0
      port map(D => \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/Q[12]_net_1\);
    
    HIEFFPLA_INST_0_53118 : MX2
      port map(A => HIEFFPLA_NET_0_117547, B => 
        HIEFFPLA_NET_0_117543, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[3]\, Y => 
        HIEFFPLA_NET_0_117463);
    
    HIEFFPLA_INST_0_42533 : OA1A
      port map(A => HIEFFPLA_NET_0_119433, B => 
        HIEFFPLA_NET_0_119010, C => \U50_PATTERNS/REG_ADDR[5]\, Y
         => HIEFFPLA_NET_0_119518);
    
    HIEFFPLA_INST_0_161262 : DFN1C0
      port map(D => \ELK0_IN_F\, CLK => CCC_160M_ADJ, CLR => 
        P_MASTER_POR_B_c_31_0, Q => HIEFFPLA_NET_0_161293);
    
    \U50_PATTERNS/ELINK_ADDRA_19[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120014, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_13, Q => 
        \U50_PATTERNS/ELINK_ADDRA_19[1]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_28[4]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116051, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_15, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_28[4]\);
    
    \U_ELK10_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2\ : IOPADN_BI
      port map(DB => \U_ELK10_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, 
        E => \U_ELK10_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET3\, PAD
         => ELK10_DAT_N, N2POUT => 
        \U_ELK10_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2_N2P\);
    
    HIEFFPLA_INST_0_63164 : AND3
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[2]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[1]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[0]\, Y => 
        HIEFFPLA_NET_0_115870);
    
    \U_MASTER_DES/U13C_MASTER_DESER/BEST_BIT_OS_VAL[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_117578, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_14, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_BIT_OS_VAL[2]\);
    
    \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[7]\ : DFN1C0
      port map(D => \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\);
    
    \U_ELK12_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]\ : DFN1C0
      port map(D => \U_ELK12_CH/U_SLAVE_1ELK/Q[8]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]_net_1\);
    
    \U_ELK10_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118649, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_6, Q => 
        \U_ELK10_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]_net_1\);
    
    \U_ELK0_CMD_TX/SER_CMD_WORD_F[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118668, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_17, Q => 
        \U_ELK0_CMD_TX/SER_CMD_WORD_F[1]_net_1\);
    
    HIEFFPLA_INST_0_37189 : NAND2B
      port map(A => \U200A_TFC/GP_PG_SM[0]_net_1\, B => 
        \U200A_TFC/GP_PG_SM[1]_net_1\, Y => HIEFFPLA_NET_0_120329);
    
    \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[7]\ : DFN1C0
      port map(D => \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\);
    
    HIEFFPLA_INST_0_61382 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_5[2]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_21[2]\, S
         => \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_1[4]_net_1\, 
        Y => HIEFFPLA_NET_0_116134);
    
    HIEFFPLA_INST_0_45664 : AO1A
      port map(A => HIEFFPLA_NET_0_119475, B => 
        \U50_PATTERNS/ELINKS_STOP_ADDR[2]\, C => 
        HIEFFPLA_NET_0_118772, Y => HIEFFPLA_NET_0_118869);
    
    \U_ELK0_CMD_TX/START_RISE\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118661, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_3, Q => 
        \U_ELK0_CMD_TX/START_RISE_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_24[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116434, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_18, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_24[0]\);
    
    HIEFFPLA_INST_0_43755 : AND3A
      port map(A => \U50_PATTERNS/RD_USB_ADBUS[3]\, B => 
        HIEFFPLA_NET_0_119594, C => 
        \U50_PATTERNS/RD_USB_ADBUS[2]\, Y => 
        HIEFFPLA_NET_0_119222);
    
    HIEFFPLA_INST_0_39326 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_1[4]\, B => 
        HIEFFPLA_NET_0_119519, S => HIEFFPLA_NET_0_119243, Y => 
        HIEFFPLA_NET_0_120003);
    
    HIEFFPLA_INST_0_51641 : MX2
      port map(A => 
        \U_EXEC_MASTER/USB_MASTER_EN/CNT_EN_60M2S_net_1\, B => 
        \U_EXEC_MASTER/USB_MASTER_EN/T_CNT60M[6]_net_1\, S => 
        HIEFFPLA_NET_0_117753, Y => HIEFFPLA_NET_0_117732);
    
    \U_ELK5_CH/U_ELK1_SERDAT_SOURCE/SERDAT[7]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118006, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i, Q => 
        \U_ELK5_CH/ELK_TX_DAT[7]\);
    
    \U50_PATTERNS/ELINK_DINA_13[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119835, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_14, Q => 
        \U50_PATTERNS/ELINK_DINA_13[4]\);
    
    \U_ELK12_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118561, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_15, Q => 
        \U_ELK12_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]_net_1\);
    
    HIEFFPLA_INST_0_56005 : MX2
      port map(A => HIEFFPLA_NET_0_116984, B => 
        HIEFFPLA_NET_0_117029, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[4]\, Y => 
        HIEFFPLA_NET_0_116962);
    
    \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM[6]\ : DFN1P0
      port map(D => HIEFFPLA_NET_0_117617, CLK => CLK_40M_GL, PRE
         => P_MASTER_POR_B_c_22_0, Q => 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM[6]_net_1\);
    
    \U50_PATTERNS/TFC_STRT_ADDR[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119167, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_13, Q => 
        \U50_PATTERNS/TFC_STRT_ADDR[5]\);
    
    \U_ELK13_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]\ : DFN1C0
      port map(D => \U_ELK13_CH/U_SLAVE_1ELK/Q[11]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]_net_1\);
    
    \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[12]\ : DFN1C0
      port map(D => 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]_net_1\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[12]_net_1\);
    
    \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[3]\ : DFN1C0
      port map(D => 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[3]_net_1\);
    
    HIEFFPLA_INST_0_61016 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_2[1]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_18[1]\, S
         => \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_4[4]_net_1\, 
        Y => HIEFFPLA_NET_0_116185);
    
    \U_ELK7_CH/U_SLAVE_1ELK/RECD_SER_WORD[6]\ : DFN1C0
      port map(D => \U_ELK7_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[6]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_7[6]\);
    
    HIEFFPLA_INST_0_46391 : AO1
      port map(A => HIEFFPLA_NET_0_119276, B => 
        \U50_PATTERNS/ELINK_DOUTA_10[3]\, C => 
        HIEFFPLA_NET_0_118850, Y => HIEFFPLA_NET_0_118700);
    
    HIEFFPLA_INST_0_41919 : AND3C
      port map(A => HIEFFPLA_NET_0_119253, B => 
        HIEFFPLA_NET_0_119262, C => \U50_PATTERNS/SM_BANK_SEL[4]\, 
        Y => HIEFFPLA_NET_0_119662);
    
    \U_ELK14_CH/U_ELK1_CMD_TX/SER_OUT_RI\ : DFN1C0
      port map(D => 
        \U_ELK14_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_10, Q
         => \U_ELK14_CH/U_ELK1_CMD_TX/SER_OUT_RI_net_1\);
    
    \U_ELK7_CH/U_SLAVE_1ELK/Q[1]\ : DFN1C0
      port map(D => \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/Q[1]_net_1\);
    
    HIEFFPLA_INST_0_52642 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_13[2]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_14[2]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_2[0]\, Y => 
        HIEFFPLA_NET_0_117534);
    
    \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[4]\ : DFN1C0
      port map(D => \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\);
    
    HIEFFPLA_INST_0_41440 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_6[6]\, B => 
        HIEFFPLA_NET_0_119566, S => HIEFFPLA_NET_0_119258, Y => 
        HIEFFPLA_NET_0_119737);
    
    \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[8]\ : DFN1C0
      port map(D => 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_115923, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_9, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[7]\);
    
    HIEFFPLA_INST_0_58266 : MX2
      port map(A => HIEFFPLA_NET_0_116815, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_12[3]\, S => 
        HIEFFPLA_NET_0_117210, Y => HIEFFPLA_NET_0_116543);
    
    \U50_PATTERNS/ELINK_DINA_9[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119719, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_19, Q => 
        \U50_PATTERNS/ELINK_DINA_9[0]\);
    
    HIEFFPLA_INST_0_54117 : MX2
      port map(A => HIEFFPLA_NET_0_116198, B => 
        HIEFFPLA_NET_0_116082, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_1[3]_net_1\, Y
         => HIEFFPLA_NET_0_117306);
    
    HIEFFPLA_INST_0_47870 : NAND2B
      port map(A => \OP_MODE_c_6[1]\, B => \PATT_ELK_DAT_15[2]\, 
        Y => HIEFFPLA_NET_0_118416);
    
    \U_MASTER_DES/U13C_MASTER_DESER/ARB_WRD_40M_FIXED[10]\ : 
        DFN1C0
      port map(D => \U_MASTER_DES/U13C_MASTER_DESER/Q[10]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_28, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_WRD_40M_FIXED[10]_net_1\);
    
    \U_ELK14_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118466, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_2, Q => 
        \U_ELK14_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]_net_1\);
    
    \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[11]\ : DFN1C0
      port map(D => \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\);
    
    \U50_PATTERNS/ELINK_ADDRA_19[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120011, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_13, Q => 
        \U50_PATTERNS/ELINK_ADDRA_19[4]\);
    
    HIEFFPLA_INST_0_55667 : MX2
      port map(A => HIEFFPLA_NET_0_115990, B => 
        HIEFFPLA_NET_0_116236, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_2[3]\, Y => 
        HIEFFPLA_NET_0_117006);
    
    HIEFFPLA_INST_0_47619 : AND2A
      port map(A => \OP_MODE_c_2[1]\, B => \PATT_ELK_DAT_14[0]\, 
        Y => HIEFFPLA_NET_0_118463);
    
    HIEFFPLA_INST_0_47374 : AND2A
      port map(A => \OP_MODE_c[1]\, B => \PATT_ELK_DAT_13[4]\, Y
         => HIEFFPLA_NET_0_118504);
    
    HIEFFPLA_INST_0_61679 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_25[2]\, B => 
        HIEFFPLA_NET_0_117181, S => HIEFFPLA_NET_0_117117, Y => 
        HIEFFPLA_NET_0_116093);
    
    HIEFFPLA_INST_0_55218 : AND2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[6]_net_1\, B => 
        HIEFFPLA_NET_0_117321, Y => HIEFFPLA_NET_0_117083);
    
    \U50_PATTERNS/U4D_REGCROSS/SAMP_TWO[0]\ : DFN1C0
      port map(D => \U50_PATTERNS/U4D_REGCROSS/SAMP_ONE[0]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_30, Q => 
        \U50_PATTERNS/U4D_REGCROSS/SAMP_TWO[0]_net_1\);
    
    HIEFFPLA_INST_0_56350 : AO1
      port map(A => HIEFFPLA_NET_0_117431, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[2]_net_1\, C => 
        HIEFFPLA_NET_0_116864, Y => HIEFFPLA_NET_0_116888);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_2[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116035, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_10, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_2[0]\);
    
    HIEFFPLA_INST_0_47845 : MX2
      port map(A => HIEFFPLA_NET_0_118425, B => 
        \U_ELK15_CH/ELK_TX_DAT[6]\, S => 
        \U_ELK15_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118424);
    
    AFLSDF_INV_39 : INV
      port map(A => DCB_SALT_SEL_c, Y => \AFLSDF_INV_39\);
    
    HIEFFPLA_INST_0_56118 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/MAX_CNT[6]\, 
        B => HIEFFPLA_NET_0_116933, S => HIEFFPLA_NET_0_117084, Y
         => HIEFFPLA_NET_0_116948);
    
    HIEFFPLA_INST_0_53062 : MX2
      port map(A => HIEFFPLA_NET_0_117562, B => 
        HIEFFPLA_NET_0_117558, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[2]\, Y => 
        HIEFFPLA_NET_0_117470);
    
    \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[13]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_WRD_40M_FIXED[13]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_32_0, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[13]_net_1\);
    
    \U_ELK18_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]\ : DFN1C0
      port map(D => \U_ELK18_CH/U_SLAVE_1ELK/Q[6]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]_net_1\);
    
    HIEFFPLA_INST_0_40558 : MX2
      port map(A => HIEFFPLA_NET_0_119570, B => 
        \U50_PATTERNS/ELINK_DINA_13[4]\, S => 
        HIEFFPLA_NET_0_119285, Y => HIEFFPLA_NET_0_119835);
    
    HIEFFPLA_INST_0_46461 : AND3C
      port map(A => HIEFFPLA_NET_0_118673, B => 
        HIEFFPLA_NET_0_119577, C => HIEFFPLA_NET_0_118678, Y => 
        HIEFFPLA_NET_0_118686);
    
    HIEFFPLA_INST_0_39281 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_19[7]\, B => 
        HIEFFPLA_NET_0_119516, S => HIEFFPLA_NET_0_119293, Y => 
        HIEFFPLA_NET_0_120008);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_19[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116481, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_20, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_19[0]\);
    
    \U_ELK15_CH/U_SLAVE_1ELK/Q[2]\ : DFN1C0
      port map(D => \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/Q[2]_net_1\);
    
    \U_ELK14_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118468, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_2, Q => 
        \U_ELK14_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]_net_1\);
    
    HIEFFPLA_INST_0_46427 : NAND3B
      port map(A => HIEFFPLA_NET_0_118695, B => 
        \U50_PATTERNS/WR_XFER_TYPE[3]_net_1\, C => 
        \U50_PATTERNS/WR_XFER_TYPE[7]_net_1\, Y => 
        HIEFFPLA_NET_0_118692);
    
    \U_MASTER_DES/U13C_MASTER_DESER/RECD_SER_WORD[4]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_116900, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_30, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/RECD_SER_WORD[4]_net_1\);
    
    \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[8]\ : DFN1C0
      port map(D => \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\);
    
    \U_ELK13_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118514, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_1, Q => 
        \U_ELK13_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_18[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116493, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_19, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_18[2]\);
    
    HIEFFPLA_INST_0_63153 : AND3
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[2]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[1]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_3[0]\, Y => 
        HIEFFPLA_NET_0_115874);
    
    \U_ELK9_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL\ : DFN1C0
      port map(D => 
        \U_ELK9_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL_net_1\);
    
    HIEFFPLA_INST_0_40141 : AOI1D
      port map(A => HIEFFPLA_NET_0_119389, B => 
        HIEFFPLA_NET_0_119464, C => 
        \U50_PATTERNS/SM_BANK_SEL[17]\, Y => 
        HIEFFPLA_NET_0_119893);
    
    \U50_PATTERNS/ELINK_DINA_4[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119753, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_13, Q => 
        \U50_PATTERNS/ELINK_DINA_4[6]\);
    
    HIEFFPLA_INST_0_52378 : MX2
      port map(A => HIEFFPLA_NET_0_117527, B => 
        HIEFFPLA_NET_0_117483, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[1]\, Y => 
        HIEFFPLA_NET_0_117571);
    
    HIEFFPLA_INST_0_51321 : NAND3C
      port map(A => \U_EXEC_MASTER/PRESCALE[0]\, B => 
        \U_EXEC_MASTER/PRESCALE[1]\, C => HIEFFPLA_NET_0_117763, 
        Y => HIEFFPLA_NET_0_117797);
    
    HIEFFPLA_INST_0_46712 : MX2
      port map(A => \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\, 
        B => \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[13]_net_1\, S => 
        \BIT_OS_SEL_6[2]\, Y => HIEFFPLA_NET_0_118624);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_29[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116042, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_16_0, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_29[3]\);
    
    HIEFFPLA_INST_0_46627 : AND2A
      port map(A => \OP_MODE_c_3[1]\, B => \PATT_ELK_DAT_10[4]\, 
        Y => HIEFFPLA_NET_0_118639);
    
    \U50_PATTERNS/ELINK_ADDRA_7[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119956, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_6, Q => 
        \U50_PATTERNS/ELINK_ADDRA_7[3]\);
    
    HIEFFPLA_INST_0_58289 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_13[2]\, B => 
        HIEFFPLA_NET_0_116535, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_1[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116540);
    
    HIEFFPLA_INST_0_51282 : MX2
      port map(A => HIEFFPLA_NET_0_117820, B => 
        HIEFFPLA_NET_0_117800, S => \BIT_OS_SEL_4[0]\, Y => 
        \U_ELK9_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[7]\);
    
    \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[3]\ : DFN1C0
      port map(D => 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[3]_net_1\);
    
    \U0A_40M_REFCLK/\\\\BIBUF_LVDS[0]\\\\/U0/U2\ : IOPADN_BI
      port map(DB => 
        \U0A_40M_REFCLK/\\\\BIBUF_LVDS[0]\\\\/U0/NET1\, E => 
        \U0A_40M_REFCLK/\\\\BIBUF_LVDS[0]\\\\/U0/NET3\, PAD => 
        BIDIR_CLK40M_N, N2POUT => 
        \U0A_40M_REFCLK/\\\\BIBUF_LVDS[0]\\\\/U0/U2_N2P\);
    
    HIEFFPLA_INST_0_55620 : MX2
      port map(A => HIEFFPLA_NET_0_116193, B => 
        HIEFFPLA_NET_0_116083, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_1[3]\, Y => 
        HIEFFPLA_NET_0_117013);
    
    HIEFFPLA_INST_0_43099 : AND2A
      port map(A => \U50_PATTERNS/REG_STATE[1]_net_1\, B => 
        \U50_PATTERNS/REG_STATE[0]_net_1\, Y => 
        HIEFFPLA_NET_0_119378);
    
    HIEFFPLA_INST_0_63097 : XA1C
      port map(A => HIEFFPLA_NET_0_115920, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[5]\, C => 
        HIEFFPLA_NET_0_117078, Y => HIEFFPLA_NET_0_115889);
    
    HIEFFPLA_INST_0_54181 : MX2
      port map(A => HIEFFPLA_NET_0_116174, B => 
        HIEFFPLA_NET_0_116063, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_1[3]_net_1\, Y
         => HIEFFPLA_NET_0_117298);
    
    HIEFFPLA_INST_0_50606 : AND2
      port map(A => CLK_40M_GL, B => 
        \U_ELK7_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0_net_1\, Y => 
        HIEFFPLA_NET_0_117924);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_3[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116008, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_11, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_3[2]\);
    
    \U_ELK13_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]\ : DFN1C0
      port map(D => \U_ELK13_CH/U_SLAVE_1ELK/Q[8]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]_net_1\);
    
    HIEFFPLA_INST_0_51933 : AND2A
      port map(A => \U_MASTER_DES/U13A_ADJ_160M/BITCNT[6]\, B => 
        HIEFFPLA_NET_0_117655, Y => HIEFFPLA_NET_0_117663);
    
    \U_ELK19_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]\ : DFN1C0
      port map(D => \U_ELK19_CH/U_SLAVE_1ELK/Q[8]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]_net_1\);
    
    AFLSDF_INV_37 : INV
      port map(A => DCB_SALT_SEL_c, Y => \AFLSDF_INV_37\);
    
    HIEFFPLA_INST_0_50568 : AND2
      port map(A => \U_ELK7_CH/ELK_TX_DAT[0]\, B => 
        \U_ELK7_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_117932);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_5[6]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116655, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_11, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_5[6]\);
    
    \U_ELK9_CH/U_ELK1_SERDAT_SOURCE/SERDAT[6]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117827, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_7, Q => 
        \U_ELK9_CH/ELK_TX_DAT[6]\);
    
    \U_ELK3_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL\ : DFN1C0
      port map(D => \U_ELK3_CH/ELK_IN_R_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL_net_1\);
    
    HIEFFPLA_INST_0_54975 : AND2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_3[6]_net_1\, B => 
        HIEFFPLA_NET_0_117214, Y => HIEFFPLA_NET_0_117150);
    
    HIEFFPLA_INST_0_38579 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_10[1]\, B => 
        HIEFFPLA_NET_0_119523, S => HIEFFPLA_NET_0_119239, Y => 
        HIEFFPLA_NET_0_120086);
    
    HIEFFPLA_INST_0_42599 : AND3B
      port map(A => HIEFFPLA_NET_0_119498, B => 
        HIEFFPLA_NET_0_119452, C => HIEFFPLA_NET_0_119509, Y => 
        HIEFFPLA_NET_0_119503);
    
    \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[13]\ : DFN1C0
      port map(D => \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\, 
        CLK => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[13]_net_1\);
    
    \U_ELK11_CH/U_SLAVE_1ELK/RECD_SER_WORD[5]\ : DFN1C0
      port map(D => \U_ELK11_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[5]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_11[5]\);
    
    HIEFFPLA_INST_0_39128 : MX2
      port map(A => HIEFFPLA_NET_0_119517, B => 
        \U50_PATTERNS/ELINK_ADDRA_17[6]\, S => 
        HIEFFPLA_NET_0_119260, Y => HIEFFPLA_NET_0_120025);
    
    \U_EXEC_MASTER/MPOR_B_15\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117787, CLK => CLK_40M_GL, CLR
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_1\, Q => 
        P_MASTER_POR_B_c_15);
    
    HIEFFPLA_INST_0_40168 : AOI1C
      port map(A => \U50_PATTERNS/ELINK_BLKA[8]\, B => 
        HIEFFPLA_NET_0_119638, C => HIEFFPLA_NET_0_119881, Y => 
        HIEFFPLA_NET_0_119882);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_16[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116212, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_5, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_16[3]\);
    
    HIEFFPLA_INST_0_54577 : AND3B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[1]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[0]_net_1\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[3]_net_1\, Y => 
        HIEFFPLA_NET_0_117242);
    
    HIEFFPLA_INST_0_38006 : MX2
      port map(A => \U200B_ELINKS/LOC_STRT_ADDR[4]\, B => 
        \ELKS_STRT_ADDR[4]\, S => 
        \U200B_ELINKS/GP_PG_SM_0[10]_net_1\, Y => 
        HIEFFPLA_NET_0_120175);
    
    HIEFFPLA_INST_0_59945 : MX2
      port map(A => HIEFFPLA_NET_0_116815, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_3[3]\, S => 
        HIEFFPLA_NET_0_117207, Y => HIEFFPLA_NET_0_116330);
    
    HIEFFPLA_INST_0_47756 : MX2
      port map(A => HIEFFPLA_NET_0_118443, B => 
        HIEFFPLA_NET_0_118440, S => \BIT_OS_SEL_4[0]\, Y => 
        \U_ELK14_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[2]\);
    
    HIEFFPLA_INST_0_46331 : AO1A
      port map(A => HIEFFPLA_NET_0_118860, B => 
        \U50_PATTERNS/SM_BANK_SEL[15]\, C => 
        HIEFFPLA_NET_0_118853, Y => HIEFFPLA_NET_0_118715);
    
    HIEFFPLA_INST_0_40594 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_14[0]\, B => 
        HIEFFPLA_NET_0_119578, S => HIEFFPLA_NET_0_119249, Y => 
        HIEFFPLA_NET_0_119831);
    
    \U_ELK14_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]\ : DFN1C0
      port map(D => \U_ELK14_CH/U_SLAVE_1ELK/Q[1]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]_net_1\);
    
    \U_EXEC_MASTER/MPOR_SALT_B_12\ : DFI1P0
      port map(D => HIEFFPLA_NET_0_117781, CLK => CLK_40M_GL, PRE
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_2\, QN => 
        MASTER_SALT_POR_B_i_0_i_12);
    
    \U_ELK13_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118516, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_1, Q => 
        \U_ELK13_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_7[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116302, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_3, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_7[1]\);
    
    \U50_PATTERNS/ELINK_DINA_6[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119743, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_16, Q => 
        \U50_PATTERNS/ELINK_DINA_6[0]\);
    
    HIEFFPLA_INST_0_56931 : NAND3C
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_1[8]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_1[7]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_1[6]\, Y => 
        HIEFFPLA_NET_0_116772);
    
    HIEFFPLA_INST_0_49756 : MX2
      port map(A => HIEFFPLA_NET_0_118080, B => 
        HIEFFPLA_NET_0_118086, S => \BIT_OS_SEL_1[0]\, Y => 
        \U_ELK3_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[3]\);
    
    \U_ELK6_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]\ : DFN1C0
      port map(D => \U_ELK6_CH/U_SLAVE_1ELK/Q[14]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]_net_1\);
    
    \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[2]\ : DFN1C0
      port map(D => 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[2]_net_1\);
    
    \U_ELK12_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]\ : DFN1C0
      port map(D => \U_ELK12_CH/U_SLAVE_1ELK/Q[11]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]_net_1\);
    
    HIEFFPLA_INST_0_48369 : NAND2B
      port map(A => \OP_MODE_c_6[1]\, B => \PATT_ELK_DAT_17[3]\, 
        Y => HIEFFPLA_NET_0_118325);
    
    \U_ELK7_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]\ : DFN1C0
      port map(D => \U_ELK7_CH/U_SLAVE_1ELK/Q[5]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]_net_1\);
    
    HIEFFPLA_INST_0_42744 : AO1A
      port map(A => HIEFFPLA_NET_0_119450, B => 
        HIEFFPLA_NET_0_119469, C => HIEFFPLA_NET_0_119452, Y => 
        HIEFFPLA_NET_0_119470);
    
    HIEFFPLA_INST_0_56206 : AOI1A
      port map(A => HIEFFPLA_NET_0_116940, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/MAX_CNT[5]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/MAX_CNT[6]\, Y => 
        HIEFFPLA_NET_0_116930);
    
    HIEFFPLA_INST_0_47188 : MX2
      port map(A => \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\, 
        B => \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[11]_net_1\, S => 
        \BIT_OS_SEL_4[2]\, Y => HIEFFPLA_NET_0_118537);
    
    HIEFFPLA_INST_0_43328 : XA1B
      port map(A => \U50_PATTERNS/SI_CNT[2]\, B => 
        HIEFFPLA_NET_0_119323, C => HIEFFPLA_NET_0_119329, Y => 
        HIEFFPLA_NET_0_119325);
    
    HIEFFPLA_INST_0_47732 : MX2
      port map(A => HIEFFPLA_NET_0_118452, B => 
        HIEFFPLA_NET_0_118449, S => \BIT_OS_SEL_2[1]\, Y => 
        HIEFFPLA_NET_0_118440);
    
    \U_ELK9_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117839, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_4, Q => 
        \U_ELK9_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]_net_1\);
    
    HIEFFPLA_INST_0_55794 : MX2
      port map(A => HIEFFPLA_NET_0_116004, B => 
        HIEFFPLA_NET_0_116260, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[3]\, Y => 
        HIEFFPLA_NET_0_116989);
    
    \U_ELK17_CH/U_SLAVE_1ELK/Q[4]\ : DFN1C0
      port map(D => \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/Q[4]_net_1\);
    
    \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[6]\ : DFN1C0
      port map(D => \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\);
    
    HIEFFPLA_INST_0_50070 : AND2
      port map(A => \U_ELK5_CH/ELK_TX_DAT[0]\, B => 
        \U_ELK5_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118022);
    
    HIEFFPLA_INST_0_46180 : AO1
      port map(A => HIEFFPLA_NET_0_119241, B => 
        \U50_PATTERNS/ELINK_DOUTA_1[5]\, C => 
        HIEFFPLA_NET_0_118925, Y => HIEFFPLA_NET_0_118748);
    
    \U_ELK16_CH/U_ELK1_SERDAT_SOURCE/SERDAT[7]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118366, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_9, Q => 
        \U_ELK16_CH/ELK_TX_DAT[7]\);
    
    HIEFFPLA_INST_0_38402 : MX2
      port map(A => \U50_PATTERNS/ELINKS_STRT_ADDR[4]\, B => 
        \U50_PATTERNS/ELINKS_STRT_ADDR_T[4]\, S => 
        HIEFFPLA_NET_0_119472, Y => HIEFFPLA_NET_0_120107);
    
    HIEFFPLA_INST_0_47848 : AND2
      port map(A => \U_ELK15_CH/ELK_TX_DAT[1]\, B => 
        \U_ELK15_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118423);
    
    HIEFFPLA_INST_0_59339 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_26[2]\, B => 
        HIEFFPLA_NET_0_116400, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_2[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116404);
    
    HIEFFPLA_INST_0_55177 : NAND2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[8]_net_1\, B => 
        \OP_MODE_c[5]\, Y => HIEFFPLA_NET_0_117104);
    
    HIEFFPLA_INST_0_51999 : MX2A
      port map(A => HIEFFPLA_NET_0_117644, B => 
        HIEFFPLA_NET_0_117643, S => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[1]\, Y => 
        HIEFFPLA_NET_0_117655);
    
    HIEFFPLA_INST_0_42387 : AO1A
      port map(A => HIEFFPLA_NET_0_119019, B => 
        \U50_PATTERNS/RD_USB_ADBUS[1]\, C => 
        HIEFFPLA_NET_0_119540, Y => HIEFFPLA_NET_0_119548);
    
    \U50_PATTERNS/U4E_REGCROSS/SAMP_ONE[1]\ : DFN1C0
      port map(D => \U50_PATTERNS/OP_MODE[1]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c, Q => 
        \U50_PATTERNS/U4E_REGCROSS/SAMP_ONE[1]_net_1\);
    
    HIEFFPLA_INST_0_44968 : AO1A
      port map(A => HIEFFPLA_NET_0_119423, B => 
        HIEFFPLA_NET_0_119632, C => HIEFFPLA_NET_0_119009, Y => 
        HIEFFPLA_NET_0_119010);
    
    HIEFFPLA_INST_0_37062 : AND3C
      port map(A => HIEFFPLA_NET_0_120336, B => 
        HIEFFPLA_NET_0_120341, C => HIEFFPLA_NET_0_120350, Y => 
        HIEFFPLA_NET_0_120354);
    
    \U_MASTER_DES/U13C_MASTER_DESER/ARB_WRD_40M_FIXED[7]\ : 
        DFN1C0
      port map(D => \U_MASTER_DES/U13C_MASTER_DESER/Q[7]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_26, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_WRD_40M_FIXED[7]_net_1\);
    
    \U_ELK15_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]\ : DFN1C0
      port map(D => \U_ELK15_CH/U_SLAVE_1ELK/Q[11]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]_net_1\);
    
    \U50_PATTERNS/U4B_REGCROSS/LOCAL_REG_VAL[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119126, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_19, Q => \TFC_STOP_ADDR[7]\);
    
    HIEFFPLA_INST_0_59567 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_29[1]\, B => 
        HIEFFPLA_NET_0_116370, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_0[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116377);
    
    HIEFFPLA_INST_0_50021 : MX2
      port map(A => HIEFFPLA_NET_0_118042, B => 
        HIEFFPLA_NET_0_118036, S => \BIT_OS_SEL_0[0]\, Y => 
        \U_ELK4_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[5]\);
    
    HIEFFPLA_INST_0_58786 : MX2
      port map(A => HIEFFPLA_NET_0_116815, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_19[3]\, S => 
        HIEFFPLA_NET_0_117205, Y => HIEFFPLA_NET_0_116476);
    
    \U_MASTER_DES/U13C_MASTER_DESER/MAX_CNT[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_116949, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_16, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/MAX_CNT[5]\);
    
    \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[11]\ : DFN1C0
      port map(D => 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[11]_net_1\);
    
    \U50_PATTERNS/U4D_REGCROSS/SAMP_TWO[7]\ : DFN1C0
      port map(D => \U50_PATTERNS/U4D_REGCROSS/SAMP_ONE[7]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_30, Q => 
        \U50_PATTERNS/U4D_REGCROSS/SAMP_TWO[7]_net_1\);
    
    HIEFFPLA_INST_0_42343 : AND2A
      port map(A => \U50_PATTERNS/RD_USB_ADBUS[0]\, B => 
        \U50_PATTERNS/RD_USB_ADBUS[1]\, Y => 
        HIEFFPLA_NET_0_119564);
    
    \U50_PATTERNS/ELINK_ADDRA_13[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120061, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_3, Q => 
        \U50_PATTERNS/ELINK_ADDRA_13[2]\);
    
    HIEFFPLA_INST_0_39056 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_16[6]\, B => 
        HIEFFPLA_NET_0_119517, S => HIEFFPLA_NET_0_119257, Y => 
        HIEFFPLA_NET_0_120033);
    
    HIEFFPLA_INST_0_49989 : MX2
      port map(A => HIEFFPLA_NET_0_118038, B => 
        HIEFFPLA_NET_0_118035, S => \BIT_OS_SEL_0[0]\, Y => 
        \U_ELK4_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[1]\);
    
    HIEFFPLA_INST_0_42430 : AND2
      port map(A => HIEFFPLA_NET_0_119473, B => 
        \U50_PATTERNS/RD_XFER_TYPE[5]_net_1\, Y => 
        HIEFFPLA_NET_0_119536);
    
    HIEFFPLA_INST_0_42402 : AO1A
      port map(A => HIEFFPLA_NET_0_119019, B => 
        \U50_PATTERNS/RD_USB_ADBUS[4]\, C => 
        HIEFFPLA_NET_0_119537, Y => HIEFFPLA_NET_0_119545);
    
    \U_ELK15_CH/U_SLAVE_1ELK/Q[10]\ : DFN1C0
      port map(D => \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/Q[10]_net_1\);
    
    \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[9]\ : DFN1C0
      port map(D => \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\);
    
    \U200B_ELINKS/RX_SER_WORD_2DEL[5]\ : DFN1C0
      port map(D => \U200B_ELINKS/RX_SER_WORD_1DEL[5]_net_1\, CLK
         => CLK_40M_GL, CLR => P_MASTER_POR_B_c_26, Q => 
        \U200B_ELINKS/RX_SER_WORD_2DEL[5]_net_1\);
    
    HIEFFPLA_INST_0_55304 : AND3
      port map(A => HIEFFPLA_NET_0_117415, B => 
        HIEFFPLA_NET_0_117359, C => HIEFFPLA_NET_0_117136, Y => 
        HIEFFPLA_NET_0_117066);
    
    HIEFFPLA_INST_0_54893 : AO1A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_0[6]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_0[8]_net_1\, C => 
        HIEFFPLA_NET_0_117177, Y => HIEFFPLA_NET_0_117178);
    
    \U50_PATTERNS/TFC_STOP_ADDR[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119182, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_8, Q => 
        \U50_PATTERNS/TFC_STOP_ADDR[6]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_5[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116322, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_1, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_5[0]\);
    
    HIEFFPLA_INST_0_50465 : MX2
      port map(A => \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\, B
         => \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[13]_net_1\, S => 
        \BIT_OS_SEL_5[2]\, Y => HIEFFPLA_NET_0_117946);
    
    HIEFFPLA_INST_0_45019 : AND3A
      port map(A => \U50_PATTERNS/USB_TXE_B\, B => 
        HIEFFPLA_NET_0_119378, C => HIEFFPLA_NET_0_119424, Y => 
        HIEFFPLA_NET_0_118998);
    
    \U_ELK16_CH/U_SLAVE_1ELK/Q[4]\ : DFN1C0
      port map(D => \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/Q[4]_net_1\);
    
    HIEFFPLA_INST_0_57115 : AND2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_2[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_2[0]\, Y => 
        HIEFFPLA_NET_0_116738);
    
    HIEFFPLA_INST_0_52884 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_27[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_28[1]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_1[0]\, Y => 
        HIEFFPLA_NET_0_117495);
    
    HIEFFPLA_INST_0_42458 : MX2
      port map(A => \U50_PATTERNS/REG_ADDR[2]\, B => 
        HIEFFPLA_NET_0_119507, S => HIEFFPLA_NET_0_119007, Y => 
        HIEFFPLA_NET_0_119531);
    
    HIEFFPLA_INST_0_40089 : AO1A
      port map(A => HIEFFPLA_NET_0_119873, B => 
        HIEFFPLA_NET_0_119240, C => HIEFFPLA_NET_0_119232, Y => 
        HIEFFPLA_NET_0_119910);
    
    HIEFFPLA_INST_0_39092 : MX2
      port map(A => HIEFFPLA_NET_0_119522, B => 
        \U50_PATTERNS/ELINK_ADDRA_17[2]\, S => 
        HIEFFPLA_NET_0_119260, Y => HIEFFPLA_NET_0_120029);
    
    \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[9]\ : DFN1C0
      port map(D => 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\);
    
    HIEFFPLA_INST_0_58151 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_10[0]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_26[0]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_2[4]_net_1\, Y
         => HIEFFPLA_NET_0_116558);
    
    HIEFFPLA_INST_0_49282 : MX2
      port map(A => HIEFFPLA_NET_0_118170, B => 
        HIEFFPLA_NET_0_118184, S => \BIT_OS_SEL_2[0]\, Y => 
        \U_ELK1_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[6]\);
    
    TFC_IN_F : DFN1C0
      port map(D => TFC_IN_DDR_F, CLK => CCC_160M_ADJ, CLR => 
        DEV_RST_B_c, Q => \TFC_IN_F\);
    
    \U_ELK5_CH/U_SLAVE_1ELK/RECD_SER_WORD[6]\ : DFN1C0
      port map(D => \U_ELK5_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[6]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_5[6]\);
    
    \U_ELK12_CH/U_SLAVE_1ELK/RECD_SER_WORD[5]\ : DFN1C0
      port map(D => \U_ELK12_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[5]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_12[5]\);
    
    \U_ELK6_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2\ : IOPADN_BI
      port map(DB => \U_ELK6_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, 
        E => \U_ELK6_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET3\, PAD => 
        ELK6_DAT_N, N2POUT => 
        \U_ELK6_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2_N2P\);
    
    HIEFFPLA_INST_0_56963 : AO1A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_1[3]\, B => 
        HIEFFPLA_NET_0_116769, C => HIEFFPLA_NET_0_117179, Y => 
        HIEFFPLA_NET_0_116764);
    
    HIEFFPLA_INST_0_47121 : AND2A
      port map(A => \OP_MODE_c_2[1]\, B => \PATT_ELK_DAT_12[0]\, 
        Y => HIEFFPLA_NET_0_118553);
    
    \U_ELK17_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL\ : DFN1C0
      port map(D => \U_ELK17_CH/ELK_IN_F_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL_net_1\);
    
    HIEFFPLA_INST_0_39452 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_3[2]\, B => 
        HIEFFPLA_NET_0_119522, S => HIEFFPLA_NET_0_119247, Y => 
        HIEFFPLA_NET_0_119989);
    
    HIEFFPLA_INST_0_111365 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_18[1]\, B => 
        HIEFFPLA_NET_0_116677, S => HIEFFPLA_NET_0_117204, Y => 
        HIEFFPLA_NET_0_116490);
    
    \U_ELK16_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]\ : DFN1C0
      port map(D => \U_ELK16_CH/U_SLAVE_1ELK/Q[7]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]_net_1\);
    
    HIEFFPLA_INST_0_63236 : AND2
      port map(A => CLK_40M_GL, B => 
        \U_TFC_CMD_TX/CLK40M_GEN_DEL0_net_1\, Y => 
        \U_TFC_CMD_TX/N_START_RISE\);
    
    HIEFFPLA_INST_0_49856 : MX2
      port map(A => 
        \U_ELK4_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]_net_1\, B => 
        \U_ELK4_CH/ELK_TX_DAT[7]\, S => 
        \U_ELK4_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118060);
    
    \U_MASTER_DES/U13C_MASTER_DESER/BEST_CLKPHASE[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117451, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_10, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_CLKPHASE[1]\);
    
    \U_EXEC_MASTER/MPOR_SALT_B_4\ : DFI1P0
      port map(D => HIEFFPLA_NET_0_117781, CLK => CLK_40M_GL, PRE
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_2\, QN => 
        MASTER_SALT_POR_B_i_0_i_4);
    
    HIEFFPLA_INST_0_50993 : MX2
      port map(A => HIEFFPLA_NET_0_117868, B => 
        HIEFFPLA_NET_0_117865, S => \BIT_OS_SEL_5[0]\, Y => 
        \U_ELK8_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[2]\);
    
    HIEFFPLA_INST_0_56761 : AND2B
      port map(A => HIEFFPLA_NET_0_116740, B => 
        HIEFFPLA_NET_0_116813, Y => HIEFFPLA_NET_0_116804);
    
    \U_ELK6_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U3\ : IOBI_ID_OD_EB
      port map(DR => \U_ELK6_CH/ELK_OUT_R\, DF => 
        \U_ELK6_CH/ELK_OUT_F\, CLR => \GND\, E => \AFLSDF_INV_45\, 
        ICLK => CCC_160M_ADJ, OCLK => CCC_160M_FXD, YIN => 
        \U_ELK6_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\, DOUT => OPEN, 
        EOUT => \U_ELK6_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET3\, YR
         => OPEN, YF => OPEN);
    
    \U50_PATTERNS/TFC_STRT_ADDR[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119172, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_13, Q => 
        \U50_PATTERNS/TFC_STRT_ADDR[0]\);
    
    HIEFFPLA_INST_0_47905 : MX2
      port map(A => \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\, 
        B => \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\, S => 
        \BIT_OS_SEL_1[2]\, Y => HIEFFPLA_NET_0_118406);
    
    \U_ELK4_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]\ : DFN1C0
      port map(D => \U_ELK4_CH/U_SLAVE_1ELK/Q[9]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]_net_1\);
    
    \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[5]\ : DFN1C0
      port map(D => \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\);
    
    HIEFFPLA_INST_0_57485 : AND2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_4[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_4[0]\, Y => 
        HIEFFPLA_NET_0_116671);
    
    \U_ELK8_CH/U_SLAVE_1ELK/RECD_SER_WORD[6]\ : DFN1C0
      port map(D => \U_ELK8_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[6]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_8[6]\);
    
    \U200B_ELINKS/RX_SER_WORD_2DEL[3]\ : DFN1C0
      port map(D => \U200B_ELINKS/RX_SER_WORD_1DEL[3]_net_1\, CLK
         => CLK_40M_GL, CLR => P_MASTER_POR_B_c_25, Q => 
        \U200B_ELINKS/RX_SER_WORD_2DEL[3]_net_1\);
    
    HIEFFPLA_INST_0_50680 : MX2
      port map(A => HIEFFPLA_NET_0_117908, B => 
        HIEFFPLA_NET_0_117904, S => \BIT_OS_SEL_4[1]\, Y => 
        HIEFFPLA_NET_0_117906);
    
    \U_ELK10_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118651, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_6, Q => 
        \U_ELK10_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]_net_1\);
    
    HIEFFPLA_INST_0_48471 : MX2
      port map(A => HIEFFPLA_NET_0_118318, B => 
        HIEFFPLA_NET_0_118316, S => \BIT_OS_SEL_1[1]\, Y => 
        HIEFFPLA_NET_0_118306);
    
    HIEFFPLA_INST_0_40123 : AOI1A
      port map(A => \U50_PATTERNS/ELINK_BLKA[18]\, B => 
        HIEFFPLA_NET_0_119231, C => HIEFFPLA_NET_0_119875, Y => 
        HIEFFPLA_NET_0_119899);
    
    \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[4]\ : DFN1C0
      port map(D => 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\);
    
    HIEFFPLA_INST_0_46026 : AND3
      port map(A => \U50_PATTERNS/TFC_DOUTA[6]\, B => 
        HIEFFPLA_NET_0_118997, C => HIEFFPLA_NET_0_119365, Y => 
        HIEFFPLA_NET_0_118783);
    
    \U200B_ELINKS/RX_SER_WORD_2DEL[1]\ : DFN1C0
      port map(D => \U200B_ELINKS/RX_SER_WORD_1DEL[1]_net_1\, CLK
         => CLK_40M_GL, CLR => P_MASTER_POR_B_c_25, Q => 
        \U200B_ELINKS/RX_SER_WORD_2DEL[1]_net_1\);
    
    HIEFFPLA_INST_0_58887 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_4[3]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_20[3]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_2[4]_net_1\, Y
         => HIEFFPLA_NET_0_116463);
    
    HIEFFPLA_INST_0_55492 : MX2
      port map(A => HIEFFPLA_NET_0_116106, B => 
        HIEFFPLA_NET_0_116012, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[3]\, Y => 
        HIEFFPLA_NET_0_117030);
    
    HIEFFPLA_INST_0_59486 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_11[2]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_27[2]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_5[4]_net_1\, Y
         => HIEFFPLA_NET_0_116388);
    
    HIEFFPLA_INST_0_50214 : MX2
      port map(A => HIEFFPLA_NET_0_118003, B => 
        HIEFFPLA_NET_0_118000, S => \BIT_OS_SEL_6[1]\, Y => 
        HIEFFPLA_NET_0_117991);
    
    \U_ELK2_CH/U_SLAVE_1ELK/Q[8]\ : DFN1C0
      port map(D => \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/Q[8]_net_1\);
    
    \U_ELK17_CH/U_ELK1_SERDAT_SOURCE/SERDAT[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118328, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_11, Q => 
        \U_ELK17_CH/ELK_TX_DAT[0]\);
    
    HIEFFPLA_INST_0_55727 : AO1
      port map(A => HIEFFPLA_NET_0_117087, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_4[0]\, C => 
        HIEFFPLA_NET_0_116997, Y => HIEFFPLA_NET_0_116998);
    
    HIEFFPLA_INST_0_45926 : AND3A
      port map(A => HIEFFPLA_NET_0_119376, B => 
        \U50_PATTERNS/TFC_STRT_ADDR[3]\, C => 
        HIEFFPLA_NET_0_119431, Y => HIEFFPLA_NET_0_118809);
    
    \U_ELK9_CH/U_SLAVE_1ELK/RECD_SER_WORD[2]\ : DFN1C0
      port map(D => \U_ELK9_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[2]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_9[2]\);
    
    HIEFFPLA_INST_0_48800 : MX2
      port map(A => HIEFFPLA_NET_0_118249, B => 
        HIEFFPLA_NET_0_118272, S => \BIT_OS_SEL_0[1]\, Y => 
        HIEFFPLA_NET_0_118251);
    
    HIEFFPLA_INST_0_50861 : AND2A
      port map(A => \OP_MODE_c_0[1]\, B => \PATT_ELK_DAT_8[5]\, Y
         => HIEFFPLA_NET_0_117873);
    
    HIEFFPLA_INST_0_56345 : AO1
      port map(A => HIEFFPLA_NET_0_117429, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[8]_net_1\, C => 
        HIEFFPLA_NET_0_116865, Y => HIEFFPLA_NET_0_116889);
    
    \EXTCLK_40MHZ_pad/U0/U1\ : IOTRI_OB_EB
      port map(D => EXTCLK_40MHZ_c, E => \VCC\, DOUT => 
        \EXTCLK_40MHZ_pad/U0/NET1\, EOUT => 
        \EXTCLK_40MHZ_pad/U0/NET2\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_3[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116723, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_7, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_3[2]\);
    
    \U_ELK16_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL\ : DFN1C0
      port map(D => 
        \U_ELK16_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL_net_1\);
    
    \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[3]\ : DFN1C0
      port map(D => 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[3]_net_1\);
    
    \U50_PATTERNS/ELINK_DINA_17[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119803, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_19, Q => 
        \U50_PATTERNS/ELINK_DINA_17[4]\);
    
    HIEFFPLA_INST_0_44652 : AND2A
      port map(A => \U50_PATTERNS/U4E_REGCROSS/DELCNT[0]_net_1\, 
        B => \U50_PATTERNS/U4E_REGCROSS/SYNC_SM[0]_net_1\, Y => 
        HIEFFPLA_NET_0_119071);
    
    HIEFFPLA_INST_0_37122 : AND3B
      port map(A => \U200A_TFC/LOC_STRT_ADDR[5]\, B => 
        HIEFFPLA_NET_0_120293, C => HIEFFPLA_NET_0_120328, Y => 
        HIEFFPLA_NET_0_120343);
    
    HIEFFPLA_INST_0_53642 : MX2
      port map(A => HIEFFPLA_NET_0_116219, B => 
        HIEFFPLA_NET_0_116112, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[3]_net_1\, Y
         => HIEFFPLA_NET_0_117379);
    
    AFLSDF_INV_61 : INV
      port map(A => \U200B_ELINKS/RX_SER_WORD_2DEL[1]_net_1\, Y
         => \AFLSDF_INV_61\);
    
    HIEFFPLA_INST_0_55699 : MX2
      port map(A => HIEFFPLA_NET_0_115973, B => 
        HIEFFPLA_NET_0_116216, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_2[3]\, Y => 
        HIEFFPLA_NET_0_117002);
    
    HIEFFPLA_INST_0_43084 : AND3A
      port map(A => \U50_PATTERNS/REG_STATE[0]_net_1\, B => 
        \U50_PATTERNS/REG_STATE[3]_net_1\, C => 
        \U50_PATTERNS/REG_STATE[5]_net_1\, Y => 
        HIEFFPLA_NET_0_119384);
    
    HIEFFPLA_INST_0_62932 : MX2
      port map(A => HIEFFPLA_NET_0_115891, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[3]\, S => 
        HIEFFPLA_NET_0_117073, Y => HIEFFPLA_NET_0_115927);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_12[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116548, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_10, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_12[0]\);
    
    \U_ELK11_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]\ : DFN1C0
      port map(D => \U_ELK11_CH/U_SLAVE_1ELK/Q[1]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]_net_1\);
    
    \U200A_TFC/LOC_STRT_ADDR[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120281, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_4, Q => \U200A_TFC/LOC_STRT_ADDR[1]\);
    
    \USBCLK60MHZ_pad/U0/U0\ : IOPAD_IN_U
      port map(PAD => USBCLK60MHZ, Y => \USBCLK60MHZ_pad/U0/NET1\);
    
    \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[9]\ : DFN1C0
      port map(D => 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\);
    
    \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[4]\ : DFN1C0
      port map(D => \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_2[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117010, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_16_0, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_2[0]\);
    
    HIEFFPLA_INST_0_56438 : AND3
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[8]_net_1\, B => 
        HIEFFPLA_NET_0_117427, C => HIEFFPLA_NET_0_117423, Y => 
        HIEFFPLA_NET_0_116867);
    
    HIEFFPLA_INST_0_50814 : MX2
      port map(A => \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\, 
        B => \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[14]_net_1\, S => 
        \BIT_OS_SEL_6[2]\, Y => HIEFFPLA_NET_0_117888);
    
    HIEFFPLA_INST_0_50603 : MX2
      port map(A => 
        \U_ELK7_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]_net_1\, B => 
        \U_ELK7_CH/ELK_TX_DAT[7]\, S => 
        \U_ELK7_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_117925);
    
    \U_ELK6_CH/U_SLAVE_1ELK/Q[5]\ : DFN1C0
      port map(D => \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/Q[5]_net_1\);
    
    HIEFFPLA_INST_0_54197 : MX2
      port map(A => HIEFFPLA_NET_0_116132, B => 
        HIEFFPLA_NET_0_116241, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_1[3]_net_1\, Y
         => HIEFFPLA_NET_0_117296);
    
    \U50_PATTERNS/TFC_DINA[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119195, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_4, Q => \U50_PATTERNS/TFC_DINA[2]\);
    
    HIEFFPLA_INST_0_63084 : XA1B
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[2]\, 
        B => HIEFFPLA_NET_0_115918, C => HIEFFPLA_NET_0_117078, Y
         => HIEFFPLA_NET_0_115892);
    
    HIEFFPLA_INST_0_37035 : AO1A
      port map(A => \TFC_STRT_ADDR[2]\, B => 
        HIEFFPLA_NET_0_120349, C => HIEFFPLA_NET_0_120346, Y => 
        HIEFFPLA_NET_0_120363);
    
    HIEFFPLA_INST_0_59035 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_6[3]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_22[3]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_2[4]_net_1\, Y
         => HIEFFPLA_NET_0_116444);
    
    HIEFFPLA_INST_0_53525 : AND3A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[2]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[4]_net_1\, C => 
        HIEFFPLA_NET_0_117318, Y => HIEFFPLA_NET_0_117394);
    
    HIEFFPLA_INST_0_47354 : MX2
      port map(A => 
        \U_ELK13_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]_net_1\, B => 
        \U_ELK13_CH/ELK_TX_DAT[3]\, S => 
        \U_ELK13_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118512);
    
    HIEFFPLA_INST_0_41674 : MX2
      port map(A => HIEFFPLA_NET_0_119691, B => 
        \U50_PATTERNS/ELINK_RWA[0]\, S => 
        \U50_PATTERNS/SM_BANK_SEL_0[20]\, Y => 
        HIEFFPLA_NET_0_119711);
    
    HIEFFPLA_INST_0_49850 : MX2
      port map(A => 
        \U_ELK4_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]_net_1\, B => 
        \U_ELK4_CH/ELK_TX_DAT[5]\, S => 
        \U_ELK4_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118061);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_14[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116233, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_2, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_14[2]\);
    
    \U_EXEC_MASTER/MPOR_B_30\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117787, CLK => CLK_40M_GL, CLR
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_0\, Q => 
        P_MASTER_POR_B_c_30);
    
    \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[1]\ : DFN1C0
      port map(D => 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[1]_net_1\);
    
    HIEFFPLA_INST_0_56611 : AND3
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[11]_net_1\, B
         => HIEFFPLA_NET_0_117424, C => HIEFFPLA_NET_0_117427, Y
         => HIEFFPLA_NET_0_116828);
    
    HIEFFPLA_INST_0_55642 : AO1
      port map(A => HIEFFPLA_NET_0_117087, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_2[0]\, C => 
        HIEFFPLA_NET_0_116997, Y => HIEFFPLA_NET_0_117010);
    
    HIEFFPLA_INST_0_40196 : AOI1D
      port map(A => HIEFFPLA_NET_0_119389, B => 
        HIEFFPLA_NET_0_119464, C => \U50_PATTERNS/SM_BANK_SEL[2]\, 
        Y => HIEFFPLA_NET_0_119876);
    
    \U_ELK19_CH/U_SLAVE_1ELK/RECD_SER_WORD[6]\ : DFN1C0
      port map(D => \U_ELK19_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[6]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_19[6]\);
    
    \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[1]\ : DFN1C0
      port map(D => 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[1]_net_1\);
    
    HIEFFPLA_INST_0_60642 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_13[4]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_29[4]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_2[4]_net_1\, Y
         => HIEFFPLA_NET_0_116239);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_19[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116179, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_11, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_19[1]\);
    
    HIEFFPLA_INST_0_39407 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_2[5]\, B => 
        HIEFFPLA_NET_0_119518, S => HIEFFPLA_NET_0_119278, Y => 
        HIEFFPLA_NET_0_119994);
    
    HIEFFPLA_INST_0_111272 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_30[0]\, B => 
        HIEFFPLA_NET_0_116735, S => HIEFFPLA_NET_0_117328, Y => 
        HIEFFPLA_NET_0_116346);
    
    \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[11]\ : DFN1C0
      port map(D => 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]_net_1\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[11]_net_1\);
    
    HIEFFPLA_INST_0_50925 : MX2
      port map(A => \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\, B
         => \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\, S => 
        \BIT_OS_SEL_3[2]\, Y => HIEFFPLA_NET_0_117862);
    
    HIEFFPLA_INST_0_47599 : AND2
      port map(A => \U_ELK14_CH/ELK_TX_DAT[1]\, B => 
        \U_ELK14_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118468);
    
    \U_ELK12_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118555, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_12, Q => 
        \U_ELK12_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]_net_1\);
    
    \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[2]\ : DFN1C0
      port map(D => \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\);
    
    HIEFFPLA_INST_0_50156 : MX2
      port map(A => \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[3]_net_1\, B
         => \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\, S => 
        \BIT_OS_SEL_6[2]\, Y => HIEFFPLA_NET_0_118000);
    
    \U50_PATTERNS/U114_PATT_ELINK_BLK/DPRT_512X9_SRAM_R0C0\ : 
        RAM4K9
      generic map(MEMORYFILE => "DPRT_512X9_SRAM_R0C0.mem")

      port map(ADDRA11 => AFLSDF_GND, ADDRA10 => AFLSDF_GND, 
        ADDRA9 => AFLSDF_GND, ADDRA8 => \GND\, ADDRA7 => 
        \U50_PATTERNS/ELINK_ADDRA_14[7]\, ADDRA6 => 
        \U50_PATTERNS/ELINK_ADDRA_14[6]\, ADDRA5 => 
        \U50_PATTERNS/ELINK_ADDRA_14[5]\, ADDRA4 => 
        \U50_PATTERNS/ELINK_ADDRA_14[4]\, ADDRA3 => 
        \U50_PATTERNS/ELINK_ADDRA_14[3]\, ADDRA2 => 
        \U50_PATTERNS/ELINK_ADDRA_14[2]\, ADDRA1 => 
        \U50_PATTERNS/ELINK_ADDRA_14[1]\, ADDRA0 => 
        \U50_PATTERNS/ELINK_ADDRA_14[0]\, ADDRB11 => AFLSDF_GND, 
        ADDRB10 => AFLSDF_GND, ADDRB9 => AFLSDF_GND, ADDRB8 => 
        \GND\, ADDRB7 => \ELKS_ADDRB[7]\, ADDRB6 => 
        \ELKS_ADDRB_0[6]\, ADDRB5 => \ELKS_ADDRB[5]\, ADDRB4 => 
        \ELKS_ADDRB_0[4]\, ADDRB3 => \ELKS_ADDRB[3]\, ADDRB2 => 
        \ELKS_ADDRB_0[2]\, ADDRB1 => \ELKS_ADDRB[1]\, ADDRB0 => 
        \ELKS_ADDRB[0]\, DINA8 => \GND\, DINA7 => 
        \U50_PATTERNS/ELINK_DINA_14[7]\, DINA6 => 
        \U50_PATTERNS/ELINK_DINA_14[6]\, DINA5 => 
        \U50_PATTERNS/ELINK_DINA_14[5]\, DINA4 => 
        \U50_PATTERNS/ELINK_DINA_14[4]\, DINA3 => 
        \U50_PATTERNS/ELINK_DINA_14[3]\, DINA2 => 
        \U50_PATTERNS/ELINK_DINA_14[2]\, DINA1 => 
        \U50_PATTERNS/ELINK_DINA_14[1]\, DINA0 => 
        \U50_PATTERNS/ELINK_DINA_14[0]\, DINB8 => \GND\, DINB7
         => \ELK_RX_SER_WORD_14[7]\, DINB6 => 
        \ELK_RX_SER_WORD_14[6]\, DINB5 => \ELK_RX_SER_WORD_14[5]\, 
        DINB4 => \ELK_RX_SER_WORD_14[4]\, DINB3 => 
        \ELK_RX_SER_WORD_14[3]\, DINB2 => \ELK_RX_SER_WORD_14[2]\, 
        DINB1 => \ELK_RX_SER_WORD_14[1]\, DINB0 => 
        \ELK_RX_SER_WORD_14[0]\, WIDTHA0 => \VCC\, WIDTHA1 => 
        \VCC\, WIDTHB0 => \VCC\, WIDTHB1 => \VCC\, PIPEA => \VCC\, 
        PIPEB => \VCC\, WMODEA => \GND\, WMODEB => \GND\, BLKA
         => \U50_PATTERNS/ELINK_BLKA[14]\, BLKB => 
        ELKS_RAM_BLKB_EN, WENA => \U50_PATTERNS/ELINK_RWA[14]\, 
        WENB => ELKS_RWB, CLKA => CLK60MHZ, CLKB => CLK_40M_GL, 
        RESET => P_USB_MASTER_EN_c_0, DOUTA8 => OPEN, DOUTA7 => 
        \U50_PATTERNS/ELINK_DOUTA_14[7]\, DOUTA6 => 
        \U50_PATTERNS/ELINK_DOUTA_14[6]\, DOUTA5 => 
        \U50_PATTERNS/ELINK_DOUTA_14[5]\, DOUTA4 => 
        \U50_PATTERNS/ELINK_DOUTA_14[4]\, DOUTA3 => 
        \U50_PATTERNS/ELINK_DOUTA_14[3]\, DOUTA2 => 
        \U50_PATTERNS/ELINK_DOUTA_14[2]\, DOUTA1 => 
        \U50_PATTERNS/ELINK_DOUTA_14[1]\, DOUTA0 => 
        \U50_PATTERNS/ELINK_DOUTA_14[0]\, DOUTB8 => OPEN, DOUTB7
         => \PATT_ELK_DAT_14[7]\, DOUTB6 => \PATT_ELK_DAT_14[6]\, 
        DOUTB5 => \PATT_ELK_DAT_14[5]\, DOUTB4 => 
        \PATT_ELK_DAT_14[4]\, DOUTB3 => \PATT_ELK_DAT_14[3]\, 
        DOUTB2 => \PATT_ELK_DAT_14[2]\, DOUTB1 => 
        \PATT_ELK_DAT_14[1]\, DOUTB0 => \PATT_ELK_DAT_14[0]\);
    
    HIEFFPLA_INST_0_56247 : AND2A
      port map(A => DCB_SALT_SEL_c, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/RECD_SER_WORD[6]_net_1\, 
        Y => \TFC_RX_SER_WORD[6]\);
    
    HIEFFPLA_INST_0_44014 : MX2
      port map(A => \U50_PATTERNS/TFC_STOP_ADDR[4]\, B => 
        \U50_PATTERNS/TFC_STOP_ADDR_T[4]\, S => 
        HIEFFPLA_NET_0_119472, Y => HIEFFPLA_NET_0_119184);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_3[5]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116720, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_7, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_3[5]\);
    
    \U_ELK16_CH/U_SLAVE_1ELK/RECD_SER_WORD[6]\ : DFN1C0
      port map(D => \U_ELK16_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[6]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_16[6]\);
    
    \U200A_TFC/RX_SER_WORD_3DEL[6]\ : DFN1C0
      port map(D => \U200A_TFC/RX_SER_WORD_2DEL[6]_net_1\, CLK
         => CLK_40M_GL, CLR => P_MASTER_POR_B_c_24, Q => 
        \U200A_TFC/RX_SER_WORD_3DEL[6]_net_1\);
    
    HIEFFPLA_INST_0_40297 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_0[7]\, B => 
        HIEFFPLA_NET_0_119560, S => HIEFFPLA_NET_0_119272, Y => 
        HIEFFPLA_NET_0_119864);
    
    \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[5]\ : DFN1C0
      port map(D => 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\);
    
    HIEFFPLA_INST_0_50527 : MX2
      port map(A => HIEFFPLA_NET_0_117960, B => 
        HIEFFPLA_NET_0_117958, S => \BIT_OS_SEL[0]\, Y => 
        \U_ELK6_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[6]\);
    
    \U_ELK1_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]\ : DFN1C0
      port map(D => \U_ELK1_CH/U_SLAVE_1ELK/Q[0]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]_net_1\);
    
    \U50_PATTERNS/ELINK_DINA_14[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119830, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_16, Q => 
        \U50_PATTERNS/ELINK_DINA_14[1]\);
    
    HIEFFPLA_INST_0_52588 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_9[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_10[1]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[0]\, Y => 
        HIEFFPLA_NET_0_117543);
    
    \U_EXEC_MASTER/USB_MASTER_EN/TERMCNT_FG60M\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117731, CLK => CLK60MHZ, CLR
         => P_MASTER_POR_B_c_27, Q => 
        \U_EXEC_MASTER/USB_MASTER_EN/TERMCNT_FG60M_net_1\);
    
    HIEFFPLA_INST_0_57580 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_5[5]\, B => 
        HIEFFPLA_NET_0_116639, S => HIEFFPLA_NET_0_117121, Y => 
        HIEFFPLA_NET_0_116656);
    
    \U50_PATTERNS/ELINK_ADDRA_6[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119962, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_4, Q => 
        \U50_PATTERNS/ELINK_ADDRA_6[5]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[12]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_WRD_40M_FIXED[12]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_32_0, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[12]_net_1\);
    
    \U_ELK6_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]\ : DFN1C0
      port map(D => \U_ELK6_CH/U_SLAVE_1ELK/Q[2]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]_net_1\);
    
    \U50_PATTERNS/ELINK_BLKA[7]/U1\ : DFN1P0
      port map(D => HIEFFPLA_NET_0_119918, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_19, Q => 
        \U50_PATTERNS/ELINK_BLKA[7]\);
    
    HIEFFPLA_INST_0_43771 : AND3A
      port map(A => HIEFFPLA_NET_0_119585, B => 
        HIEFFPLA_NET_0_119564, C => HIEFFPLA_NET_0_119597, Y => 
        HIEFFPLA_NET_0_119217);
    
    \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_4[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_116998, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_16_0, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_4[0]\);
    
    \U_ELK1_CH/U_ELK1_SERDAT_SOURCE/SERDAT[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118190, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_11, Q => 
        \U_ELK1_CH/ELK_TX_DAT[3]\);
    
    HIEFFPLA_INST_0_53694 : AND3
      port map(A => HIEFFPLA_NET_0_116708, B => 
        HIEFFPLA_NET_0_117360, C => HIEFFPLA_NET_0_117415, Y => 
        HIEFFPLA_NET_0_117371);
    
    HIEFFPLA_INST_0_51702 : MX2
      port map(A => \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[50]\, B
         => \U_MASTER_DES/PHASE_ADJ_160_L[4]\, S => 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM_0[4]_net_1\, Y => 
        HIEFFPLA_NET_0_117722);
    
    HIEFFPLA_INST_0_51517 : AX1E
      port map(A => \U_EXEC_MASTER/PRESCALE[1]\, B => 
        \U_EXEC_MASTER/PRESCALE[0]\, C => 
        \U_EXEC_MASTER/PRESCALE[2]\, Y => HIEFFPLA_NET_0_117756);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_13[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116247, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_1, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_13[3]\);
    
    HIEFFPLA_INST_0_57802 : NAND3A
      port map(A => HIEFFPLA_NET_0_116622, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_6[6]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_6[5]\, Y => 
        HIEFFPLA_NET_0_116618);
    
    HIEFFPLA_INST_0_44360 : MX2
      port map(A => \TFC_STOP_ADDR[2]\, B => 
        \U50_PATTERNS/U4B_REGCROSS/SAMP_TWO[2]_net_1\, S => 
        HIEFFPLA_NET_0_119135, Y => HIEFFPLA_NET_0_119131);
    
    \U_ELK5_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]\ : DFN1C0
      port map(D => \U_ELK5_CH/U_SLAVE_1ELK/Q[10]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]_net_1\);
    
    \U_ELK17_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]\ : DFN1C0
      port map(D => \U_ELK17_CH/U_SLAVE_1ELK/Q[0]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]_net_1\);
    
    \U_ELK11_CH/U_ELK1_SERDAT_SOURCE/SERDAT[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118596, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_0, Q => 
        \U_ELK11_CH/ELK_TX_DAT[2]\);
    
    HIEFFPLA_INST_0_52093 : MX2C
      port map(A => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[76]_net_1\, B => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[77]_net_1\, S => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[0]\, Y => 
        HIEFFPLA_NET_0_117638);
    
    HIEFFPLA_INST_0_44837 : NOR3B
      port map(A => HIEFFPLA_NET_0_119596, B => 
        \U50_PATTERNS/USB_RXF_B\, C => HIEFFPLA_NET_0_119037, Y
         => HIEFFPLA_NET_0_119038);
    
    \U50_PATTERNS/U111_PATT_ELINK_BLK/DPRT_512X9_SRAM_R0C0\ : 
        RAM4K9
      generic map(MEMORYFILE => "DPRT_512X9_SRAM_R0C0.mem")

      port map(ADDRA11 => AFLSDF_GND, ADDRA10 => AFLSDF_GND, 
        ADDRA9 => AFLSDF_GND, ADDRA8 => \GND\, ADDRA7 => 
        \U50_PATTERNS/ELINK_ADDRA_11[7]\, ADDRA6 => 
        \U50_PATTERNS/ELINK_ADDRA_11[6]\, ADDRA5 => 
        \U50_PATTERNS/ELINK_ADDRA_11[5]\, ADDRA4 => 
        \U50_PATTERNS/ELINK_ADDRA_11[4]\, ADDRA3 => 
        \U50_PATTERNS/ELINK_ADDRA_11[3]\, ADDRA2 => 
        \U50_PATTERNS/ELINK_ADDRA_11[2]\, ADDRA1 => 
        \U50_PATTERNS/ELINK_ADDRA_11[1]\, ADDRA0 => 
        \U50_PATTERNS/ELINK_ADDRA_11[0]\, ADDRB11 => AFLSDF_GND, 
        ADDRB10 => AFLSDF_GND, ADDRB9 => AFLSDF_GND, ADDRB8 => 
        \GND\, ADDRB7 => \ELKS_ADDRB[7]\, ADDRB6 => 
        \ELKS_ADDRB_0[6]\, ADDRB5 => \ELKS_ADDRB[5]\, ADDRB4 => 
        \ELKS_ADDRB_0[4]\, ADDRB3 => \ELKS_ADDRB[3]\, ADDRB2 => 
        \ELKS_ADDRB_0[2]\, ADDRB1 => \ELKS_ADDRB[1]\, ADDRB0 => 
        \ELKS_ADDRB[0]\, DINA8 => \GND\, DINA7 => 
        \U50_PATTERNS/ELINK_DINA_11[7]\, DINA6 => 
        \U50_PATTERNS/ELINK_DINA_11[6]\, DINA5 => 
        \U50_PATTERNS/ELINK_DINA_11[5]\, DINA4 => 
        \U50_PATTERNS/ELINK_DINA_11[4]\, DINA3 => 
        \U50_PATTERNS/ELINK_DINA_11[3]\, DINA2 => 
        \U50_PATTERNS/ELINK_DINA_11[2]\, DINA1 => 
        \U50_PATTERNS/ELINK_DINA_11[1]\, DINA0 => 
        \U50_PATTERNS/ELINK_DINA_11[0]\, DINB8 => \GND\, DINB7
         => \ELK_RX_SER_WORD_11[7]\, DINB6 => 
        \ELK_RX_SER_WORD_11[6]\, DINB5 => \ELK_RX_SER_WORD_11[5]\, 
        DINB4 => \ELK_RX_SER_WORD_11[4]\, DINB3 => 
        \ELK_RX_SER_WORD_11[3]\, DINB2 => \ELK_RX_SER_WORD_11[2]\, 
        DINB1 => \ELK_RX_SER_WORD_11[1]\, DINB0 => 
        \ELK_RX_SER_WORD_11[0]\, WIDTHA0 => \VCC\, WIDTHA1 => 
        \VCC\, WIDTHB0 => \VCC\, WIDTHB1 => \VCC\, PIPEA => \VCC\, 
        PIPEB => \VCC\, WMODEA => \GND\, WMODEB => \GND\, BLKA
         => \U50_PATTERNS/ELINK_BLKA[11]\, BLKB => 
        ELKS_RAM_BLKB_EN, WENA => \U50_PATTERNS/ELINK_RWA[11]\, 
        WENB => ELKS_RWB, CLKA => CLK60MHZ, CLKB => CLK_40M_GL, 
        RESET => P_USB_MASTER_EN_c_0, DOUTA8 => OPEN, DOUTA7 => 
        \U50_PATTERNS/ELINK_DOUTA_11[7]\, DOUTA6 => 
        \U50_PATTERNS/ELINK_DOUTA_11[6]\, DOUTA5 => 
        \U50_PATTERNS/ELINK_DOUTA_11[5]\, DOUTA4 => 
        \U50_PATTERNS/ELINK_DOUTA_11[4]\, DOUTA3 => 
        \U50_PATTERNS/ELINK_DOUTA_11[3]\, DOUTA2 => 
        \U50_PATTERNS/ELINK_DOUTA_11[2]\, DOUTA1 => 
        \U50_PATTERNS/ELINK_DOUTA_11[1]\, DOUTA0 => 
        \U50_PATTERNS/ELINK_DOUTA_11[0]\, DOUTB8 => OPEN, DOUTB7
         => \PATT_ELK_DAT_11[7]\, DOUTB6 => \PATT_ELK_DAT_11[6]\, 
        DOUTB5 => \PATT_ELK_DAT_11[5]\, DOUTB4 => 
        \PATT_ELK_DAT_11[4]\, DOUTB3 => \PATT_ELK_DAT_11[3]\, 
        DOUTB2 => \PATT_ELK_DAT_11[2]\, DOUTB1 => 
        \PATT_ELK_DAT_11[1]\, DOUTB0 => \PATT_ELK_DAT_11[0]\);
    
    HIEFFPLA_INST_0_43172 : AND3B
      port map(A => HIEFFPLA_NET_0_119352, B => 
        HIEFFPLA_NET_0_119411, C => HIEFFPLA_NET_0_119353, Y => 
        HIEFFPLA_NET_0_119355);
    
    \U_EXEC_MASTER/MPOR_SALT_B_3\ : DFI1P0
      port map(D => HIEFFPLA_NET_0_117781, CLK => CLK_40M_GL, PRE
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_2\, QN => 
        MASTER_SALT_POR_B_i_0_i_3);
    
    \U50_PATTERNS/ELINK_BLKA[13]/U1\ : DFN1P0
      port map(D => HIEFFPLA_NET_0_119931, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_20, Q => 
        \U50_PATTERNS/ELINK_BLKA[13]\);
    
    \U_ELK14_CH/U_SLAVE_1ELK/Q[9]\ : DFN1C0
      port map(D => \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/Q[9]_net_1\);
    
    HIEFFPLA_INST_0_56285 : NAND3C
      port map(A => HIEFFPLA_NET_0_116876, B => 
        HIEFFPLA_NET_0_116884, C => HIEFFPLA_NET_0_116892, Y => 
        HIEFFPLA_NET_0_116900);
    
    \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[0]\ : DFN1C0
      port map(D => 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[0]_net_1\);
    
    \U_ELK1_CH/U_SLAVE_1ELK/Q[1]\ : DFN1C0
      port map(D => \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/Q[1]_net_1\);
    
    HIEFFPLA_INST_0_43627 : AND2A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/SM_BANK_SEL[11]\, Y => 
        HIEFFPLA_NET_0_119263);
    
    \U_ELK12_CH/U_ELK1_CMD_TX/SER_OUT_RDEL\ : DFN1C0
      port map(D => \U_ELK12_CH/U_ELK1_CMD_TX/SER_OUT_RI_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_8, Q
         => \U_ELK12_CH/ELK_OUT_R\);
    
    \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[9]\ : DFN1C0
      port map(D => 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\);
    
    \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[8]\ : DFN1C0
      port map(D => \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\);
    
    \U200A_TFC/ADDR_POINTER[4]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120360, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_30, Q => \TFC_ADDRB[4]\);
    
    \U50_PATTERNS/U4A_REGCROSS/LOCAL_REG_VAL[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119148, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_17, Q => \TFC_STRT_ADDR[6]\);
    
    HIEFFPLA_INST_0_50858 : NAND2B
      port map(A => \OP_MODE_c_0[1]\, B => \PATT_ELK_DAT_8[2]\, Y
         => HIEFFPLA_NET_0_117876);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_5[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_115994, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_15, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_5[1]\);
    
    \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[2]\ : DFN1C0
      port map(D => 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[2]_net_1\);
    
    \U200B_ELINKS/GP_PG_SM[4]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120212, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_29, Q => 
        \U200B_ELINKS/GP_PG_SM[4]_net_1\);
    
    HIEFFPLA_INST_0_42897 : AND2
      port map(A => \U50_PATTERNS/REG_STATE[4]_net_1\, B => 
        \U50_PATTERNS/REG_STATE[3]_net_1\, Y => 
        HIEFFPLA_NET_0_119431);
    
    \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[5]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[3]_net_1\, CLK => 
        CCC_160M_ADJ, CLR => P_MASTER_POR_B_c_34_0, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[5]_net_1\);
    
    \U_ELK3_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0\ : DFN1C0
      port map(D => CLK_40M_GL, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_8, Q => 
        \U_ELK3_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0_net_1\);
    
    HIEFFPLA_INST_0_42889 : AND3B
      port map(A => \U50_PATTERNS/REG_STATE[1]_net_1\, B => 
        \U50_PATTERNS/REG_STATE[3]_net_1\, C => 
        \U50_PATTERNS/REG_STATE[4]_net_1\, Y => 
        HIEFFPLA_NET_0_119434);
    
    HIEFFPLA_INST_0_38338 : MX2
      port map(A => \U50_PATTERNS/ELINKS_STOP_ADDR_T[4]\, B => 
        \U50_PATTERNS/RD_USB_ADBUS[4]\, S => 
        HIEFFPLA_NET_0_119413, Y => HIEFFPLA_NET_0_120115);
    
    AFLSDF_INV_53 : INV
      port map(A => \U200A_TFC/RX_SER_WORD_2DEL[2]_net_1\, Y => 
        \AFLSDF_INV_53\);
    
    HIEFFPLA_INST_0_62556 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_7[0]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_8[0]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[0]\, Y => 
        HIEFFPLA_NET_0_115975);
    
    HIEFFPLA_INST_0_61232 : MX2
      port map(A => HIEFFPLA_NET_0_117166, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_20[4]\, S => 
        HIEFFPLA_NET_0_117141, Y => HIEFFPLA_NET_0_116156);
    
    \U_ELK9_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]\ : DFN1C0
      port map(D => \U_ELK9_CH/U_SLAVE_1ELK/Q[0]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]_net_1\);
    
    HIEFFPLA_INST_0_58184 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_11[1]\, B => 
        HIEFFPLA_NET_0_116677, S => HIEFFPLA_NET_0_117163, Y => 
        HIEFFPLA_NET_0_116553);
    
    HIEFFPLA_INST_0_53334 : AND2B
      port map(A => \BIT_OS_SEL[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_SEL[3]_net_1\, Y
         => HIEFFPLA_NET_0_117425);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_11[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116262, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_20, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_11[3]\);
    
    HIEFFPLA_INST_0_41921 : AO1A
      port map(A => \U50_PATTERNS/SM_BANK_SEL[0]\, B => 
        HIEFFPLA_NET_0_119240, C => \U50_PATTERNS/ELINK_RWA[11]\, 
        Y => HIEFFPLA_NET_0_119661);
    
    \U200A_TFC/LOC_STOP_ADDR[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120289, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_1, Q => \U200A_TFC/LOC_STOP_ADDR[1]\);
    
    HIEFFPLA_INST_0_61046 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_19[0]\, B => 
        HIEFFPLA_NET_0_117096, S => HIEFFPLA_NET_0_117170, Y => 
        HIEFFPLA_NET_0_116180);
    
    HIEFFPLA_INST_0_47571 : MX2
      port map(A => \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[0]_net_1\, 
        B => \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\, S => 
        \BIT_OS_SEL_2[2]\, Y => HIEFFPLA_NET_0_118474);
    
    \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[7]\ : DFN1C0
      port map(D => 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\);
    
    HIEFFPLA_INST_0_58503 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_31[3]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_15[3]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_3[4]_net_1\, Y
         => HIEFFPLA_NET_0_116513);
    
    HIEFFPLA_INST_0_43797 : AND3
      port map(A => HIEFFPLA_NET_0_119593, B => 
        \U50_PATTERNS/RD_USB_ADBUS[2]\, C => 
        \U50_PATTERNS/RD_USB_ADBUS[3]\, Y => 
        HIEFFPLA_NET_0_119212);
    
    \U_EXEC_MASTER/USB_MASTER_EN/T_CNT60M[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117741, CLK => CLK60MHZ, CLR
         => P_MASTER_POR_B_c_28, Q => 
        \U_EXEC_MASTER/USB_MASTER_EN/T_CNT60M[2]_net_1\);
    
    \U_ELK8_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]\ : DFN1C0
      port map(D => \U_ELK8_CH/U_SLAVE_1ELK/Q[4]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]_net_1\);
    
    \U_ELK4_CH/U_SLAVE_1ELK/RECD_SER_WORD[3]\ : DFN1C0
      port map(D => \U_ELK4_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[3]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_4[3]\);
    
    \U_ELK3_CH/U_SLAVE_1ELK/Q[7]\ : DFN1C0
      port map(D => \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/Q[7]_net_1\);
    
    HIEFFPLA_INST_0_37477 : MX2
      port map(A => \U200A_TFC/LOC_STRT_ADDR[4]\, B => 
        \TFC_STRT_ADDR[4]\, S => \U200A_TFC/GP_PG_SM_0[10]_net_1\, 
        Y => HIEFFPLA_NET_0_120278);
    
    \U200A_TFC/RX_SER_WORD_2DEL[2]\ : DFN1C0
      port map(D => \U200A_TFC/RX_SER_WORD_1DEL[2]_net_1\, CLK
         => CLK_40M_GL, CLR => P_MASTER_POR_B_c, Q => 
        \U200A_TFC/RX_SER_WORD_2DEL[2]_net_1\);
    
    HIEFFPLA_INST_0_45723 : AO1
      port map(A => HIEFFPLA_NET_0_119236, B => 
        \U50_PATTERNS/ELINK_DOUTA_0[3]\, C => 
        HIEFFPLA_NET_0_118785, Y => HIEFFPLA_NET_0_118858);
    
    \U_ELK3_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]\ : DFN1C0
      port map(D => \U_ELK3_CH/U_SLAVE_1ELK/Q[1]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]_net_1\);
    
    \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[12]\ : DFN1C0
      port map(D => \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\, 
        CLK => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\);
    
    HIEFFPLA_INST_0_37833 : AO1D
      port map(A => \OP_MODE_c[6]\, B => HIEFFPLA_NET_0_120190, C
         => HIEFFPLA_NET_0_120235, Y => HIEFFPLA_NET_0_120195);
    
    HIEFFPLA_INST_0_56643 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_0[1]\, B => 
        HIEFFPLA_NET_0_116799, S => HIEFFPLA_NET_0_117602, Y => 
        HIEFFPLA_NET_0_116823);
    
    HIEFFPLA_INST_0_55810 : MX2
      port map(A => HIEFFPLA_NET_0_116003, B => 
        HIEFFPLA_NET_0_116259, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[3]\, Y => 
        HIEFFPLA_NET_0_116987);
    
    HIEFFPLA_INST_0_41242 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_4[0]\, B => 
        HIEFFPLA_NET_0_119578, S => HIEFFPLA_NET_0_119284, Y => 
        HIEFFPLA_NET_0_119759);
    
    \U_ELK8_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]\ : DFN1C0
      port map(D => \U_ELK8_CH/U_SLAVE_1ELK/Q[12]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]_net_1\);
    
    HIEFFPLA_INST_0_53432 : MX2
      port map(A => HIEFFPLA_NET_0_117239, B => 
        HIEFFPLA_NET_0_117418, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[2]_net_1\, Y
         => HIEFFPLA_NET_0_117409);
    
    HIEFFPLA_INST_0_38024 : MX2
      port map(A => \U200B_ELINKS/LOC_STRT_ADDR[7]\, B => 
        \ELKS_STRT_ADDR[7]\, S => 
        \U200B_ELINKS/GP_PG_SM[10]_net_1\, Y => 
        HIEFFPLA_NET_0_120172);
    
    \U_ELK7_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]\ : DFN1C0
      port map(D => \U_ELK7_CH/U_SLAVE_1ELK/Q[14]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]_net_1\);
    
    \U50_PATTERNS/ELINK_DINA_8[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119726, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_18, Q => 
        \U50_PATTERNS/ELINK_DINA_8[1]\);
    
    HIEFFPLA_INST_0_50862 : AND2A
      port map(A => \OP_MODE_c_0[1]\, B => \PATT_ELK_DAT_8[6]\, Y
         => HIEFFPLA_NET_0_117872);
    
    HIEFFPLA_INST_0_43793 : AND3
      port map(A => HIEFFPLA_NET_0_119592, B => 
        \U50_PATTERNS/RD_USB_ADBUS[2]\, C => 
        \U50_PATTERNS/RD_USB_ADBUS[3]\, Y => 
        HIEFFPLA_NET_0_119213);
    
    HIEFFPLA_INST_0_43699 : NAND3C
      port map(A => HIEFFPLA_NET_0_119234, B => 
        HIEFFPLA_NET_0_119259, C => HIEFFPLA_NET_0_119287, Y => 
        HIEFFPLA_NET_0_119238);
    
    \U50_PATTERNS/REG_ADDR[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119526, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_10, Q => \U50_PATTERNS/REG_ADDR[7]\);
    
    \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[7]\ : DFN1C0
      port map(D => 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\);
    
    \U50_PATTERNS/REG_ADDR[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119533, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_10, Q => \U50_PATTERNS/REG_ADDR[0]\);
    
    HIEFFPLA_INST_0_58440 : MX2
      port map(A => HIEFFPLA_NET_0_116815, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_14[3]\, S => 
        HIEFFPLA_NET_0_117219, Y => HIEFFPLA_NET_0_116521);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_5[4]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116657, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_11, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_5[4]\);
    
    HIEFFPLA_INST_0_40118 : AOI1C
      port map(A => \U50_PATTERNS/ELINK_BLKA[17]\, B => 
        HIEFFPLA_NET_0_119233, C => HIEFFPLA_NET_0_119876, Y => 
        HIEFFPLA_NET_0_119900);
    
    \U50_PATTERNS/ELINK_DINA_2[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119772, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_9, Q => 
        \U50_PATTERNS/ELINK_DINA_2[3]\);
    
    HIEFFPLA_INST_0_48865 : NAND2B
      port map(A => \OP_MODE_c_5[1]\, B => \PATT_ELK_DAT_19[1]\, 
        Y => HIEFFPLA_NET_0_118237);
    
    HIEFFPLA_INST_0_43990 : MX2
      port map(A => \U50_PATTERNS/TFC_STOP_ADDR[1]\, B => 
        \U50_PATTERNS/TFC_STOP_ADDR_T[1]\, S => 
        HIEFFPLA_NET_0_119472, Y => HIEFFPLA_NET_0_119187);
    
    \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[14]\ : DFN1C0
      port map(D => \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\, 
        CLK => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[14]_net_1\);
    
    \U50_PATTERNS/SM_BANK_SEL[15]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119316, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_1_0, Q => 
        \U50_PATTERNS/SM_BANK_SEL[15]\);
    
    \U50_PATTERNS/ELINK_RWA[8]/U1\ : DFN1P0
      port map(D => HIEFFPLA_NET_0_119693, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_6, Q => \U50_PATTERNS/ELINK_RWA[8]\);
    
    HIEFFPLA_INST_0_41494 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_7[4]\, B => 
        HIEFFPLA_NET_0_119570, S => HIEFFPLA_NET_0_119289, Y => 
        HIEFFPLA_NET_0_119731);
    
    \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[14]\ : DFN1C0
      port map(D => \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[14]_net_1\);
    
    HIEFFPLA_INST_0_52316 : AND3B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[5]_net_1\, B => 
        HIEFFPLA_NET_0_117582, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[4]_net_1\, Y => 
        HIEFFPLA_NET_0_117583);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_18[4]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116186, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_8, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_18[4]\);
    
    \U50_PATTERNS/U4B_REGCROSS/SAMP_TWO[1]\ : DFN1C0
      port map(D => \U50_PATTERNS/U4B_REGCROSS/SAMP_ONE[1]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_29, Q => 
        \U50_PATTERNS/U4B_REGCROSS/SAMP_TWO[1]_net_1\);
    
    AFLSDF_INV_56 : INV
      port map(A => \U_ELK3_CH/U_DDR_ELK1/ELK_IN_DDR_R\, Y => 
        \AFLSDF_INV_56\);
    
    \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[2]\ : DFN1C0
      port map(D => \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\);
    
    HIEFFPLA_INST_0_40819 : MX2
      port map(A => HIEFFPLA_NET_0_119576, B => 
        \U50_PATTERNS/ELINK_DINA_17[1]\, S => 
        HIEFFPLA_NET_0_119260, Y => HIEFFPLA_NET_0_119806);
    
    HIEFFPLA_INST_0_42938 : AOI1A
      port map(A => HIEFFPLA_NET_0_119432, B => 
        HIEFFPLA_NET_0_119466, C => HIEFFPLA_NET_0_119403, Y => 
        HIEFFPLA_NET_0_119419);
    
    HIEFFPLA_INST_0_52866 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_19[2]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_20[2]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_1[0]\, Y => 
        HIEFFPLA_NET_0_117498);
    
    HIEFFPLA_INST_0_51837 : XA1
      port map(A => \U_MASTER_DES/U13A_ADJ_160M/BITCNT[0]\, B => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[1]\, C => 
        HIEFFPLA_NET_0_117674, Y => HIEFFPLA_NET_0_117680);
    
    HIEFFPLA_INST_0_43706 : AND2A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/SM_BANK_SEL[19]\, Y => 
        HIEFFPLA_NET_0_119236);
    
    HIEFFPLA_INST_0_47547 : MX2
      port map(A => HIEFFPLA_NET_0_118487, B => 
        HIEFFPLA_NET_0_118475, S => \BIT_OS_SEL_5[0]\, Y => 
        \U_ELK13_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[7]\);
    
    \U_ELK10_CH/U_SLAVE_1ELK/RECD_SER_WORD[3]\ : DFN1C0
      port map(D => \U_ELK10_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[3]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_10[3]\);
    
    HIEFFPLA_INST_0_58029 : AOI1A
      port map(A => HIEFFPLA_NET_0_116592, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_7[3]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_7[4]\, Y => 
        HIEFFPLA_NET_0_116575);
    
    HIEFFPLA_INST_0_43964 : MX2
      port map(A => HIEFFPLA_NET_0_119560, B => 
        \U50_PATTERNS/TFC_DINA[7]\, S => HIEFFPLA_NET_0_119294, Y
         => HIEFFPLA_NET_0_119190);
    
    HIEFFPLA_INST_0_56997 : AOI1A
      port map(A => HIEFFPLA_NET_0_116775, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_1[4]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_1[5]\, Y => 
        HIEFFPLA_NET_0_116757);
    
    \U50_PATTERNS/ELINK_DINA_1[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119783, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_7, Q => 
        \U50_PATTERNS/ELINK_DINA_1[0]\);
    
    \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_2S_3\ : DFN1C0
      port map(D => 
        \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_1S_net_1\, CLK
         => CLK60MHZ, CLR => P_MASTER_POR_B_c_0_0, Q => 
        P_USB_MASTER_EN_c_3);
    
    HIEFFPLA_INST_0_45458 : AO1
      port map(A => HIEFFPLA_NET_0_119250, B => 
        \U50_PATTERNS/ELINK_DOUTA_5[3]\, C => 
        HIEFFPLA_NET_0_118817, Y => HIEFFPLA_NET_0_118910);
    
    \U_ELK1_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL\ : DFN1C0
      port map(D => 
        \U_ELK1_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL_net_1\);
    
    HIEFFPLA_INST_0_43729 : NAND3C
      port map(A => \U50_PATTERNS/SM_BANK_SEL[0]\, B => 
        \U50_PATTERNS/SM_BANK_SEL[2]\, C => 
        \U50_PATTERNS/SM_BANK_SEL[1]\, Y => HIEFFPLA_NET_0_119229);
    
    \U_ELK10_CH/U_SLAVE_1ELK/Q[8]\ : DFN1C0
      port map(D => \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/Q[8]_net_1\);
    
    HIEFFPLA_INST_0_51715 : NAND2B
      port map(A => 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM[4]_net_1\, B => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[41]_net_1\, Y => 
        HIEFFPLA_NET_0_117711);
    
    \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[0]\ : DFN1C0
      port map(D => 
        \U_ELK8_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\);
    
    \U_ELK15_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U0\ : IOPADP_BI
      port map(N2PIN => 
        \U_ELK15_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2_N2P\, D => 
        \U_ELK15_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, E => 
        \U_ELK15_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET2\, PAD => 
        ELK15_DAT_P, Y => 
        \U_ELK15_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/TUNE_CLKPHASE[0]/U1\ : DFN1P0
      port map(D => HIEFFPLA_NET_0_115949, CLK => CLK_40M_GL, PRE
         => P_MASTER_POR_B_c_12, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/TUNE_CLKPHASE[0]\);
    
    HIEFFPLA_INST_0_60292 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_9[0]\, B => 
        HIEFFPLA_NET_0_116680, S => HIEFFPLA_NET_0_117130, Y => 
        HIEFFPLA_NET_0_116285);
    
    \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[12]\ : DFN1C0
      port map(D => 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]_net_1\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[12]_net_1\);
    
    \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[11]\ : DFN1C0
      port map(D => 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[11]_net_1\);
    
    \U50_PATTERNS/ELINK_DINA_18[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119793, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_21, Q => 
        \U50_PATTERNS/ELINK_DINA_18[6]\);
    
    \U50_PATTERNS/ELINK_BLKA[0]/U1\ : DFN1P0
      port map(D => HIEFFPLA_NET_0_119935, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_19, Q => 
        \U50_PATTERNS/ELINK_BLKA[0]\);
    
    \U200B_ELINKS/LOC_STOP_ADDR[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120186, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_7, Q => 
        \U200B_ELINKS/LOC_STOP_ADDR[1]\);
    
    HIEFFPLA_INST_0_59242 : MX2
      port map(A => HIEFFPLA_NET_0_116411, B => 
        HIEFFPLA_NET_0_116409, S => HIEFFPLA_NET_0_117366, Y => 
        HIEFFPLA_NET_0_116416);
    
    HIEFFPLA_INST_0_49339 : MX2
      port map(A => 
        \U_ELK2_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]_net_1\, B => 
        \U_ELK2_CH/ELK_TX_DAT[6]\, S => 
        \U_ELK2_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118154);
    
    HIEFFPLA_INST_0_62817 : MX2
      port map(A => HIEFFPLA_NET_0_115877, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/TUNE_CLKPHASE[3]\, S => 
        HIEFFPLA_NET_0_117102, Y => HIEFFPLA_NET_0_115942);
    
    HIEFFPLA_INST_0_59429 : MX2B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_26[3]\, B => 
        HIEFFPLA_NET_0_116774, S => HIEFFPLA_NET_0_117337, Y => 
        HIEFFPLA_NET_0_116395);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_6[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116313, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_2, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_6[1]\);
    
    \U50_PATTERNS/TFC_BLKA/U1\ : DFN1P0
      port map(D => HIEFFPLA_NET_0_119199, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_13, Q => \U50_PATTERNS/TFC_BLKA\);
    
    \U_ELK9_CH/U_ELK1_SERDAT_SOURCE/SERDAT[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117833, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_7, Q => 
        \U_ELK9_CH/ELK_TX_DAT[0]\);
    
    HIEFFPLA_INST_0_45221 : NAND3C
      port map(A => HIEFFPLA_NET_0_118741, B => 
        HIEFFPLA_NET_0_118920, C => HIEFFPLA_NET_0_118751, Y => 
        HIEFFPLA_NET_0_118963);
    
    \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[13]\ : DFN1C0
      port map(D => 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]_net_1\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[13]_net_1\);
    
    \U50_PATTERNS/U4B_REGCROSS/SAMP_TWO[4]\ : DFN1C0
      port map(D => \U50_PATTERNS/U4B_REGCROSS/SAMP_ONE[4]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_29, Q => 
        \U50_PATTERNS/U4B_REGCROSS/SAMP_TWO[4]_net_1\);
    
    HIEFFPLA_INST_0_57809 : NAND2B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_6[7]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_6[6]\, Y => 
        HIEFFPLA_NET_0_116616);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_6[7]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116625, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_12, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_6[7]\);
    
    \U_ELK6_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]\ : DFN1C0
      port map(D => \U_ELK6_CH/U_SLAVE_1ELK/Q[6]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]_net_1\);
    
    HIEFFPLA_INST_0_54714 : NAND3B
      port map(A => HIEFFPLA_NET_0_117238, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[0]_net_1\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[3]_net_1\, Y => 
        HIEFFPLA_NET_0_117219);
    
    \U50_PATTERNS/ELINK_ADDRA_4[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119978, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_2_0, Q => 
        \U50_PATTERNS/ELINK_ADDRA_4[5]\);
    
    HIEFFPLA_INST_0_44812 : NAND3C
      port map(A => HIEFFPLA_NET_0_119041, B => 
        HIEFFPLA_NET_0_119421, C => HIEFFPLA_NET_0_119588, Y => 
        HIEFFPLA_NET_0_119043);
    
    HIEFFPLA_INST_0_56766 : AO1
      port map(A => HIEFFPLA_NET_0_116813, B => 
        HIEFFPLA_NET_0_117354, C => HIEFFPLA_NET_0_117406, Y => 
        HIEFFPLA_NET_0_116803);
    
    \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_2S_12\ : DFN1C0
      port map(D => 
        \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_1S_0_net_1\, CLK
         => CLK60MHZ, CLR => \U_EXEC_MASTER/P_MASTER_POR_B_c_0\, 
        Q => P_USB_MASTER_EN_c_12);
    
    HIEFFPLA_INST_0_54567 : NAND2A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[4]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[2]_net_1\, Y => 
        HIEFFPLA_NET_0_117246);
    
    HIEFFPLA_INST_0_48868 : AND2A
      port map(A => \OP_MODE_c_6[1]\, B => \PATT_ELK_DAT_19[4]\, 
        Y => HIEFFPLA_NET_0_118234);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_6[8]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116624, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_12, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_6[8]\);
    
    HIEFFPLA_INST_0_51852 : AND2
      port map(A => HIEFFPLA_NET_0_117673, B => 
        HIEFFPLA_NET_0_117674, Y => HIEFFPLA_NET_0_117677);
    
    HIEFFPLA_INST_0_59262 : NOR3A
      port map(A => HIEFFPLA_NET_0_116407, B => 
        HIEFFPLA_NET_0_116410, C => HIEFFPLA_NET_0_116412, Y => 
        HIEFFPLA_NET_0_116413);
    
    \U_ELK1_CH/U_SLAVE_1ELK/Q[4]\ : DFN1C0
      port map(D => \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/Q[4]_net_1\);
    
    HIEFFPLA_INST_0_39047 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_16[5]\, B => 
        HIEFFPLA_NET_0_119518, S => HIEFFPLA_NET_0_119257, Y => 
        HIEFFPLA_NET_0_120034);
    
    HIEFFPLA_INST_0_40783 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_16[5]\, B => 
        HIEFFPLA_NET_0_119567, S => HIEFFPLA_NET_0_119257, Y => 
        HIEFFPLA_NET_0_119810);
    
    HIEFFPLA_INST_0_43291 : MX2
      port map(A => \U50_PATTERNS/SI_CNT[2]\, B => 
        HIEFFPLA_NET_0_119325, S => HIEFFPLA_NET_0_119439, Y => 
        HIEFFPLA_NET_0_119332);
    
    \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[10]\ : DFN1C0
      port map(D => \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\);
    
    HIEFFPLA_INST_0_51041 : MX2
      port map(A => HIEFFPLA_NET_0_117844, B => 
        HIEFFPLA_NET_0_117864, S => \BIT_OS_SEL_3[1]\, Y => 
        HIEFFPLA_NET_0_117846);
    
    HIEFFPLA_INST_0_42673 : AO1D
      port map(A => \U50_PATTERNS/REG_STATE_0[5]_net_1\, B => 
        HIEFFPLA_NET_0_119368, C => HIEFFPLA_NET_0_119402, Y => 
        HIEFFPLA_NET_0_119486);
    
    \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[11]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[9]_net_1\, CLK => 
        CCC_160M_ADJ, CLR => P_MASTER_POR_B_c_26, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[11]_net_1\);
    
    HIEFFPLA_INST_0_37752 : AOI1
      port map(A => \OP_MODE_c[6]\, B => HIEFFPLA_NET_0_120234, C
         => HIEFFPLA_NET_0_120215, Y => HIEFFPLA_NET_0_120216);
    
    \U62_TS_OE_BUF/\\\\TRIBUFF_F_24U[0]\\\\/U0/U0\ : IOPAD_TRI_U
      port map(D => 
        \U62_TS_OE_BUF/\\\\TRIBUFF_F_24U[0]\\\\/U0/NET1\, E => 
        \U62_TS_OE_BUF/\\\\TRIBUFF_F_24U[0]\\\\/U0/NET2\, PAD => 
        USB_OE_B);
    
    HIEFFPLA_INST_0_37809 : AND3
      port map(A => HIEFFPLA_NET_0_120228, B => 
        \U200B_ELINKS/GP_PG_SM[8]_net_1\, C => \OP_MODE[4]\, Y
         => HIEFFPLA_NET_0_120203);
    
    \U_ELK9_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]\ : DFN1C0
      port map(D => \U_ELK9_CH/U_SLAVE_1ELK/Q[6]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]_net_1\);
    
    \U_ELK12_CH/ELK_IN_F\ : DFN1C0
      port map(D => \U_ELK12_CH/ELK_IN_DDR_F\, CLK => 
        CCC_160M_ADJ, CLR => DEV_RST_B_c, Q => 
        \U_ELK12_CH/ELK_IN_F_net_1\);
    
    HIEFFPLA_INST_0_47306 : MX2
      port map(A => HIEFFPLA_NET_0_118519, B => 
        HIEFFPLA_NET_0_118530, S => \BIT_OS_SEL_4[1]\, Y => 
        HIEFFPLA_NET_0_118521);
    
    \U_ELK10_CH/U_SLAVE_1ELK/Q[14]\ : DFN1C0
      port map(D => \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[14]_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/Q[14]_net_1\);
    
    \U50_PATTERNS/U4D_REGCROSS/SAMP_TWO[2]\ : DFN1C0
      port map(D => \U50_PATTERNS/U4D_REGCROSS/SAMP_ONE[2]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_30, Q => 
        \U50_PATTERNS/U4D_REGCROSS/SAMP_TWO[2]_net_1\);
    
    HIEFFPLA_INST_0_57077 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_2[7]\, B => 
        HIEFFPLA_NET_0_116728, S => HIEFFPLA_NET_0_117601, Y => 
        HIEFFPLA_NET_0_116748);
    
    \U50_PATTERNS/ELINK_ADDRA_11[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120075, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_2, Q => 
        \U50_PATTERNS/ELINK_ADDRA_11[4]\);
    
    HIEFFPLA_INST_0_42232 : AND3A
      port map(A => HIEFFPLA_NET_0_119559, B => 
        \U50_PATTERNS/RD_USB_ADBUS[5]\, C => 
        \U50_PATTERNS/RD_USB_ADBUS[4]\, Y => 
        HIEFFPLA_NET_0_119597);
    
    HIEFFPLA_INST_0_46110 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_19[4]\, C => 
        \U50_PATTERNS/SM_BANK_SEL[0]\, Y => HIEFFPLA_NET_0_118763);
    
    HIEFFPLA_INST_0_37668 : AND3B
      port map(A => HIEFFPLA_NET_0_120147, B => 
        \U200B_ELINKS/GP_PG_SM[10]_net_1\, C => 
        HIEFFPLA_NET_0_120220, Y => HIEFFPLA_NET_0_120236);
    
    HIEFFPLA_INST_0_44094 : MX2
      port map(A => \U50_PATTERNS/TFC_STOP_ADDR_T[6]\, B => 
        \U50_PATTERNS/RD_USB_ADBUS[6]\, S => 
        HIEFFPLA_NET_0_119492, Y => HIEFFPLA_NET_0_119174);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_19[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116177, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_11, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_19[3]\);
    
    HIEFFPLA_INST_0_62914 : MX2
      port map(A => HIEFFPLA_NET_0_115893, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[1]\, S => 
        HIEFFPLA_NET_0_117073, Y => HIEFFPLA_NET_0_115929);
    
    HIEFFPLA_INST_0_63108 : AND2B
      port map(A => HIEFFPLA_NET_0_117078, B => 
        HIEFFPLA_NET_0_115880, Y => HIEFFPLA_NET_0_115886);
    
    HIEFFPLA_INST_0_46443 : AND3C
      port map(A => HIEFFPLA_NET_0_118672, B => 
        HIEFFPLA_NET_0_118676, C => HIEFFPLA_NET_0_118681, Y => 
        HIEFFPLA_NET_0_118689);
    
    \U_ELK5_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]\ : DFN1C0
      port map(D => \U_ELK5_CH/U_SLAVE_1ELK/Q[2]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]_net_1\);
    
    HIEFFPLA_INST_0_45145 : MX2
      port map(A => HIEFFPLA_NET_0_118968, B => 
        \U50_PATTERNS/WR_USB_ADBUS[7]\, S => 
        HIEFFPLA_NET_0_119486, Y => HIEFFPLA_NET_0_118978);
    
    HIEFFPLA_INST_0_56937 : OA1A
      port map(A => HIEFFPLA_NET_0_116776, B => 
        HIEFFPLA_NET_0_116594, C => HIEFFPLA_NET_0_116679, Y => 
        HIEFFPLA_NET_0_116770);
    
    HIEFFPLA_INST_0_111286 : NAND3C
      port map(A => HIEFFPLA_NET_0_116806, B => 
        HIEFFPLA_NET_0_116742, C => HIEFFPLA_NET_0_116687, Y => 
        HIEFFPLA_NET_0_115843);
    
    \U_ELK0_SERDAT_SOURCE/SERDAT[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118658, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_10, Q => \ELK0_TX_DAT[2]\);
    
    \U_ELK2_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL\ : DFN1C0
      port map(D => 
        \U_ELK2_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL_net_1\);
    
    HIEFFPLA_INST_0_60450 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_11[1]\, B => 
        HIEFFPLA_NET_0_117114, S => HIEFFPLA_NET_0_117348, Y => 
        HIEFFPLA_NET_0_116264);
    
    HIEFFPLA_INST_0_51924 : MX2A
      port map(A => HIEFFPLA_NET_0_117657, B => 
        HIEFFPLA_NET_0_117656, S => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[5]\, Y => 
        HIEFFPLA_NET_0_117665);
    
    HIEFFPLA_INST_0_43431 : MX2
      port map(A => \U50_PATTERNS/SM_BANK_SEL[19]\, B => 
        HIEFFPLA_NET_0_119218, S => HIEFFPLA_NET_0_118691, Y => 
        HIEFFPLA_NET_0_119312);
    
    HIEFFPLA_INST_0_47897 : MX2
      port map(A => HIEFFPLA_NET_0_118406, B => 
        HIEFFPLA_NET_0_118403, S => \BIT_OS_SEL_2[1]\, Y => 
        HIEFFPLA_NET_0_118407);
    
    \U_EXEC_MASTER/SYNC_BRD_RST_BI\ : DFI1P0
      port map(D => \U_EXEC_MASTER/DEV_RST_1B_i\, CLK => 
        CCC_160M_FXD, PRE => DEV_RST_B_c, QN => 
        \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i\);
    
    \U200A_TFC/LOC_STOP_ADDR[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120290, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_1, Q => \U200A_TFC/LOC_STOP_ADDR[0]\);
    
    \U50_PATTERNS/ELINK_ADDRA_0[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120089, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_18, Q => 
        \U50_PATTERNS/ELINK_ADDRA_0[6]\);
    
    HIEFFPLA_INST_0_46768 : MX2
      port map(A => HIEFFPLA_NET_0_118625, B => 
        HIEFFPLA_NET_0_118622, S => \BIT_OS_SEL_0[0]\, Y => 
        \U_ELK10_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[3]\);
    
    HIEFFPLA_INST_0_43919 : MX2
      port map(A => HIEFFPLA_NET_0_119575, B => 
        \U50_PATTERNS/TFC_DINA[2]\, S => HIEFFPLA_NET_0_119294, Y
         => HIEFFPLA_NET_0_119195);
    
    HIEFFPLA_INST_0_37226 : NAND3C
      port map(A => \U200A_TFC/GP_PG_SM[0]_net_1\, B => 
        \U200A_TFC/GP_PG_SM[1]_net_1\, C => HIEFFPLA_NET_0_120325, 
        Y => HIEFFPLA_NET_0_120320);
    
    \U_ELK11_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]\ : DFN1C0
      port map(D => \U_ELK11_CH/U_SLAVE_1ELK/Q[9]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]_net_1\);
    
    HIEFFPLA_INST_0_62834 : AOI1D
      port map(A => HIEFFPLA_NET_0_115944, B => 
        HIEFFPLA_NET_0_115943, C => HIEFFPLA_NET_0_117104, Y => 
        HIEFFPLA_NET_0_115939);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_23[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116118, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_6, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_23[2]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_8[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116291, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_5, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_8[2]\);
    
    \U_ELK6_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117976, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_9, Q => 
        \U_ELK6_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]_net_1\);
    
    HIEFFPLA_INST_0_53078 : MX2
      port map(A => HIEFFPLA_NET_0_117556, B => 
        HIEFFPLA_NET_0_117552, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[2]\, Y => 
        HIEFFPLA_NET_0_117468);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_5[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116320, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_1, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_5[2]\);
    
    \U50_PATTERNS/ELINK_ADDRA_11[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120072, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_2, Q => 
        \U50_PATTERNS/ELINK_ADDRA_11[7]\);
    
    HIEFFPLA_INST_0_60552 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_12[4]\, B => 
        HIEFFPLA_NET_0_117100, S => HIEFFPLA_NET_0_117133, Y => 
        HIEFFPLA_NET_0_116251);
    
    HIEFFPLA_INST_0_41143 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_2[5]\, B => 
        HIEFFPLA_NET_0_119567, S => HIEFFPLA_NET_0_119278, Y => 
        HIEFFPLA_NET_0_119770);
    
    \U_ELK5_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U1\ : IOBI_ID_OD_EB
      port map(DR => \U_ELK5_CH/ELK_OUT_R\, DF => 
        \U_ELK5_CH/ELK_OUT_F\, CLR => \GND\, E => \AFLSDF_INV_42\, 
        ICLK => CCC_160M_ADJ, OCLK => CCC_160M_FXD, YIN => 
        \U_ELK5_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\, DOUT => 
        \U_ELK5_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, EOUT => 
        \U_ELK5_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET2\, YR => 
        \U_ELK5_CH/ELK_IN_DDR_R\, YF => \U_ELK5_CH/ELK_IN_DDR_F\);
    
    HIEFFPLA_INST_0_61406 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_22[0]\, B => 
        HIEFFPLA_NET_0_117190, S => HIEFFPLA_NET_0_117080, Y => 
        HIEFFPLA_NET_0_116130);
    
    \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[11]\ : DFN1C0
      port map(D => 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]_net_1\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[11]_net_1\);
    
    HIEFFPLA_INST_0_44547 : AND2
      port map(A => \U50_PATTERNS/U4D_REGCROSS/DELCNT[0]_net_1\, 
        B => \U50_PATTERNS/U4D_REGCROSS/DELCNT[1]_net_1\, Y => 
        HIEFFPLA_NET_0_119093);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_4[8]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116688, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_9, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_4[8]\);
    
    HIEFFPLA_INST_0_45922 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_15[2]\, C => 
        \U50_PATTERNS/SM_BANK_SEL[4]\, Y => HIEFFPLA_NET_0_118810);
    
    HIEFFPLA_INST_0_40495 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_12[5]\, B => 
        HIEFFPLA_NET_0_119567, S => HIEFFPLA_NET_0_119295, Y => 
        HIEFFPLA_NET_0_119842);
    
    \U_ELK2_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]\ : DFN1C0
      port map(D => \U_ELK2_CH/U_SLAVE_1ELK/Q[1]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_13[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116541, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_12, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_13[1]\);
    
    \U_ELK11_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]\ : DFN1C0
      port map(D => \U_ELK11_CH/U_SLAVE_1ELK/Q[11]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]_net_1\);
    
    HIEFFPLA_INST_0_63244 : NAND2B
      port map(A => \OP_MODE_c_0[1]\, B => \PATT_TFC_DAT[7]\, Y
         => \U_TFC_SERDAT_SOURCE/N_SERDAT[7]\);
    
    HIEFFPLA_INST_0_58662 : MX2
      port map(A => HIEFFPLA_NET_0_116486, B => 
        HIEFFPLA_NET_0_116484, S => HIEFFPLA_NET_0_117231, Y => 
        HIEFFPLA_NET_0_116491);
    
    HIEFFPLA_INST_0_53379 : MX2
      port map(A => HIEFFPLA_NET_0_116451, B => 
        HIEFFPLA_NET_0_116372, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[3]_net_1\, Y
         => HIEFFPLA_NET_0_117418);
    
    HIEFFPLA_INST_0_46808 : MX2
      port map(A => HIEFFPLA_NET_0_118609, B => 
        HIEFFPLA_NET_0_118621, S => \BIT_OS_SEL_5[1]\, Y => 
        HIEFFPLA_NET_0_118611);
    
    \U_ELK11_CH/ELK_IN_R\ : DFN1C0
      port map(D => \U_ELK11_CH/ELK_IN_DDR_R\, CLK => 
        CCC_160M_ADJ, CLR => DEV_RST_B_c, Q => 
        \U_ELK11_CH/ELK_IN_R_net_1\);
    
    HIEFFPLA_INST_0_45756 : AO1
      port map(A => HIEFFPLA_NET_0_119263, B => 
        \U50_PATTERNS/ELINK_DOUTA_8[2]\, C => 
        HIEFFPLA_NET_0_118768, Y => HIEFFPLA_NET_0_118851);
    
    HIEFFPLA_INST_0_40855 : MX2
      port map(A => HIEFFPLA_NET_0_119567, B => 
        \U50_PATTERNS/ELINK_DINA_17[5]\, S => 
        HIEFFPLA_NET_0_119260, Y => HIEFFPLA_NET_0_119802);
    
    HIEFFPLA_INST_0_45872 : AO1
      port map(A => HIEFFPLA_NET_0_119283, B => 
        \U50_PATTERNS/ELINK_DOUTA_13[5]\, C => 
        HIEFFPLA_NET_0_118776, Y => HIEFFPLA_NET_0_118823);
    
    HIEFFPLA_INST_0_61337 : MX2
      port map(A => HIEFFPLA_NET_0_117166, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_21[4]\, S => 
        HIEFFPLA_NET_0_117144, Y => HIEFFPLA_NET_0_116141);
    
    HIEFFPLA_INST_0_51408 : AND2
      port map(A => \U_EXEC_MASTER/DEL_CNT[3]\, B => 
        \U_EXEC_MASTER/DEL_CNT[2]\, Y => HIEFFPLA_NET_0_117783);
    
    HIEFFPLA_INST_0_44102 : MX2
      port map(A => \U50_PATTERNS/TFC_STOP_ADDR_T[7]\, B => 
        \U50_PATTERNS/RD_USB_ADBUS[7]\, S => 
        HIEFFPLA_NET_0_119492, Y => HIEFFPLA_NET_0_119173);
    
    \U_ELK7_CH/U_SLAVE_1ELK/Q[4]\ : DFN1C0
      port map(D => \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/Q[4]_net_1\);
    
    \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[0]\ : DFN1C0
      port map(D => 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[0]_net_1\);
    
    HIEFFPLA_INST_0_56459 : AOI1D
      port map(A => HIEFFPLA_NET_0_117432, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_SEL[3]_net_1\, C
         => \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[3]_net_1\, Y
         => HIEFFPLA_NET_0_116861);
    
    HIEFFPLA_INST_0_54357 : MX2
      port map(A => HIEFFPLA_NET_0_116444, B => 
        HIEFFPLA_NET_0_116351, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_2[3]_net_1\, Y
         => HIEFFPLA_NET_0_117276);
    
    \U_ELK16_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118382, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_14, Q => 
        \U_ELK16_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]_net_1\);
    
    HIEFFPLA_INST_0_57889 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_7[2]\, B => 
        HIEFFPLA_NET_0_116582, S => HIEFFPLA_NET_0_117113, Y => 
        HIEFFPLA_NET_0_116601);
    
    HIEFFPLA_INST_0_59785 : AO1C
      port map(A => HIEFFPLA_NET_0_117328, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_30[2]\, C => 
        HIEFFPLA_NET_0_117357, Y => HIEFFPLA_NET_0_116348);
    
    HIEFFPLA_INST_0_47917 : MX2
      port map(A => HIEFFPLA_NET_0_118405, B => 
        HIEFFPLA_NET_0_118401, S => \BIT_OS_SEL_2[1]\, Y => 
        HIEFFPLA_NET_0_118404);
    
    HIEFFPLA_INST_0_62622 : MX2
      port map(A => HIEFFPLA_NET_0_117100, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_8[4]\, S => 
        HIEFFPLA_NET_0_117153, Y => HIEFFPLA_NET_0_115966);
    
    \U50_PATTERNS/U4C_REGCROSS/DELCNT[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119094, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_28, Q => 
        \U50_PATTERNS/U4C_REGCROSS/DELCNT[1]_net_1\);
    
    HIEFFPLA_INST_0_39227 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_19[1]\, B => 
        HIEFFPLA_NET_0_119523, S => HIEFFPLA_NET_0_119293, Y => 
        HIEFFPLA_NET_0_120014);
    
    HIEFFPLA_INST_0_39218 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_19[0]\, B => 
        HIEFFPLA_NET_0_119524, S => HIEFFPLA_NET_0_119293, Y => 
        HIEFFPLA_NET_0_120015);
    
    \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[9]\ : DFN1C0
      port map(D => \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\);
    
    \U_ELK16_CH/U_SLAVE_1ELK/Q[11]\ : DFN1C0
      port map(D => \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/Q[11]_net_1\);
    
    \U_ELK13_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U3\ : IOBI_ID_OD_EB
      port map(DR => \U_ELK13_CH/ELK_OUT_R\, DF => 
        \U_ELK13_CH/ELK_OUT_F\, CLR => \GND\, E => 
        \AFLSDF_INV_21\, ICLK => CCC_160M_ADJ, OCLK => 
        CCC_160M_FXD, YIN => 
        \U_ELK13_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\, DOUT => 
        OPEN, EOUT => 
        \U_ELK13_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET3\, YR => OPEN, 
        YF => OPEN);
    
    HIEFFPLA_INST_0_42994 : AND3A
      port map(A => \U50_PATTERNS/REG_STATE[4]_net_1\, B => 
        HIEFFPLA_NET_0_119017, C => HIEFFPLA_NET_0_119370, Y => 
        HIEFFPLA_NET_0_119406);
    
    HIEFFPLA_INST_0_37706 : AND3B
      port map(A => \U200B_ELINKS/GP_PG_SM[9]_net_1\, B => 
        \U200B_ELINKS/GP_PG_SM[1]_net_1\, C => 
        HIEFFPLA_NET_0_120233, Y => HIEFFPLA_NET_0_120224);
    
    \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_2S_21\ : DFN1C0
      port map(D => 
        \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_1S_0_net_1\, CLK
         => CLK60MHZ, CLR => \U_EXEC_MASTER/P_MASTER_POR_B_c_0\, 
        Q => P_USB_MASTER_EN_c_21);
    
    HIEFFPLA_INST_0_60129 : NAND3A
      port map(A => HIEFFPLA_NET_0_117211, B => 
        HIEFFPLA_NET_0_116620, C => HIEFFPLA_NET_0_116649, Y => 
        HIEFFPLA_NET_0_116306);
    
    HIEFFPLA_INST_0_60702 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_14[4]\, B => 
        HIEFFPLA_NET_0_117166, S => HIEFFPLA_NET_0_117228, Y => 
        HIEFFPLA_NET_0_116231);
    
    HIEFFPLA_INST_0_58880 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_20[3]\, B => 
        HIEFFPLA_NET_0_116457, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_1[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116464);
    
    \U_MASTER_DES/U13C_MASTER_DESER/ARB_WRD_40M_FIXED[11]\ : 
        DFN1C0
      port map(D => \U_MASTER_DES/U13C_MASTER_DESER/Q[11]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_28, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_WRD_40M_FIXED[11]_net_1\);
    
    HIEFFPLA_INST_0_111643 : MX2B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[0]_net_1\, B => 
        \OP_MODE_c[5]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_0[8]_net_1\, Y => 
        HIEFFPLA_NET_0_115837);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_31[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116017, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_10, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_31[3]\);
    
    HIEFFPLA_INST_0_48124 : NAND2B
      port map(A => \OP_MODE_c_2[1]\, B => \PATT_ELK_DAT_16[7]\, 
        Y => HIEFFPLA_NET_0_118366);
    
    \U_ELK7_CH/U_SLAVE_1ELK/Q[8]\ : DFN1C0
      port map(D => \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/Q[8]_net_1\);
    
    HIEFFPLA_INST_0_53224 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_CLKPHASE[2]\, B => 
        HIEFFPLA_NET_0_117445, S => HIEFFPLA_NET_0_117111, Y => 
        HIEFFPLA_NET_0_117450);
    
    HIEFFPLA_INST_0_52454 : MX2
      port map(A => HIEFFPLA_NET_0_117513, B => 
        HIEFFPLA_NET_0_117509, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[3]\, Y => 
        HIEFFPLA_NET_0_117561);
    
    \U_ELK5_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]\ : DFN1C0
      port map(D => \U_ELK5_CH/U_SLAVE_1ELK/Q[13]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/MAX_CNT[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_116952, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_16, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/MAX_CNT[2]\);
    
    \U_EXEC_MASTER/MPOR_B_28\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117787, CLK => CLK_40M_GL, CLR
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_0\, Q => 
        P_MASTER_POR_B_c_28);
    
    \U50_PATTERNS/ELINK_ADDRA_0[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120092, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_18, Q => 
        \U50_PATTERNS/ELINK_ADDRA_0[3]\);
    
    HIEFFPLA_INST_0_55115 : AOI1D
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[6]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[8]_net_1\, C => 
        HIEFFPLA_NET_0_116740, Y => HIEFFPLA_NET_0_117119);
    
    \U_ELK7_CH/U_ELK1_SERDAT_SOURCE/SERDAT[6]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117917, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_3, Q => 
        \U_ELK7_CH/ELK_TX_DAT[6]\);
    
    HIEFFPLA_INST_0_61706 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_25[0]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_26[0]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_4[0]\, Y => 
        HIEFFPLA_NET_0_116090);
    
    HIEFFPLA_INST_0_59972 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_4[2]\, B => 
        HIEFFPLA_NET_0_116324, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_2[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116327);
    
    HIEFFPLA_INST_0_54039 : MX2
      port map(A => HIEFFPLA_NET_0_116122, B => 
        HIEFFPLA_NET_0_116025, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[3]_net_1\, Y
         => HIEFFPLA_NET_0_117316);
    
    HIEFFPLA_INST_0_53215 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_CLKPHASE[1]\, B => 
        HIEFFPLA_NET_0_117446, S => HIEFFPLA_NET_0_117111, Y => 
        HIEFFPLA_NET_0_117451);
    
    HIEFFPLA_INST_0_45325 : AO1A
      port map(A => HIEFFPLA_NET_0_118831, B => 
        \U50_PATTERNS/SM_BANK_SEL[5]\, C => HIEFFPLA_NET_0_118939, 
        Y => HIEFFPLA_NET_0_118940);
    
    \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[1]\ : DFN1C0
      port map(D => 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[1]_net_1\);
    
    HIEFFPLA_INST_0_52031 : MX2
      port map(A => HIEFFPLA_NET_0_117635, B => 
        HIEFFPLA_NET_0_117634, S => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[3]\, Y => 
        HIEFFPLA_NET_0_117648);
    
    \U200A_TFC/ADDR_POINTER[7]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120354, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_30, Q => \TFC_ADDRB[7]\);
    
    HIEFFPLA_INST_0_58564 : AND2A
      port map(A => HIEFFPLA_NET_0_117215, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_16[0]\, Y => 
        HIEFFPLA_NET_0_116504);
    
    \U_ELK16_CH/U_SLAVE_1ELK/RECD_SER_WORD[1]\ : DFN1C0
      port map(D => \U_ELK16_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[1]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_16[1]\);
    
    HIEFFPLA_INST_0_60588 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_13[3]\, B => 
        HIEFFPLA_NET_0_117186, S => HIEFFPLA_NET_0_117137, Y => 
        HIEFFPLA_NET_0_116247);
    
    \U50_PATTERNS/OP_MODE[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119616, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_15, Q => \U50_PATTERNS/OP_MODE[1]\);
    
    HIEFFPLA_INST_0_54765 : NAND3B
      port map(A => HIEFFPLA_NET_0_117245, B => 
        HIEFFPLA_NET_0_117252, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[1]_net_1\, Y => 
        HIEFFPLA_NET_0_117206);
    
    HIEFFPLA_INST_0_39245 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_19[3]\, B => 
        HIEFFPLA_NET_0_119520, S => HIEFFPLA_NET_0_119293, Y => 
        HIEFFPLA_NET_0_120012);
    
    \U50_PATTERNS/U115_PATT_ELINK_BLK/DPRT_512X9_SRAM_R0C0\ : 
        RAM4K9
      generic map(MEMORYFILE => "DPRT_512X9_SRAM_R0C0.mem")

      port map(ADDRA11 => AFLSDF_GND, ADDRA10 => AFLSDF_GND, 
        ADDRA9 => AFLSDF_GND, ADDRA8 => \GND\, ADDRA7 => 
        \U50_PATTERNS/ELINK_ADDRA_15[7]\, ADDRA6 => 
        \U50_PATTERNS/ELINK_ADDRA_15[6]\, ADDRA5 => 
        \U50_PATTERNS/ELINK_ADDRA_15[5]\, ADDRA4 => 
        \U50_PATTERNS/ELINK_ADDRA_15[4]\, ADDRA3 => 
        \U50_PATTERNS/ELINK_ADDRA_15[3]\, ADDRA2 => 
        \U50_PATTERNS/ELINK_ADDRA_15[2]\, ADDRA1 => 
        \U50_PATTERNS/ELINK_ADDRA_15[1]\, ADDRA0 => 
        \U50_PATTERNS/ELINK_ADDRA_15[0]\, ADDRB11 => AFLSDF_GND, 
        ADDRB10 => AFLSDF_GND, ADDRB9 => AFLSDF_GND, ADDRB8 => 
        \GND\, ADDRB7 => \ELKS_ADDRB[7]\, ADDRB6 => 
        \ELKS_ADDRB[6]\, ADDRB5 => \ELKS_ADDRB[5]\, ADDRB4 => 
        \ELKS_ADDRB[4]\, ADDRB3 => \ELKS_ADDRB[3]\, ADDRB2 => 
        \ELKS_ADDRB[2]\, ADDRB1 => \ELKS_ADDRB[1]\, ADDRB0 => 
        \ELKS_ADDRB[0]\, DINA8 => \GND\, DINA7 => 
        \U50_PATTERNS/ELINK_DINA_15[7]\, DINA6 => 
        \U50_PATTERNS/ELINK_DINA_15[6]\, DINA5 => 
        \U50_PATTERNS/ELINK_DINA_15[5]\, DINA4 => 
        \U50_PATTERNS/ELINK_DINA_15[4]\, DINA3 => 
        \U50_PATTERNS/ELINK_DINA_15[3]\, DINA2 => 
        \U50_PATTERNS/ELINK_DINA_15[2]\, DINA1 => 
        \U50_PATTERNS/ELINK_DINA_15[1]\, DINA0 => 
        \U50_PATTERNS/ELINK_DINA_15[0]\, DINB8 => \GND\, DINB7
         => \ELK_RX_SER_WORD_15[7]\, DINB6 => 
        \ELK_RX_SER_WORD_15[6]\, DINB5 => \ELK_RX_SER_WORD_15[5]\, 
        DINB4 => \ELK_RX_SER_WORD_15[4]\, DINB3 => 
        \ELK_RX_SER_WORD_15[3]\, DINB2 => \ELK_RX_SER_WORD_15[2]\, 
        DINB1 => \ELK_RX_SER_WORD_15[1]\, DINB0 => 
        \ELK_RX_SER_WORD_15[0]\, WIDTHA0 => \VCC\, WIDTHA1 => 
        \VCC\, WIDTHB0 => \VCC\, WIDTHB1 => \VCC\, PIPEA => \VCC\, 
        PIPEB => \VCC\, WMODEA => \GND\, WMODEB => \GND\, BLKA
         => \U50_PATTERNS/ELINK_BLKA[15]\, BLKB => 
        ELKS_RAM_BLKB_EN, WENA => \U50_PATTERNS/ELINK_RWA[15]\, 
        WENB => ELKS_RWB, CLKA => CLK60MHZ, CLKB => CLK_40M_GL, 
        RESET => P_USB_MASTER_EN_c_0, DOUTA8 => OPEN, DOUTA7 => 
        \U50_PATTERNS/ELINK_DOUTA_15[7]\, DOUTA6 => 
        \U50_PATTERNS/ELINK_DOUTA_15[6]\, DOUTA5 => 
        \U50_PATTERNS/ELINK_DOUTA_15[5]\, DOUTA4 => 
        \U50_PATTERNS/ELINK_DOUTA_15[4]\, DOUTA3 => 
        \U50_PATTERNS/ELINK_DOUTA_15[3]\, DOUTA2 => 
        \U50_PATTERNS/ELINK_DOUTA_15[2]\, DOUTA1 => 
        \U50_PATTERNS/ELINK_DOUTA_15[1]\, DOUTA0 => 
        \U50_PATTERNS/ELINK_DOUTA_15[0]\, DOUTB8 => OPEN, DOUTB7
         => \PATT_ELK_DAT_15[7]\, DOUTB6 => \PATT_ELK_DAT_15[6]\, 
        DOUTB5 => \PATT_ELK_DAT_15[5]\, DOUTB4 => 
        \PATT_ELK_DAT_15[4]\, DOUTB3 => \PATT_ELK_DAT_15[3]\, 
        DOUTB2 => \PATT_ELK_DAT_15[2]\, DOUTB1 => 
        \PATT_ELK_DAT_15[1]\, DOUTB0 => \PATT_ELK_DAT_15[0]\);
    
    \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[11]\ : DFN1C0
      port map(D => 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[11]_net_1\);
    
    HIEFFPLA_INST_0_52099 : MX2C
      port map(A => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[78]_net_1\, B => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[79]_net_1\, S => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[0]\, Y => 
        HIEFFPLA_NET_0_117637);
    
    \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[6]\ : DFN1C0
      port map(D => 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\);
    
    \U_ELK13_CH/U_SLAVE_1ELK/Q[2]\ : DFN1C0
      port map(D => \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/Q[2]_net_1\);
    
    \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[0]\ : DFN1C0
      port map(D => 
        \U_ELK14_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\);
    
    HIEFFPLA_INST_0_43705 : NAND3C
      port map(A => HIEFFPLA_NET_0_119234, B => 
        HIEFFPLA_NET_0_119259, C => HIEFFPLA_NET_0_119286, Y => 
        HIEFFPLA_NET_0_119237);
    
    \U_MASTER_DES/U13C_MASTER_DESER/Q[6]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[6]_net_1\, CLK => 
        CCC_160M_FXD, CLR => P_MASTER_POR_B_c_34, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/Q[6]_net_1\);
    
    \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[14]\ : DFN1C0
      port map(D => 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[14]_net_1\);
    
    HIEFFPLA_INST_0_53843 : NAND3C
      port map(A => HIEFFPLA_NET_0_117370, B => 
        HIEFFPLA_NET_0_117310, C => HIEFFPLA_NET_0_117407, Y => 
        HIEFFPLA_NET_0_117344);
    
    HIEFFPLA_INST_0_50222 : MX2
      port map(A => HIEFFPLA_NET_0_117995, B => 
        HIEFFPLA_NET_0_117993, S => \BIT_OS_SEL_6[1]\, Y => 
        HIEFFPLA_NET_0_117990);
    
    \U_ELK7_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL\ : DFN1C0
      port map(D => 
        \U_ELK7_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL_net_1\);
    
    HIEFFPLA_INST_0_51630 : MX2
      port map(A => 
        \U_EXEC_MASTER/USB_MASTER_EN/CNT_EN_60M2S_net_1\, B => 
        \U_EXEC_MASTER/USB_MASTER_EN/T_CNT60M[4]_net_1\, S => 
        HIEFFPLA_NET_0_117753, Y => HIEFFPLA_NET_0_117733);
    
    HIEFFPLA_INST_0_45384 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_7[6]\, C => 
        \U50_PATTERNS/SM_BANK_SEL[12]\, Y => 
        HIEFFPLA_NET_0_118924);
    
    HIEFFPLA_INST_0_48720 : MX2
      port map(A => HIEFFPLA_NET_0_118266, B => 
        HIEFFPLA_NET_0_118263, S => \BIT_OS_SEL_1[1]\, Y => 
        HIEFFPLA_NET_0_118261);
    
    HIEFFPLA_INST_0_43395 : MX2
      port map(A => \U50_PATTERNS/SM_BANK_SEL[15]\, B => 
        HIEFFPLA_NET_0_119222, S => HIEFFPLA_NET_0_118691, Y => 
        HIEFFPLA_NET_0_119316);
    
    \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[10]\ : DFN1C0
      port map(D => \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\);
    
    \U50_PATTERNS/ELINK_DINA_6[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119738, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_16, Q => 
        \U50_PATTERNS/ELINK_DINA_6[5]\);
    
    HIEFFPLA_INST_0_43616 : AOI1B
      port map(A => \U50_PATTERNS/REG_STATE[2]_net_1\, B => 
        \U50_PATTERNS/REG_STATE[1]_net_1\, C => 
        \U50_PATTERNS/SM_BANK_SEL[20]\, Y => 
        HIEFFPLA_NET_0_119267);
    
    \U_ELK9_CH/U_ELK1_CMD_TX/SER_OUT_RDEL\ : DFN1C0
      port map(D => \U_ELK9_CH/U_ELK1_CMD_TX/SER_OUT_RI_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_13, Q
         => \U_ELK9_CH/ELK_OUT_R\);
    
    HIEFFPLA_INST_0_43310 : NAND3
      port map(A => \U50_PATTERNS/SI_CNT[2]\, B => 
        \U50_PATTERNS/SI_CNT[1]\, C => \U50_PATTERNS/SI_CNT[0]\, 
        Y => HIEFFPLA_NET_0_119330);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_24[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116433, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_18, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_24[1]\);
    
    HIEFFPLA_INST_0_38561 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_0[7]\, B => 
        HIEFFPLA_NET_0_119516, S => HIEFFPLA_NET_0_119272, Y => 
        HIEFFPLA_NET_0_120088);
    
    HIEFFPLA_INST_0_51816 : NAND2B
      port map(A => \U_MASTER_DES/U13A_ADJ_160M/BITCNT[4]\, B => 
        HIEFFPLA_NET_0_117685, Y => HIEFFPLA_NET_0_117688);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_4[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116328, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_20, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_4[1]\);
    
    \U50_PATTERNS/ELINK_RWA[9]/U1\ : DFN1P0
      port map(D => HIEFFPLA_NET_0_119692, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_6, Q => \U50_PATTERNS/ELINK_RWA[9]\);
    
    \U200B_ELINKS/RX_SER_WORD_1DEL[0]\ : DFN1C0
      port map(D => \ELK_RX_SER_WORD_0[0]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_23, Q => 
        \U200B_ELINKS/RX_SER_WORD_1DEL[0]_net_1\);
    
    HIEFFPLA_INST_0_53989 : MX2
      port map(A => HIEFFPLA_NET_0_117227, B => 
        HIEFFPLA_NET_0_117358, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[2]_net_1\, Y
         => HIEFFPLA_NET_0_117323);
    
    HIEFFPLA_INST_0_48097 : AND2
      port map(A => \U_ELK16_CH/ELK_TX_DAT[1]\, B => 
        \U_ELK16_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118378);
    
    HIEFFPLA_INST_0_51298 : MX2
      port map(A => HIEFFPLA_NET_0_117810, B => 
        HIEFFPLA_NET_0_117798, S => \BIT_OS_SEL_5[1]\, Y => 
        HIEFFPLA_NET_0_117800);
    
    HIEFFPLA_INST_0_44622 : NAND3C
      port map(A => HIEFFPLA_NET_0_119079, B => 
        HIEFFPLA_NET_0_119080, C => HIEFFPLA_NET_0_119081, Y => 
        HIEFFPLA_NET_0_119082);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_3[6]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116719, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_7, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_3[6]\);
    
    HIEFFPLA_INST_0_61289 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_4[2]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_20[2]\, S
         => \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_5[4]_net_1\, 
        Y => HIEFFPLA_NET_0_116147);
    
    HIEFFPLA_INST_0_46843 : MX2
      port map(A => 
        \U_ELK11_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]_net_1\, B => 
        \U_ELK11_CH/ELK_TX_DAT[4]\, S => 
        \U_ELK11_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118605);
    
    \U50_PATTERNS/U3_USB_DAT_BUS/_BIBUF_F_24U[2]_/U0/U1\ : 
        IOBI_IRC_OB_EB
      port map(D => \U50_PATTERNS/WR_USB_ADBUS[2]\, CLR => 
        \AFLSDF_INV_6\, E => \U50_PATTERNS/TrienAux\, ICLK => 
        CLK60MHZ, YIN => 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[2]\\\\/U0/NET3\, 
        DOUT => 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[2]\\\\/U0/NET1\, 
        EOUT => 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[2]\\\\/U0/NET2\, 
        Y => \U50_PATTERNS/RD_USB_ADBUS[2]\);
    
    HIEFFPLA_INST_0_46529 : AOI1A
      port map(A => HIEFFPLA_NET_0_119571, B => 
        HIEFFPLA_NET_0_119587, C => 
        \U50_PATTERNS/WR_XFER_TYPE[1]_net_1\, Y => 
        HIEFFPLA_NET_0_118671);
    
    \U_ELK17_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118334, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_17, Q => 
        \U_ELK17_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]_net_1\);
    
    \U200B_ELINKS/LOC_STOP_ADDR[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120180, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_7, Q => 
        \U200B_ELINKS/LOC_STOP_ADDR[7]\);
    
    \U_ELK1_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]\ : DFN1C0
      port map(D => \U_ELK1_CH/U_SLAVE_1ELK/Q[3]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]_net_1\);
    
    \U50_PATTERNS/ELINK_ADDRA_0[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120088, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_19, Q => 
        \U50_PATTERNS/ELINK_ADDRA_0[7]\);
    
    HIEFFPLA_INST_0_42133 : MX2
      port map(A => \U50_PATTERNS/OP_MODE[5]\, B => 
        \U50_PATTERNS/OP_MODE_T[5]\, S => HIEFFPLA_NET_0_119472, 
        Y => HIEFFPLA_NET_0_119612);
    
    HIEFFPLA_INST_0_43760 : AND3C
      port map(A => HIEFFPLA_NET_0_119590, B => 
        HIEFFPLA_NET_0_119596, C => HIEFFPLA_NET_0_119559, Y => 
        HIEFFPLA_NET_0_119221);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_0[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116572, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_15, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_0[0]\);
    
    HIEFFPLA_INST_0_45785 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/SM_BANK_SEL[19]\, C => 
        \U50_PATTERNS/ELINK_DOUTA_0[2]\, Y => 
        HIEFFPLA_NET_0_118843);
    
    \U_ELK7_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117930, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_14, Q => 
        \U_ELK7_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]_net_1\);
    
    HIEFFPLA_INST_0_50393 : MX2
      port map(A => \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[1]_net_1\, B
         => \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\, S => 
        \BIT_OS_SEL_5[2]\, Y => HIEFFPLA_NET_0_117957);
    
    HIEFFPLA_INST_0_47939 : MX2
      port map(A => \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\, 
        B => \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[11]_net_1\, S => 
        \BIT_OS_SEL_1[2]\, Y => HIEFFPLA_NET_0_118401);
    
    \U50_PATTERNS/SM_BANK_SEL[11]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119320, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_1_0, Q => 
        \U50_PATTERNS/SM_BANK_SEL[11]\);
    
    HIEFFPLA_INST_0_52932 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_31[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_0[1]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_3[0]\, Y => 
        HIEFFPLA_NET_0_117487);
    
    HIEFFPLA_INST_0_42887 : AO1B
      port map(A => \U50_PATTERNS/REG_STATE[2]_net_1\, B => 
        \U50_PATTERNS/REG_STATE[1]_net_1\, C => 
        \U50_PATTERNS/REG_STATE[5]_net_1\, Y => 
        HIEFFPLA_NET_0_119435);
    
    \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[2]\ : DFN1C0
      port map(D => 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[2]_net_1\);
    
    \U50_PATTERNS/U100_PATT_ELINK_BLK/DPRT_512X9_SRAM_R0C0\ : 
        RAM4K9
      generic map(MEMORYFILE => "DPRT_512X9_SRAM_R0C0.mem")

      port map(ADDRA11 => AFLSDF_GND, ADDRA10 => AFLSDF_GND, 
        ADDRA9 => AFLSDF_GND, ADDRA8 => \GND\, ADDRA7 => 
        \U50_PATTERNS/ELINK_ADDRA_0[7]\, ADDRA6 => 
        \U50_PATTERNS/ELINK_ADDRA_0[6]\, ADDRA5 => 
        \U50_PATTERNS/ELINK_ADDRA_0[5]\, ADDRA4 => 
        \U50_PATTERNS/ELINK_ADDRA_0[4]\, ADDRA3 => 
        \U50_PATTERNS/ELINK_ADDRA_0[3]\, ADDRA2 => 
        \U50_PATTERNS/ELINK_ADDRA_0[2]\, ADDRA1 => 
        \U50_PATTERNS/ELINK_ADDRA_0[1]\, ADDRA0 => 
        \U50_PATTERNS/ELINK_ADDRA_0[0]\, ADDRB11 => AFLSDF_GND, 
        ADDRB10 => AFLSDF_GND, ADDRB9 => AFLSDF_GND, ADDRB8 => 
        \GND\, ADDRB7 => \ELKS_ADDRB[7]\, ADDRB6 => 
        \ELKS_ADDRB[6]\, ADDRB5 => \ELKS_ADDRB[5]\, ADDRB4 => 
        \ELKS_ADDRB[4]\, ADDRB3 => \ELKS_ADDRB[3]\, ADDRB2 => 
        \ELKS_ADDRB[2]\, ADDRB1 => \ELKS_ADDRB[1]\, ADDRB0 => 
        \ELKS_ADDRB[0]\, DINA8 => \GND\, DINA7 => 
        \U50_PATTERNS/ELINK_DINA_0[7]\, DINA6 => 
        \U50_PATTERNS/ELINK_DINA_0[6]\, DINA5 => 
        \U50_PATTERNS/ELINK_DINA_0[5]\, DINA4 => 
        \U50_PATTERNS/ELINK_DINA_0[4]\, DINA3 => 
        \U50_PATTERNS/ELINK_DINA_0[3]\, DINA2 => 
        \U50_PATTERNS/ELINK_DINA_0[2]\, DINA1 => 
        \U50_PATTERNS/ELINK_DINA_0[1]\, DINA0 => 
        \U50_PATTERNS/ELINK_DINA_0[0]\, DINB8 => \GND\, DINB7 => 
        \ELK_RX_SER_WORD_0[7]\, DINB6 => \ELK_RX_SER_WORD_0[6]\, 
        DINB5 => \ELK_RX_SER_WORD_0[5]\, DINB4 => 
        \ELK_RX_SER_WORD_0[4]\, DINB3 => \ELK_RX_SER_WORD_0[3]\, 
        DINB2 => \ELK_RX_SER_WORD_0[2]\, DINB1 => 
        \ELK_RX_SER_WORD_0[1]\, DINB0 => \ELK_RX_SER_WORD_0[0]\, 
        WIDTHA0 => \VCC\, WIDTHA1 => \VCC\, WIDTHB0 => \VCC\, 
        WIDTHB1 => \VCC\, PIPEA => \VCC\, PIPEB => \VCC\, WMODEA
         => \GND\, WMODEB => \GND\, BLKA => 
        \U50_PATTERNS/ELINK_BLKA[0]\, BLKB => ELKS_RAM_BLKB_EN, 
        WENA => \U50_PATTERNS/ELINK_RWA[0]\, WENB => ELKS_RWB, 
        CLKA => CLK60MHZ, CLKB => CLK_40M_GL, RESET => 
        P_USB_MASTER_EN_c_0, DOUTA8 => OPEN, DOUTA7 => 
        \U50_PATTERNS/ELINK_DOUTA_0[7]\, DOUTA6 => 
        \U50_PATTERNS/ELINK_DOUTA_0[6]\, DOUTA5 => 
        \U50_PATTERNS/ELINK_DOUTA_0[5]\, DOUTA4 => 
        \U50_PATTERNS/ELINK_DOUTA_0[4]\, DOUTA3 => 
        \U50_PATTERNS/ELINK_DOUTA_0[3]\, DOUTA2 => 
        \U50_PATTERNS/ELINK_DOUTA_0[2]\, DOUTA1 => 
        \U50_PATTERNS/ELINK_DOUTA_0[1]\, DOUTA0 => 
        \U50_PATTERNS/ELINK_DOUTA_0[0]\, DOUTB8 => OPEN, DOUTB7
         => \PATT_ELK_DAT_0[7]\, DOUTB6 => \PATT_ELK_DAT_0[6]\, 
        DOUTB5 => \PATT_ELK_DAT_0[5]\, DOUTB4 => 
        \PATT_ELK_DAT_0[4]\, DOUTB3 => \PATT_ELK_DAT_0[3]\, 
        DOUTB2 => \PATT_ELK_DAT_0[2]\, DOUTB1 => 
        \PATT_ELK_DAT_0[1]\, DOUTB0 => \PATT_ELK_DAT_0[0]\);
    
    \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[5]\ : DFN1C0
      port map(D => 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_0[7]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116817, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_3, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_0[7]\);
    
    \U_ELK18_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118291, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_3, Q => 
        \U_ELK18_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]_net_1\);
    
    \U_ELK17_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U1\ : IOBI_ID_OD_EB
      port map(DR => \U_ELK17_CH/ELK_OUT_R\, DF => 
        \U_ELK17_CH/ELK_OUT_F\, CLR => \GND\, E => 
        \AFLSDF_INV_28\, ICLK => CCC_160M_ADJ, OCLK => 
        CCC_160M_FXD, YIN => 
        \U_ELK17_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\, DOUT => 
        \U_ELK17_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, EOUT => 
        \U_ELK17_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET2\, YR => 
        \U_ELK17_CH/ELK_IN_DDR_R\, YF => 
        \U_ELK17_CH/ELK_IN_DDR_F\);
    
    \U50_PATTERNS/ELINK_ADDRA_7[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119957, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_6, Q => 
        \U50_PATTERNS/ELINK_ADDRA_7[2]\);
    
    \U50_PATTERNS/ELINKS_STRT_ADDR[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120109, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_17, Q => 
        \U50_PATTERNS/ELINKS_STRT_ADDR[2]\);
    
    \U_ELK14_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]\ : DFN1C0
      port map(D => \U_ELK14_CH/U_SLAVE_1ELK/Q[7]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]_net_1\);
    
    HIEFFPLA_INST_0_61997 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_12[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_28[1]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_3[4]_net_1\, Y
         => HIEFFPLA_NET_0_116049);
    
    HIEFFPLA_INST_0_51111 : AND2A
      port map(A => \OP_MODE_c_3[1]\, B => \PATT_ELK_DAT_9[6]\, Y
         => HIEFFPLA_NET_0_117827);
    
    \U_ELK8_CH/U_SLAVE_1ELK/Q[14]\ : DFN1C0
      port map(D => \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[14]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/Q[14]_net_1\);
    
    HIEFFPLA_INST_0_59307 : MX2B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_25[3]\, B => 
        HIEFFPLA_NET_0_116774, S => HIEFFPLA_NET_0_117394, Y => 
        HIEFFPLA_NET_0_116407);
    
    \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_2S_1_0\ : DFN1C0
      port map(D => 
        \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_1S_0_net_1\, CLK
         => CLK60MHZ, CLR => P_MASTER_POR_B_c_0_0, Q => 
        P_USB_MASTER_EN_c_1_0);
    
    HIEFFPLA_INST_0_58628 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_1[2]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_17[2]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[4]_net_1\, Y
         => HIEFFPLA_NET_0_116496);
    
    \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[13]\ : DFN1C0
      port map(D => 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]_net_1\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[13]_net_1\);
    
    HIEFFPLA_INST_0_49654 : MX2
      port map(A => HIEFFPLA_NET_0_118087, B => 
        HIEFFPLA_NET_0_118083, S => \BIT_OS_SEL[1]\, Y => 
        HIEFFPLA_NET_0_118090);
    
    HIEFFPLA_INST_0_37786 : AOI1D
      port map(A => HIEFFPLA_NET_0_120192, B => 
        HIEFFPLA_NET_0_120200, C => HIEFFPLA_NET_0_120218, Y => 
        HIEFFPLA_NET_0_120207);
    
    \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[11]\ : DFN1C0
      port map(D => \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\);
    
    \U_ELK0_CMD_TX/SER_CMD_WORD_F[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118669, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_17, Q => 
        \U_ELK0_CMD_TX/SER_CMD_WORD_F[0]_net_1\);
    
    \U_ELK17_CH/U_ELK1_SERDAT_SOURCE/SERDAT[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118325, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_11, Q => 
        \U_ELK17_CH/ELK_TX_DAT[3]\);
    
    HIEFFPLA_INST_0_161275 : DFN1C0
      port map(D => \U_ELK0_CMD_TX/SER_CMD_WORD_F[1]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_17, Q
         => HIEFFPLA_NET_0_161280);
    
    HIEFFPLA_INST_0_39713 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_6[7]\, B => 
        HIEFFPLA_NET_0_119516, S => HIEFFPLA_NET_0_119258, Y => 
        HIEFFPLA_NET_0_119960);
    
    \U_ELK8_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL\ : DFN1C0
      port map(D => 
        \U_ELK8_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL_net_1\);
    
    \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[6]\ : DFN1C0
      port map(D => \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\);
    
    \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[3]\ : DFN1C0
      port map(D => \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\);
    
    HIEFFPLA_INST_0_61469 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_6[4]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_22[4]\, S
         => \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_5[4]_net_1\, 
        Y => HIEFFPLA_NET_0_116122);
    
    \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[6]\ : DFN1C0
      port map(D => 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_19[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116480, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_20, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_19[1]\);
    
    HIEFFPLA_INST_0_55267 : AND3C
      port map(A => HIEFFPLA_NET_0_117102, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[3]_net_1\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[2]_net_1\, Y => 
        HIEFFPLA_NET_0_117073);
    
    \EXTCLK_40MHZ_pad/U0/U0\ : IOPAD_TRI_U
      port map(D => \EXTCLK_40MHZ_pad/U0/NET1\, E => 
        \EXTCLK_40MHZ_pad/U0/NET2\, PAD => EXTCLK_40MHZ);
    
    \U_REFCLKBUF/\\\\BIBUF_LVDS[0]\\\\/U0/U2\ : IOPADN_BI
      port map(DB => \U_REFCLKBUF/\\\\BIBUF_LVDS[0]\\\\/U0/NET1\, 
        E => \U_REFCLKBUF/\\\\BIBUF_LVDS[0]\\\\/U0/NET3\, PAD => 
        REF_CLK_0N, N2POUT => 
        \U_REFCLKBUF/\\\\BIBUF_LVDS[0]\\\\/U0/U2_N2P\);
    
    \U_ELK19_CH/U_SLAVE_1ELK/Q[14]\ : DFN1C0
      port map(D => \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[14]_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/Q[14]_net_1\);
    
    HIEFFPLA_INST_0_113037 : AO13
      port map(A => HIEFFPLA_NET_0_115812, B => 
        \U200B_ELINKS/LOC_STOP_ADDR[6]\, C => \ELKS_ADDRB[6]\, Y
         => HIEFFPLA_NET_0_115820);
    
    \U_ELK6_CH/U_ELK1_CMD_TX/SER_OUT_FDEL\ : DFN1C0
      port map(D => \U_ELK6_CH/U_ELK1_CMD_TX/SER_OUT_FI_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_1, Q
         => \U_ELK6_CH/ELK_OUT_F\);
    
    AFLSDF_INV_34 : INV
      port map(A => DCB_SALT_SEL_c, Y => \AFLSDF_INV_34\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_0[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116571, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_15, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_0[1]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_SEL_3[0]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_BIT_OS_VAL[0]\, CLK
         => CLK_40M_GL, CLR => P_MASTER_POR_B_c_27_0, Q => 
        \BIT_OS_SEL_3[0]\);
    
    HIEFFPLA_INST_0_57057 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_2[5]\, B => 
        HIEFFPLA_NET_0_116730, S => HIEFFPLA_NET_0_117601, Y => 
        HIEFFPLA_NET_0_116750);
    
    \U_ELK3_CH/U_ELK1_SERDAT_SOURCE/SERDAT[7]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118096, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_15, Q => 
        \U_ELK3_CH/ELK_TX_DAT[7]\);
    
    HIEFFPLA_INST_0_45850 : NAND2A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_15[0]\, Y => 
        HIEFFPLA_NET_0_118828);
    
    HIEFFPLA_INST_0_63062 : XA1B
      port map(A => HIEFFPLA_NET_0_115884, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[10]\, C => 
        HIEFFPLA_NET_0_117078, Y => HIEFFPLA_NET_0_115898);
    
    HIEFFPLA_INST_0_55199 : AND3B
      port map(A => HIEFFPLA_NET_0_117252, B => 
        HIEFFPLA_NET_0_117237, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[6]_net_1\, Y => 
        HIEFFPLA_NET_0_117095);
    
    HIEFFPLA_INST_0_48119 : NAND2B
      port map(A => \OP_MODE_c_2[1]\, B => \PATT_ELK_DAT_16[2]\, 
        Y => HIEFFPLA_NET_0_118371);
    
    \U_ELK6_CH/U_ELK1_SERDAT_SOURCE/SERDAT[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117967, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_1, Q => 
        \U_ELK6_CH/ELK_TX_DAT[1]\);
    
    \U50_PATTERNS/ELINK_DINA_14[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119831, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_16, Q => 
        \U50_PATTERNS/ELINK_DINA_14[0]\);
    
    HIEFFPLA_INST_0_40846 : MX2
      port map(A => HIEFFPLA_NET_0_119570, B => 
        \U50_PATTERNS/ELINK_DINA_17[4]\, S => 
        HIEFFPLA_NET_0_119260, Y => HIEFFPLA_NET_0_119803);
    
    \U_ELK17_CH/U_SLAVE_1ELK/Q[0]\ : DFN1C0
      port map(D => \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/Q[0]_net_1\);
    
    \U50_PATTERNS/U4E_REGCROSS/SAMP_ONE[2]\ : DFN1C0
      port map(D => \U50_PATTERNS/OP_MODE[2]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c, Q => 
        \U50_PATTERNS/U4E_REGCROSS/SAMP_ONE[2]_net_1\);
    
    HIEFFPLA_INST_0_56244 : AND2
      port map(A => DCB_SALT_SEL_c, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/RECD_SER_WORD[5]_net_1\, 
        Y => \ELK_RX_SER_WORD_0[5]\);
    
    HIEFFPLA_INST_0_53404 : MX2
      port map(A => HIEFFPLA_NET_0_116221, B => 
        HIEFFPLA_NET_0_116115, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[3]_net_1\, Y
         => HIEFFPLA_NET_0_117413);
    
    HIEFFPLA_INST_0_41161 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_2[7]\, B => 
        HIEFFPLA_NET_0_119560, S => HIEFFPLA_NET_0_119278, Y => 
        HIEFFPLA_NET_0_119768);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_7[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116303, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_3, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_7[0]\);
    
    HIEFFPLA_INST_0_45354 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_18[5]\, C => 
        \U50_PATTERNS/SM_BANK_SEL[1]\, Y => HIEFFPLA_NET_0_118932);
    
    HIEFFPLA_INST_0_55210 : AND2A
      port map(A => HIEFFPLA_NET_0_117210, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[6]_net_1\, Y => 
        HIEFFPLA_NET_0_117089);
    
    HIEFFPLA_INST_0_45264 : AO1
      port map(A => HIEFFPLA_NET_0_119263, B => 
        \U50_PATTERNS/ELINK_DOUTA_8[3]\, C => 
        HIEFFPLA_NET_0_118842, Y => HIEFFPLA_NET_0_118955);
    
    HIEFFPLA_INST_0_50931 : MX2
      port map(A => \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\, B
         => \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\, S => 
        \BIT_OS_SEL_3[2]\, Y => HIEFFPLA_NET_0_117861);
    
    \U_ELK19_CH/U_ELK1_CMD_TX/SER_OUT_FI\ : DFN1C0
      port map(D => 
        \U_ELK19_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_0, Q => 
        \U_ELK19_CH/U_ELK1_CMD_TX/SER_OUT_FI_net_1\);
    
    HIEFFPLA_INST_0_54954 : AND2A
      port map(A => HIEFFPLA_NET_0_117216, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_3[6]_net_1\, Y => 
        HIEFFPLA_NET_0_117158);
    
    HIEFFPLA_INST_0_40774 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_16[4]\, B => 
        HIEFFPLA_NET_0_119570, S => HIEFFPLA_NET_0_119257, Y => 
        HIEFFPLA_NET_0_119811);
    
    HIEFFPLA_INST_0_56236 : AND2
      port map(A => DCB_SALT_SEL_c, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/RECD_SER_WORD[1]_net_1\, 
        Y => \ELK_RX_SER_WORD_0[1]\);
    
    HIEFFPLA_INST_0_46704 : MX2
      port map(A => HIEFFPLA_NET_0_118620, B => 
        HIEFFPLA_NET_0_118633, S => \BIT_OS_SEL_5[1]\, Y => 
        HIEFFPLA_NET_0_118625);
    
    \U_ELK19_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]\ : DFN1C0
      port map(D => \U_ELK19_CH/U_SLAVE_1ELK/Q[3]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]_net_1\);
    
    HIEFFPLA_INST_0_50013 : MX2
      port map(A => HIEFFPLA_NET_0_118043, B => 
        HIEFFPLA_NET_0_118042, S => \BIT_OS_SEL_0[0]\, Y => 
        \U_ELK4_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[4]\);
    
    \U_ELK4_CH/U_ELK1_SERDAT_SOURCE/SERDAT[6]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118052, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_16, Q => 
        \U_ELK4_CH/ELK_TX_DAT[6]\);
    
    HIEFFPLA_INST_0_52974 : MX2
      port map(A => HIEFFPLA_NET_0_117469, B => 
        HIEFFPLA_NET_0_117465, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[4]\, Y => 
        HIEFFPLA_NET_0_117481);
    
    HIEFFPLA_INST_0_43422 : MX2
      port map(A => \U50_PATTERNS/SM_BANK_SEL[18]\, B => 
        HIEFFPLA_NET_0_119219, S => HIEFFPLA_NET_0_118691, Y => 
        HIEFFPLA_NET_0_119313);
    
    HIEFFPLA_INST_0_38134 : AND3
      port map(A => HIEFFPLA_NET_0_120145, B => \ELKS_ADDRB[3]\, 
        C => \ELKS_ADDRB[2]\, Y => HIEFFPLA_NET_0_120146);
    
    \U_EXEC_MASTER/USB_MASTER_EN/TERMCNT_FG40M2S\ : DFN1C0
      port map(D => 
        \U_EXEC_MASTER/USB_MASTER_EN/TERMCNT_FG40M1S_net_1\, CLK
         => CLK_40M_GL, CLR => P_MASTER_POR_B_c_32_0, Q => 
        \U_EXEC_MASTER/USB_MASTER_EN/TERMCNT_FG40M2S_net_1\);
    
    \U50_PATTERNS/U4D_REGCROSS/SAMP_TWO[5]\ : DFN1C0
      port map(D => \U50_PATTERNS/U4D_REGCROSS/SAMP_ONE[5]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_30, Q => 
        \U50_PATTERNS/U4D_REGCROSS/SAMP_TWO[5]_net_1\);
    
    HIEFFPLA_INST_0_53743 : AND2
      port map(A => HIEFFPLA_NET_0_117391, B => 
        HIEFFPLA_NET_0_117392, Y => HIEFFPLA_NET_0_117361);
    
    \U_ELK11_CH/U_SLAVE_1ELK/Q[12]\ : DFN1C0
      port map(D => \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/Q[12]_net_1\);
    
    HIEFFPLA_INST_0_111370 : NAND3C
      port map(A => HIEFFPLA_NET_0_116806, B => 
        HIEFFPLA_NET_0_116742, C => HIEFFPLA_NET_0_116687, Y => 
        HIEFFPLA_NET_0_115839);
    
    HIEFFPLA_INST_0_46406 : AO1
      port map(A => HIEFFPLA_NET_0_119244, B => 
        \U50_PATTERNS/ELINK_DOUTA_2[6]\, C => 
        HIEFFPLA_NET_0_118847, Y => HIEFFPLA_NET_0_118697);
    
    HIEFFPLA_INST_0_56291 : NAND3C
      port map(A => HIEFFPLA_NET_0_116875, B => 
        HIEFFPLA_NET_0_116883, C => HIEFFPLA_NET_0_116891, Y => 
        HIEFFPLA_NET_0_116899);
    
    \U50_PATTERNS/CHKSUM[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120138, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_3, Q => \U50_PATTERNS/CHKSUM[5]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_10[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116560, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_6, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_10[2]\);
    
    \U_ELK13_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118515, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_1, Q => 
        \U_ELK13_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]_net_1\);
    
    HIEFFPLA_INST_0_39668 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_6[2]\, B => 
        HIEFFPLA_NET_0_119522, S => HIEFFPLA_NET_0_119258, Y => 
        HIEFFPLA_NET_0_119965);
    
    \U_ELK14_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2\ : IOPADN_BI
      port map(DB => \U_ELK14_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, 
        E => \U_ELK14_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET3\, PAD
         => ELK14_DAT_N, N2POUT => 
        \U_ELK14_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2_N2P\);
    
    \U_EXEC_MASTER/USB_MASTER_EN/T_CNT60M[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117740, CLK => CLK60MHZ, CLR
         => P_MASTER_POR_B_c_28, Q => 
        \U_EXEC_MASTER/USB_MASTER_EN/T_CNT60M[3]_net_1\);
    
    \U50_PATTERNS/ELINKS_STOP_ADDR[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120124, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_14, Q => 
        \U50_PATTERNS/ELINKS_STOP_ADDR[3]\);
    
    HIEFFPLA_INST_0_58535 : NAND3C
      port map(A => HIEFFPLA_NET_0_116502, B => 
        HIEFFPLA_NET_0_116503, C => HIEFFPLA_NET_0_116504, Y => 
        HIEFFPLA_NET_0_116508);
    
    \U_ELK17_CH/U_ELK1_CMD_TX/START_RISE\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118329, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_8, Q => 
        \U_ELK17_CH/U_ELK1_CMD_TX/START_RISE_net_1\);
    
    HIEFFPLA_INST_0_58848 : MX2
      port map(A => HIEFFPLA_NET_0_116815, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_1[3]\, S => 
        HIEFFPLA_NET_0_117216, Y => HIEFFPLA_NET_0_116468);
    
    HIEFFPLA_INST_0_47726 : MX2
      port map(A => \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\, 
        B => \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[13]_net_1\, S => 
        \BIT_OS_SEL_2[2]\, Y => HIEFFPLA_NET_0_118441);
    
    HIEFFPLA_INST_0_38930 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_15[0]\, B => 
        HIEFFPLA_NET_0_119524, S => HIEFFPLA_NET_0_119297, Y => 
        HIEFFPLA_NET_0_120047);
    
    HIEFFPLA_INST_0_42535 : OA1A
      port map(A => HIEFFPLA_NET_0_119433, B => 
        HIEFFPLA_NET_0_119010, C => \U50_PATTERNS/REG_ADDR[6]\, Y
         => HIEFFPLA_NET_0_119517);
    
    \U_ELK8_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117886, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]_net_1\);
    
    HIEFFPLA_INST_0_58216 : MX2
      port map(A => HIEFFPLA_NET_0_116815, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_11[3]\, S => 
        HIEFFPLA_NET_0_117329, Y => HIEFFPLA_NET_0_116549);
    
    HIEFFPLA_INST_0_48567 : MX2
      port map(A => \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[0]_net_1\, 
        B => \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\, S => 
        \BIT_OS_SEL_0[2]\, Y => HIEFFPLA_NET_0_118294);
    
    HIEFFPLA_INST_0_55484 : MX2
      port map(A => HIEFFPLA_NET_0_116965, B => 
        HIEFFPLA_NET_0_117028, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[2]\, Y => 
        HIEFFPLA_NET_0_117031);
    
    HIEFFPLA_INST_0_61097 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_3[2]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_19[2]\, S
         => \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_1[4]_net_1\, 
        Y => HIEFFPLA_NET_0_116174);
    
    HIEFFPLA_INST_0_44134 : MX2
      port map(A => \U50_PATTERNS/TFC_STRT_ADDR[3]\, B => 
        \U50_PATTERNS/TFC_STRT_ADDR_T[3]\, S => 
        HIEFFPLA_NET_0_119472, Y => HIEFFPLA_NET_0_119169);
    
    \U50_PATTERNS/ELINK_ADDRA_12[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120070, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_2_0, Q => 
        \U50_PATTERNS/ELINK_ADDRA_12[1]\);
    
    HIEFFPLA_INST_0_39308 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_1[2]\, B => 
        HIEFFPLA_NET_0_119522, S => HIEFFPLA_NET_0_119243, Y => 
        HIEFFPLA_NET_0_120005);
    
    \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_115934, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_9, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[0]\);
    
    \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[6]\ : DFN1C0
      port map(D => 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\);
    
    \U50_PATTERNS/ELINKS_STRT_ADDR[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120111, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_17, Q => 
        \U50_PATTERNS/ELINKS_STRT_ADDR[0]\);
    
    HIEFFPLA_INST_0_53528 : AND3B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[4]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[2]_net_1\, C => 
        HIEFFPLA_NET_0_117318, Y => HIEFFPLA_NET_0_117393);
    
    HIEFFPLA_INST_0_37544 : MX2
      port map(A => TFC_RWB, B => \U200A_TFC/N_232_li\, S => 
        \U200A_TFC/GP_PG_SM[10]_net_1\, Y => 
        HIEFFPLA_NET_0_120263);
    
    \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[4]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117057, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_27, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[4]_net_1\);
    
    \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[3]\ : DFN1C0
      port map(D => 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[3]_net_1\);
    
    HIEFFPLA_INST_0_47636 : MX2
      port map(A => \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[2]_net_1\, 
        B => \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\, S => 
        \BIT_OS_SEL_2[2]\, Y => HIEFFPLA_NET_0_118454);
    
    HIEFFPLA_INST_0_62673 : NAND2A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_CLKPHASE[0]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_SEQCNT[1]\, Y => 
        HIEFFPLA_NET_0_115960);
    
    HIEFFPLA_INST_0_41224 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_3[6]\, B => 
        HIEFFPLA_NET_0_119566, S => HIEFFPLA_NET_0_119247, Y => 
        HIEFFPLA_NET_0_119761);
    
    HIEFFPLA_INST_0_111247 : NAND3C
      port map(A => HIEFFPLA_NET_0_116806, B => 
        HIEFFPLA_NET_0_116742, C => HIEFFPLA_NET_0_116687, Y => 
        HIEFFPLA_NET_0_115847);
    
    \U50_PATTERNS/REG_STATE[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119461, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_22_0, Q => 
        \U50_PATTERNS/REG_STATE[2]_net_1\);
    
    HIEFFPLA_INST_0_58770 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_19[3]\, B => 
        HIEFFPLA_NET_0_116476, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_2[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116478);
    
    HIEFFPLA_INST_0_51690 : MX2
      port map(A => \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[48]\, B
         => \U_MASTER_DES/PHASE_ADJ_160_L[2]\, S => 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM_0[4]_net_1\, Y => 
        HIEFFPLA_NET_0_117724);
    
    HIEFFPLA_INST_0_43128 : AND2A
      port map(A => \U50_PATTERNS/REG_STATE[3]_net_1\, B => 
        \U50_PATTERNS/REG_STATE[0]_net_1\, Y => 
        HIEFFPLA_NET_0_119365);
    
    HIEFFPLA_INST_0_46903 : MX2
      port map(A => \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\, 
        B => \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\, S => 
        \BIT_OS_SEL_4[2]\, Y => HIEFFPLA_NET_0_118587);
    
    \U50_PATTERNS/U103_PATT_ELINK_BLK/DPRT_512X9_SRAM_R0C0\ : 
        RAM4K9
      generic map(MEMORYFILE => "DPRT_512X9_SRAM_R0C0.mem")

      port map(ADDRA11 => AFLSDF_GND, ADDRA10 => AFLSDF_GND, 
        ADDRA9 => AFLSDF_GND, ADDRA8 => \GND\, ADDRA7 => 
        \U50_PATTERNS/ELINK_ADDRA_3[7]\, ADDRA6 => 
        \U50_PATTERNS/ELINK_ADDRA_3[6]\, ADDRA5 => 
        \U50_PATTERNS/ELINK_ADDRA_3[5]\, ADDRA4 => 
        \U50_PATTERNS/ELINK_ADDRA_3[4]\, ADDRA3 => 
        \U50_PATTERNS/ELINK_ADDRA_3[3]\, ADDRA2 => 
        \U50_PATTERNS/ELINK_ADDRA_3[2]\, ADDRA1 => 
        \U50_PATTERNS/ELINK_ADDRA_3[1]\, ADDRA0 => 
        \U50_PATTERNS/ELINK_ADDRA_3[0]\, ADDRB11 => AFLSDF_GND, 
        ADDRB10 => AFLSDF_GND, ADDRB9 => AFLSDF_GND, ADDRB8 => 
        \GND\, ADDRB7 => \ELKS_ADDRB[7]\, ADDRB6 => 
        \ELKS_ADDRB_0[6]\, ADDRB5 => \ELKS_ADDRB[5]\, ADDRB4 => 
        \ELKS_ADDRB_0[4]\, ADDRB3 => \ELKS_ADDRB[3]\, ADDRB2 => 
        \ELKS_ADDRB_0[2]\, ADDRB1 => \ELKS_ADDRB[1]\, ADDRB0 => 
        \ELKS_ADDRB[0]\, DINA8 => \GND\, DINA7 => 
        \U50_PATTERNS/ELINK_DINA_3[7]\, DINA6 => 
        \U50_PATTERNS/ELINK_DINA_3[6]\, DINA5 => 
        \U50_PATTERNS/ELINK_DINA_3[5]\, DINA4 => 
        \U50_PATTERNS/ELINK_DINA_3[4]\, DINA3 => 
        \U50_PATTERNS/ELINK_DINA_3[3]\, DINA2 => 
        \U50_PATTERNS/ELINK_DINA_3[2]\, DINA1 => 
        \U50_PATTERNS/ELINK_DINA_3[1]\, DINA0 => 
        \U50_PATTERNS/ELINK_DINA_3[0]\, DINB8 => \GND\, DINB7 => 
        \ELK_RX_SER_WORD_3[7]\, DINB6 => \ELK_RX_SER_WORD_3[6]\, 
        DINB5 => \ELK_RX_SER_WORD_3[5]\, DINB4 => 
        \ELK_RX_SER_WORD_3[4]\, DINB3 => \ELK_RX_SER_WORD_3[3]\, 
        DINB2 => \ELK_RX_SER_WORD_3[2]\, DINB1 => 
        \ELK_RX_SER_WORD_3[1]\, DINB0 => \ELK_RX_SER_WORD_3[0]\, 
        WIDTHA0 => \VCC\, WIDTHA1 => \VCC\, WIDTHB0 => \VCC\, 
        WIDTHB1 => \VCC\, PIPEA => \VCC\, PIPEB => \VCC\, WMODEA
         => \GND\, WMODEB => \GND\, BLKA => 
        \U50_PATTERNS/ELINK_BLKA[3]\, BLKB => ELKS_RAM_BLKB_EN, 
        WENA => \U50_PATTERNS/ELINK_RWA[3]\, WENB => ELKS_RWB, 
        CLKA => CLK60MHZ, CLKB => CLK_40M_GL, RESET => 
        P_USB_MASTER_EN_c_0, DOUTA8 => OPEN, DOUTA7 => 
        \U50_PATTERNS/ELINK_DOUTA_3[7]\, DOUTA6 => 
        \U50_PATTERNS/ELINK_DOUTA_3[6]\, DOUTA5 => 
        \U50_PATTERNS/ELINK_DOUTA_3[5]\, DOUTA4 => 
        \U50_PATTERNS/ELINK_DOUTA_3[4]\, DOUTA3 => 
        \U50_PATTERNS/ELINK_DOUTA_3[3]\, DOUTA2 => 
        \U50_PATTERNS/ELINK_DOUTA_3[2]\, DOUTA1 => 
        \U50_PATTERNS/ELINK_DOUTA_3[1]\, DOUTA0 => 
        \U50_PATTERNS/ELINK_DOUTA_3[0]\, DOUTB8 => OPEN, DOUTB7
         => \PATT_ELK_DAT_3[7]\, DOUTB6 => \PATT_ELK_DAT_3[6]\, 
        DOUTB5 => \PATT_ELK_DAT_3[5]\, DOUTB4 => 
        \PATT_ELK_DAT_3[4]\, DOUTB3 => \PATT_ELK_DAT_3[3]\, 
        DOUTB2 => \PATT_ELK_DAT_3[2]\, DOUTB1 => 
        \PATT_ELK_DAT_3[1]\, DOUTB0 => \PATT_ELK_DAT_3[0]\);
    
    \U_ELK5_CH/U_ELK1_SERDAT_SOURCE/SERDAT[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118010, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_17, Q => 
        \U_ELK5_CH/ELK_TX_DAT[3]\);
    
    \U_ELK18_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U0\ : IOPADP_BI
      port map(N2PIN => 
        \U_ELK18_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2_N2P\, D => 
        \U_ELK18_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, E => 
        \U_ELK18_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET2\, PAD => 
        ELK18_DAT_P, Y => 
        \U_ELK18_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\);
    
    \U50_PATTERNS/ELINK_DINA_10[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119863, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_9, Q => 
        \U50_PATTERNS/ELINK_DINA_10[0]\);
    
    HIEFFPLA_INST_0_53308 : AND2A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[8]_net_1\, B => 
        HIEFFPLA_NET_0_116978, Y => HIEFFPLA_NET_0_117434);
    
    \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[12]\ : DFN1C0
      port map(D => \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\);
    
    HIEFFPLA_INST_0_41954 : NAND2B
      port map(A => \U50_PATTERNS/ELINK_RWA[2]\, B => 
        HIEFFPLA_NET_0_119646, Y => HIEFFPLA_NET_0_119647);
    
    HIEFFPLA_INST_0_62340 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_3[3]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_4[3]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_4[0]\, Y => 
        HIEFFPLA_NET_0_116001);
    
    HIEFFPLA_INST_0_45708 : NAND2A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_4[7]\, Y => 
        HIEFFPLA_NET_0_118861);
    
    HIEFFPLA_INST_0_44730 : MX2
      port map(A => \OP_MODE_c_2[1]\, B => 
        \U50_PATTERNS/U4E_REGCROSS/SAMP_TWO[1]_net_1\, S => 
        HIEFFPLA_NET_0_119072, Y => HIEFFPLA_NET_0_119060);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_25[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116094, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_10, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_25[1]\);
    
    \U_ELK6_CH/U_ELK1_SERDAT_SOURCE/SERDAT[4]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117964, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_1, Q => 
        \U_ELK6_CH/ELK_TX_DAT[4]\);
    
    HIEFFPLA_INST_0_51400 : AND3A
      port map(A => HIEFFPLA_NET_0_117784, B => 
        \U_EXEC_MASTER/DEL_CNT[5]\, C => HIEFFPLA_NET_0_117780, Y
         => HIEFFPLA_NET_0_117787);
    
    HIEFFPLA_INST_0_48437 : MX2
      port map(A => \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\, 
        B => \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[11]_net_1\, S => 
        \BIT_OS_SEL_0[2]\, Y => HIEFFPLA_NET_0_118311);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_4[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116000, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_13, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_4[0]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/BEST_SEQCNT[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117442, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_8, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_SEQCNT[0]\);
    
    HIEFFPLA_INST_0_57099 : AND2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_2[5]\, B => 
        HIEFFPLA_NET_0_116736, Y => HIEFFPLA_NET_0_116744);
    
    HIEFFPLA_INST_0_53070 : MX2
      port map(A => HIEFFPLA_NET_0_117561, B => 
        HIEFFPLA_NET_0_117557, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[2]\, Y => 
        HIEFFPLA_NET_0_117469);
    
    \U_ELK14_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]\ : DFN1C0
      port map(D => \U_ELK14_CH/U_SLAVE_1ELK/Q[10]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_11[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116552, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_8, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_11[2]\);
    
    HIEFFPLA_INST_0_54309 : MX2
      port map(A => HIEFFPLA_NET_0_116516, B => 
        HIEFFPLA_NET_0_116299, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_2[3]_net_1\, Y
         => HIEFFPLA_NET_0_117282);
    
    HIEFFPLA_INST_0_43515 : MX2
      port map(A => \U50_PATTERNS/SM_BANK_SEL[8]\, B => 
        HIEFFPLA_NET_0_119210, S => HIEFFPLA_NET_0_118691, Y => 
        HIEFFPLA_NET_0_119302);
    
    HIEFFPLA_INST_0_59181 : MX2
      port map(A => HIEFFPLA_NET_0_116708, B => 
        HIEFFPLA_NET_0_116421, S => HIEFFPLA_NET_0_117264, Y => 
        HIEFFPLA_NET_0_116423);
    
    \U_EXEC_MASTER/MPOR_B_23\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117787, CLK => CLK_40M_GL, CLR
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_1\, Q => 
        P_MASTER_POR_B_c_23);
    
    \U_ELK3_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]\ : DFN1C0
      port map(D => \U_ELK3_CH/U_SLAVE_1ELK/Q[9]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]_net_1\);
    
    HIEFFPLA_INST_0_61595 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_24[1]\, B => 
        HIEFFPLA_NET_0_117167, S => HIEFFPLA_NET_0_117074, Y => 
        HIEFFPLA_NET_0_116104);
    
    HIEFFPLA_INST_0_59074 : AND2A
      port map(A => HIEFFPLA_NET_0_117214, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_3[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116438);
    
    \U200A_TFC/GP_PG_SM[6]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120314, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_28, Q => 
        \U200A_TFC/GP_PG_SM[6]_net_1\);
    
    HIEFFPLA_INST_0_62427 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_5[4]\, 
        B => HIEFFPLA_NET_0_117100, S => HIEFFPLA_NET_0_117172, Y
         => HIEFFPLA_NET_0_115991);
    
    HIEFFPLA_INST_0_56136 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/MAX_CNT[8]\, 
        B => HIEFFPLA_NET_0_116931, S => HIEFFPLA_NET_0_117084, Y
         => HIEFFPLA_NET_0_116946);
    
    HIEFFPLA_INST_0_37127 : AND3B
      port map(A => \U200A_TFC/LOC_STRT_ADDR[6]\, B => 
        HIEFFPLA_NET_0_120293, C => HIEFFPLA_NET_0_120328, Y => 
        HIEFFPLA_NET_0_120342);
    
    \U_ELK18_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118292, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_3, Q => 
        \U_ELK18_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]_net_1\);
    
    AFLSDF_INV_19 : INV
      port map(A => DCB_SALT_SEL_c, Y => \AFLSDF_INV_19\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_25[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116418, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_20, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_25[2]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_7[4]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116599, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_14, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_7[4]\);
    
    HIEFFPLA_INST_0_42428 : AND2
      port map(A => HIEFFPLA_NET_0_119473, B => 
        \U50_PATTERNS/RD_XFER_TYPE[4]_net_1\, Y => 
        HIEFFPLA_NET_0_119537);
    
    \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[12]\ : DFN1C0
      port map(D => \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\);
    
    HIEFFPLA_INST_0_56231 : AND3
      port map(A => HIEFFPLA_NET_0_116907, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/RECD_SER_WORD[2]_net_1\, 
        C => 
        \U_MASTER_DES/U13C_MASTER_DESER/RECD_SER_WORD[1]_net_1\, 
        Y => HIEFFPLA_NET_0_116924);
    
    HIEFFPLA_INST_0_55427 : AO1
      port map(A => HIEFFPLA_NET_0_117087, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[2]\, C => 
        HIEFFPLA_NET_0_117038, Y => HIEFFPLA_NET_0_117039);
    
    HIEFFPLA_INST_0_113075 : AO18
      port map(A => \U200A_TFC/LOC_STOP_ADDR[5]\, B => 
        \TFC_ADDRB[5]\, C => HIEFFPLA_NET_0_120294, Y => 
        HIEFFPLA_NET_0_115810);
    
    \U_ELK1_CH/ELK_IN_F\ : DFN1C0
      port map(D => \AFLSDF_INV_55\, CLK => CCC_160M_ADJ, CLR => 
        DEV_RST_B_c, Q => \U_ELK1_CH/ELK_IN_F_net_1\);
    
    HIEFFPLA_INST_0_47826 : MX2
      port map(A => \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\, 
        B => \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[14]_net_1\, S => 
        \BIT_OS_SEL_5[2]\, Y => HIEFFPLA_NET_0_118428);
    
    HIEFFPLA_INST_0_53190 : MX2
      port map(A => HIEFFPLA_NET_0_117530, B => 
        HIEFFPLA_NET_0_117522, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[3]\, Y => 
        HIEFFPLA_NET_0_117454);
    
    \U50_PATTERNS/ELINK_DINA_13[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119836, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_14, Q => 
        \U50_PATTERNS/ELINK_DINA_13[3]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[8]\ : DFN1P0
      port map(D => HIEFFPLA_NET_0_117188, CLK => CLK_40M_GL, PRE
         => P_MASTER_POR_B_c_27, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[8]_net_1\);
    
    HIEFFPLA_INST_0_55038 : AOI1D
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[6]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[8]_net_1\, C => 
        HIEFFPLA_NET_0_116774, Y => HIEFFPLA_NET_0_117136);
    
    HIEFFPLA_INST_0_43640 : NAND2B
      port map(A => \U50_PATTERNS/SM_BANK_SEL[21]\, B => 
        \U50_PATTERNS/SM_BANK_SEL[3]\, Y => HIEFFPLA_NET_0_119257);
    
    HIEFFPLA_INST_0_44488 : MX2
      port map(A => \ELKS_STRT_ADDR[5]\, B => 
        \U50_PATTERNS/U4C_REGCROSS/SAMP_TWO[5]_net_1\, S => 
        HIEFFPLA_NET_0_119114, Y => HIEFFPLA_NET_0_119107);
    
    AFLSDF_INV_17 : INV
      port map(A => DCB_SALT_SEL_c, Y => \AFLSDF_INV_17\);
    
    HIEFFPLA_INST_0_54743 : NAND3A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[4]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[2]_net_1\, C => 
        HIEFFPLA_NET_0_117242, Y => HIEFFPLA_NET_0_117210);
    
    \U50_PATTERNS/TFC_STOP_ADDR_T[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119176, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_15, Q => 
        \U50_PATTERNS/TFC_STOP_ADDR_T[4]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_2[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116755, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_5, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_2[0]\);
    
    \U_ELK10_CH/ELK_IN_F\ : DFN1C0
      port map(D => \U_ELK10_CH/ELK_IN_DDR_F\, CLK => 
        CCC_160M_ADJ, CLR => DEV_RST_B_c, Q => 
        \U_ELK10_CH/ELK_IN_F_net_1\);
    
    \U50_PATTERNS/ELINK_ADDRA_16[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120034, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_9, Q => 
        \U50_PATTERNS/ELINK_ADDRA_16[5]\);
    
    \P_TFC_SYNC_DET_pad/U0/U0\ : IOPAD_TRI_U
      port map(D => \P_TFC_SYNC_DET_pad/U0/NET1\, E => 
        \P_TFC_SYNC_DET_pad/U0/NET2\, PAD => P_TFC_SYNC_DET);
    
    HIEFFPLA_INST_0_47615 : MX2
      port map(A => 
        \U_ELK14_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]_net_1\, B => 
        \U_ELK14_CH/ELK_TX_DAT[7]\, S => 
        \U_ELK14_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118465);
    
    HIEFFPLA_INST_0_42449 : MX2
      port map(A => \U50_PATTERNS/REG_ADDR[1]\, B => 
        HIEFFPLA_NET_0_119508, S => HIEFFPLA_NET_0_119007, Y => 
        HIEFFPLA_NET_0_119532);
    
    \U_ELK7_CH/U_SLAVE_1ELK/RECD_SER_WORD[4]\ : DFN1C0
      port map(D => \U_ELK7_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[4]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_7[4]\);
    
    \U50_PATTERNS/U4A_REGCROSS/LOCAL_REG_VAL[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119151, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_17, Q => \TFC_STRT_ADDR[3]\);
    
    \U_ELK10_CH/U_SLAVE_1ELK/Q[2]\ : DFN1C0
      port map(D => \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/Q[2]_net_1\);
    
    HIEFFPLA_INST_0_54638 : MX2
      port map(A => HIEFFPLA_NET_0_117194, B => 
        HIEFFPLA_NET_0_117352, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[1]_net_1\, Y => 
        HIEFFPLA_NET_0_117229);
    
    \U_ELK2_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118154, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_12, Q => 
        \U_ELK2_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]_net_1\);
    
    HIEFFPLA_INST_0_55339 : AND2A
      port map(A => HIEFFPLA_NET_0_117269, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_3[6]_net_1\, Y => 
        HIEFFPLA_NET_0_117056);
    
    HIEFFPLA_INST_0_51525 : AOI1B
      port map(A => HIEFFPLA_NET_0_117747, B => 
        HIEFFPLA_NET_0_117745, C => 
        \U_EXEC_MASTER/USB_MASTER_EN/CNT_EN_60M2S_net_1\, Y => 
        HIEFFPLA_NET_0_117753);
    
    \U_ELK10_CH/U_SLAVE_1ELK/Q[0]\ : DFN1C0
      port map(D => \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/Q[0]_net_1\);
    
    HIEFFPLA_INST_0_55208 : AND2A
      port map(A => HIEFFPLA_NET_0_117206, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[6]_net_1\, Y => 
        HIEFFPLA_NET_0_117090);
    
    HIEFFPLA_INST_0_49097 : MX2
      port map(A => HIEFFPLA_NET_0_118198, B => 
        \U_ELK1_CH/ELK_TX_DAT[3]\, S => 
        \U_ELK1_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118197);
    
    HIEFFPLA_INST_0_45640 : NAND3C
      port map(A => HIEFFPLA_NET_0_118718, B => 
        HIEFFPLA_NET_0_118892, C => HIEFFPLA_NET_0_118708, Y => 
        HIEFFPLA_NET_0_118875);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_7[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116601, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_14, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_7[2]\);
    
    \U_ELK3_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]\ : DFN1C0
      port map(D => \U_ELK3_CH/U_SLAVE_1ELK/Q[0]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]_net_1\);
    
    \U50_PATTERNS/ELINKS_STOP_ADDR[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120126, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_14, Q => 
        \U50_PATTERNS/ELINKS_STOP_ADDR[1]\);
    
    \U_ELK3_CH/U_SLAVE_1ELK/Q[6]\ : DFN1C0
      port map(D => \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/Q[6]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_23[4]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116116, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_6, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_23[4]\);
    
    HIEFFPLA_INST_0_41737 : MX2
      port map(A => HIEFFPLA_NET_0_119681, B => 
        \U50_PATTERNS/ELINK_RWA[18]\, S => 
        \U50_PATTERNS/SM_BANK_SEL_0[20]\, Y => 
        HIEFFPLA_NET_0_119702);
    
    HIEFFPLA_INST_0_37632 : AND3B
      port map(A => \U200B_ELINKS/LOC_STRT_ADDR[0]\, B => 
        HIEFFPLA_NET_0_120190, C => HIEFFPLA_NET_0_120234, Y => 
        HIEFFPLA_NET_0_120243);
    
    \U50_PATTERNS/RD_XFER_TYPE[4]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119545, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c, Q => 
        \U50_PATTERNS/RD_XFER_TYPE[4]_net_1\);
    
    HIEFFPLA_INST_0_48246 : MX2
      port map(A => HIEFFPLA_NET_0_118356, B => 
        HIEFFPLA_NET_0_118352, S => \BIT_OS_SEL_3[0]\, Y => 
        \U_ELK16_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[1]\);
    
    HIEFFPLA_INST_0_37540 : AND2B
      port map(A => \U200A_TFC/GP_PG_SM[10]_net_1\, B => 
        \U200A_TFC/GP_PG_SM[1]_net_1\, Y => HIEFFPLA_NET_0_120264);
    
    HIEFFPLA_INST_0_37249 : AND3A
      port map(A => HIEFFPLA_NET_0_120305, B => 
        \U200A_TFC/GP_PG_SM[8]_net_1\, C => HIEFFPLA_NET_0_120330, 
        Y => HIEFFPLA_NET_0_120315);
    
    \U_ELK11_CH/U_ELK1_SERDAT_SOURCE/SERDAT[5]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118593, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_0, Q => 
        \U_ELK11_CH/ELK_TX_DAT[5]\);
    
    HIEFFPLA_INST_0_54918 : AO1C
      port map(A => HIEFFPLA_NET_0_117205, B => 
        HIEFFPLA_NET_0_117116, C => HIEFFPLA_NET_0_117180, Y => 
        HIEFFPLA_NET_0_117170);
    
    \U50_PATTERNS/SM_BANK_SEL[21]/U1\ : DFN1P0
      port map(D => HIEFFPLA_NET_0_119309, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_2, Q => 
        \U50_PATTERNS/SM_BANK_SEL[21]\);
    
    HIEFFPLA_INST_0_55973 : MX2
      port map(A => HIEFFPLA_NET_0_116005, B => 
        HIEFFPLA_NET_0_116256, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[3]\, Y => 
        HIEFFPLA_NET_0_116966);
    
    \U_ELK5_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U0\ : IOPADP_BI
      port map(N2PIN => 
        \U_ELK5_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2_N2P\, D => 
        \U_ELK5_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, E => 
        \U_ELK5_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET2\, PAD => 
        ELK5_DAT_P, Y => 
        \U_ELK5_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\);
    
    \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[7]\ : DFN1C0
      port map(D => \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\);
    
    \U_ELK18_CH/U_SLAVE_1ELK/RECD_SER_WORD[7]\ : DFN1C0
      port map(D => \U_ELK18_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[7]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_18[7]\);
    
    HIEFFPLA_INST_0_56181 : XA1C
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/MAX_CNT[4]\, 
        B => HIEFFPLA_NET_0_116941, C => HIEFFPLA_NET_0_117112, Y
         => HIEFFPLA_NET_0_116935);
    
    \U_ELK9_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]\ : DFN1C0
      port map(D => \U_ELK9_CH/U_SLAVE_1ELK/Q[1]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]_net_1\);
    
    HIEFFPLA_INST_0_53821 : MX2
      port map(A => HIEFFPLA_NET_0_116192, B => 
        HIEFFPLA_NET_0_116088, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[3]_net_1\, Y
         => HIEFFPLA_NET_0_117347);
    
    \U_ELK9_CH/U_SLAVE_1ELK/Q[2]\ : DFN1C0
      port map(D => \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/Q[2]_net_1\);
    
    \U_ELK14_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL\ : DFN1C0
      port map(D => 
        \U_ELK14_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL_net_1\);
    
    HIEFFPLA_INST_0_54999 : NAND2B
      port map(A => HIEFFPLA_NET_0_117182, B => 
        HIEFFPLA_NET_0_117143, Y => HIEFFPLA_NET_0_117144);
    
    HIEFFPLA_INST_0_46296 : NAND3C
      port map(A => HIEFFPLA_NET_0_118792, B => 
        HIEFFPLA_NET_0_118895, C => HIEFFPLA_NET_0_118722, Y => 
        HIEFFPLA_NET_0_118723);
    
    \U_ELK2_CH/U_ELK1_SERDAT_SOURCE/SERDAT[6]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118142, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_13, Q => 
        \U_ELK2_CH/ELK_TX_DAT[6]\);
    
    HIEFFPLA_INST_0_111249 : NAND3C
      port map(A => HIEFFPLA_NET_0_116806, B => 
        HIEFFPLA_NET_0_116742, C => HIEFFPLA_NET_0_116687, Y => 
        HIEFFPLA_NET_0_115846);
    
    \ALL_PLL_LOCK_pad/U0/U0\ : IOPAD_TRI_U
      port map(D => \ALL_PLL_LOCK_pad/U0/NET1\, E => 
        \ALL_PLL_LOCK_pad/U0/NET2\, PAD => ALL_PLL_LOCK);
    
    HIEFFPLA_INST_0_47820 : MX2
      port map(A => \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[0]_net_1\, 
        B => \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\, S => 
        \BIT_OS_SEL_2[2]\, Y => HIEFFPLA_NET_0_118429);
    
    HIEFFPLA_INST_0_39614 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_5[4]\, B => 
        HIEFFPLA_NET_0_119519, S => HIEFFPLA_NET_0_119251, Y => 
        HIEFFPLA_NET_0_119971);
    
    \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[11]\ : DFN1C0
      port map(D => 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[11]_net_1\);
    
    \U50_PATTERNS/ELINK_BLKA[14]/U1\ : DFN1P0
      port map(D => HIEFFPLA_NET_0_119930, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_20, Q => 
        \U50_PATTERNS/ELINK_BLKA[14]\);
    
    HIEFFPLA_INST_0_55326 : AOI1
      port map(A => HIEFFPLA_NET_0_115919, B => 
        HIEFFPLA_NET_0_117054, C => HIEFFPLA_NET_0_117051, Y => 
        HIEFFPLA_NET_0_117059);
    
    HIEFFPLA_INST_0_37696 : AO1A
      port map(A => \OP_MODE_c[6]\, B => 
        \U200B_ELINKS/GP_PG_SM[0]_net_1\, C => 
        HIEFFPLA_NET_0_120230, Y => HIEFFPLA_NET_0_120227);
    
    \U50_PATTERNS/ELINK_ADDRA_6[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119965, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_4, Q => 
        \U50_PATTERNS/ELINK_ADDRA_6[2]\);
    
    HIEFFPLA_INST_0_46856 : MX2
      port map(A => 
        \U_ELK11_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]_net_1\, B => 
        \U_ELK11_CH/ELK_TX_DAT[3]\, S => 
        \U_ELK11_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118602);
    
    \U_ELK4_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]\ : DFN1C0
      port map(D => \U_ELK4_CH/U_SLAVE_1ELK/Q[11]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]_net_1\);
    
    \U_ELK3_CH/ELK_IN_R\ : DFN1C0
      port map(D => \AFLSDF_INV_56\, CLK => CCC_160M_ADJ, CLR => 
        DEV_RST_B_c, Q => \U_ELK3_CH/ELK_IN_R_net_1\);
    
    HIEFFPLA_INST_0_57608 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_5[8]\, B => 
        HIEFFPLA_NET_0_116636, S => HIEFFPLA_NET_0_117121, Y => 
        HIEFFPLA_NET_0_116653);
    
    HIEFFPLA_INST_0_51797 : MX2
      port map(A => \U_MASTER_DES/U13A_ADJ_160M/BITCNT[7]\, B => 
        HIEFFPLA_NET_0_117675, S => HIEFFPLA_NET_0_117630, Y => 
        HIEFFPLA_NET_0_117691);
    
    HIEFFPLA_INST_0_42814 : AND3A
      port map(A => HIEFFPLA_NET_0_119379, B => 
        HIEFFPLA_NET_0_119432, C => HIEFFPLA_NET_0_119393, Y => 
        HIEFFPLA_NET_0_119458);
    
    \U50_PATTERNS/ELINK_ADDRA_9[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119938, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_10, Q => 
        \U50_PATTERNS/ELINK_ADDRA_9[5]\);
    
    \U200A_TFC/GP_PG_SM[9]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120310, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_28, Q => 
        \U200A_TFC/GP_PG_SM[9]_net_1\);
    
    HIEFFPLA_INST_0_55110 : AO1
      port map(A => HIEFFPLA_NET_0_117128, B => 
        HIEFFPLA_NET_0_117586, C => HIEFFPLA_NET_0_117179, Y => 
        HIEFFPLA_NET_0_117120);
    
    HIEFFPLA_INST_0_53878 : MX2
      port map(A => HIEFFPLA_NET_0_117381, B => 
        HIEFFPLA_NET_0_117200, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[0]_net_1\, Y
         => HIEFFPLA_NET_0_117338);
    
    HIEFFPLA_INST_0_38687 : MX2
      port map(A => HIEFFPLA_NET_0_119518, B => 
        \U50_PATTERNS/ELINK_ADDRA_11[5]\, S => 
        HIEFFPLA_NET_0_119280, Y => HIEFFPLA_NET_0_120074);
    
    \U50_PATTERNS/ELINK_ADDRA_3[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119984, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_1_0, Q => 
        \U50_PATTERNS/ELINK_ADDRA_3[7]\);
    
    \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[13]\ : DFN1C0
      port map(D => \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[13]_net_1\);
    
    HIEFFPLA_INST_0_45463 : AO1
      port map(A => HIEFFPLA_NET_0_119263, B => 
        \U50_PATTERNS/ELINK_DOUTA_8[4]\, C => 
        HIEFFPLA_NET_0_118808, Y => HIEFFPLA_NET_0_118909);
    
    \U_ELK17_CH/U_SLAVE_1ELK/Q[8]\ : DFN1C0
      port map(D => \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/Q[8]_net_1\);
    
    \U0A_40M_REFCLK/_BIBUF_LVDS[0]_/U0/U3\ : IOBI_IB_OB_EB
      port map(D => CLK40M_10NS_REF, E => \AFLSDF_INV_3\, YIN => 
        \U0A_40M_REFCLK/\\\\BIBUF_LVDS[0]\\\\/U0/NET4\, DOUT => 
        OPEN, EOUT => 
        \U0A_40M_REFCLK/\\\\BIBUF_LVDS[0]\\\\/U0/NET3\, Y => OPEN);
    
    HIEFFPLA_INST_0_62355 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_4[1]\, 
        B => HIEFFPLA_NET_0_117114, S => HIEFFPLA_NET_0_117148, Y
         => HIEFFPLA_NET_0_115999);
    
    HIEFFPLA_INST_0_45581 : AO1A
      port map(A => HIEFFPLA_NET_0_119428, B => 
        \U50_PATTERNS/ELINKS_STRT_ADDR[3]\, C => 
        HIEFFPLA_NET_0_118791, Y => HIEFFPLA_NET_0_118886);
    
    HIEFFPLA_INST_0_53014 : MX2
      port map(A => HIEFFPLA_NET_0_117456, B => 
        HIEFFPLA_NET_0_117568, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[2]\, Y => 
        HIEFFPLA_NET_0_117476);
    
    HIEFFPLA_INST_0_55358 : AOI1D
      port map(A => HIEFFPLA_NET_0_116941, B => 
        HIEFFPLA_NET_0_116943, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[7]_net_1\, Y => 
        HIEFFPLA_NET_0_117052);
    
    HIEFFPLA_INST_0_46849 : MX2
      port map(A => 
        \U_ELK11_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]_net_1\, B => 
        \U_ELK11_CH/ELK_TX_DAT[6]\, S => 
        \U_ELK11_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118604);
    
    \U50_PATTERNS/ELINK_DINA_15[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119821, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_16, Q => 
        \U50_PATTERNS/ELINK_DINA_15[2]\);
    
    HIEFFPLA_INST_0_55393 : MX2
      port map(A => HIEFFPLA_NET_0_116956, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[1]\, S => 
        HIEFFPLA_NET_0_117087, Y => HIEFFPLA_NET_0_117044);
    
    HIEFFPLA_INST_0_48385 : MX2
      port map(A => \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[1]_net_1\, 
        B => \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\, S => 
        \BIT_OS_SEL_0[2]\, Y => HIEFFPLA_NET_0_118319);
    
    HIEFFPLA_INST_0_55194 : AND2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[6]_net_1\, B => 
        HIEFFPLA_NET_0_117335, Y => HIEFFPLA_NET_0_117097);
    
    HIEFFPLA_INST_0_55104 : AO1
      port map(A => HIEFFPLA_NET_0_117128, B => 
        HIEFFPLA_NET_0_117583, C => HIEFFPLA_NET_0_117179, Y => 
        HIEFFPLA_NET_0_117121);
    
    HIEFFPLA_INST_0_50543 : MX2
      port map(A => HIEFFPLA_NET_0_117934, B => 
        HIEFFPLA_NET_0_117955, S => \BIT_OS_SEL_5[1]\, Y => 
        HIEFFPLA_NET_0_117936);
    
    HIEFFPLA_INST_0_42842 : NAND2A
      port map(A => \U50_PATTERNS/REG_STATE[4]_net_1\, B => 
        \U50_PATTERNS/REG_STATE[0]_net_1\, Y => 
        HIEFFPLA_NET_0_119450);
    
    \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[14]\ : DFN1C0
      port map(D => \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[14]_net_1\);
    
    HIEFFPLA_INST_0_44640 : XO1
      port map(A => \ELKS_STOP_ADDR[4]\, B => 
        \U50_PATTERNS/U4D_REGCROSS/SAMP_TWO[4]_net_1\, C => 
        HIEFFPLA_NET_0_119075, Y => HIEFFPLA_NET_0_119078);
    
    HIEFFPLA_INST_0_42378 : AND2B
      port map(A => \U50_PATTERNS/RD_XFER_TYPE[2]_net_1\, B => 
        \U50_PATTERNS/RD_XFER_TYPE[5]_net_1\, Y => 
        HIEFFPLA_NET_0_119550);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_15[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116519, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_15, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_15[1]\);
    
    HIEFFPLA_INST_0_59534 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_12[0]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_28[0]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[4]_net_1\, Y
         => HIEFFPLA_NET_0_116382);
    
    HIEFFPLA_INST_0_50487 : MX2
      port map(A => HIEFFPLA_NET_0_117945, B => 
        HIEFFPLA_NET_0_117959, S => \BIT_OS_SEL[0]\, Y => 
        \U_ELK6_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[1]\);
    
    \U_ELK17_CH/U_ELK1_SERDAT_SOURCE/SERDAT[6]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118322, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_11, Q => 
        \U_ELK17_CH/ELK_TX_DAT[6]\);
    
    \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[13]\ : DFN1C0
      port map(D => \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[13]_net_1\);
    
    HIEFFPLA_INST_0_45011 : AO1
      port map(A => HIEFFPLA_NET_0_119372, B => 
        HIEFFPLA_NET_0_118999, C => HIEFFPLA_NET_0_119454, Y => 
        HIEFFPLA_NET_0_119000);
    
    \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[8]\ : DFN1C0
      port map(D => 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\);
    
    \U_ELK12_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]\ : DFN1C0
      port map(D => \U_ELK12_CH/U_SLAVE_1ELK/Q[6]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]_net_1\);
    
    HIEFFPLA_INST_0_40081 : AOI1C
      port map(A => \U50_PATTERNS/ELINK_BLKA[10]\, B => 
        HIEFFPLA_NET_0_119662, C => HIEFFPLA_NET_0_119912, Y => 
        HIEFFPLA_NET_0_119913);
    
    \U_ELK4_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0\ : DFN1C0
      port map(D => CLK_40M_GL, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_9, Q => 
        \U_ELK4_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0_net_1\);
    
    \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[11]\ : DFN1C0
      port map(D => 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]_net_1\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[11]_net_1\);
    
    \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[7]\ : DFN1C0
      port map(D => \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\);
    
    \U50_PATTERNS/U107_PATT_ELINK_BLK/DPRT_512X9_SRAM_R0C0\ : 
        RAM4K9
      generic map(MEMORYFILE => "DPRT_512X9_SRAM_R0C0.mem")

      port map(ADDRA11 => AFLSDF_GND, ADDRA10 => AFLSDF_GND, 
        ADDRA9 => AFLSDF_GND, ADDRA8 => \GND\, ADDRA7 => 
        \U50_PATTERNS/ELINK_ADDRA_7[7]\, ADDRA6 => 
        \U50_PATTERNS/ELINK_ADDRA_7[6]\, ADDRA5 => 
        \U50_PATTERNS/ELINK_ADDRA_7[5]\, ADDRA4 => 
        \U50_PATTERNS/ELINK_ADDRA_7[4]\, ADDRA3 => 
        \U50_PATTERNS/ELINK_ADDRA_7[3]\, ADDRA2 => 
        \U50_PATTERNS/ELINK_ADDRA_7[2]\, ADDRA1 => 
        \U50_PATTERNS/ELINK_ADDRA_7[1]\, ADDRA0 => 
        \U50_PATTERNS/ELINK_ADDRA_7[0]\, ADDRB11 => AFLSDF_GND, 
        ADDRB10 => AFLSDF_GND, ADDRB9 => AFLSDF_GND, ADDRB8 => 
        \GND\, ADDRB7 => \ELKS_ADDRB[7]\, ADDRB6 => 
        \ELKS_ADDRB_0[6]\, ADDRB5 => \ELKS_ADDRB[5]\, ADDRB4 => 
        \ELKS_ADDRB_0[4]\, ADDRB3 => \ELKS_ADDRB[3]\, ADDRB2 => 
        \ELKS_ADDRB_0[2]\, ADDRB1 => \ELKS_ADDRB[1]\, ADDRB0 => 
        \ELKS_ADDRB[0]\, DINA8 => \GND\, DINA7 => 
        \U50_PATTERNS/ELINK_DINA_7[7]\, DINA6 => 
        \U50_PATTERNS/ELINK_DINA_7[6]\, DINA5 => 
        \U50_PATTERNS/ELINK_DINA_7[5]\, DINA4 => 
        \U50_PATTERNS/ELINK_DINA_7[4]\, DINA3 => 
        \U50_PATTERNS/ELINK_DINA_7[3]\, DINA2 => 
        \U50_PATTERNS/ELINK_DINA_7[2]\, DINA1 => 
        \U50_PATTERNS/ELINK_DINA_7[1]\, DINA0 => 
        \U50_PATTERNS/ELINK_DINA_7[0]\, DINB8 => \GND\, DINB7 => 
        \ELK_RX_SER_WORD_7[7]\, DINB6 => \ELK_RX_SER_WORD_7[6]\, 
        DINB5 => \ELK_RX_SER_WORD_7[5]\, DINB4 => 
        \ELK_RX_SER_WORD_7[4]\, DINB3 => \ELK_RX_SER_WORD_7[3]\, 
        DINB2 => \ELK_RX_SER_WORD_7[2]\, DINB1 => 
        \ELK_RX_SER_WORD_7[1]\, DINB0 => \ELK_RX_SER_WORD_7[0]\, 
        WIDTHA0 => \VCC\, WIDTHA1 => \VCC\, WIDTHB0 => \VCC\, 
        WIDTHB1 => \VCC\, PIPEA => \VCC\, PIPEB => \VCC\, WMODEA
         => \GND\, WMODEB => \GND\, BLKA => 
        \U50_PATTERNS/ELINK_BLKA[7]\, BLKB => ELKS_RAM_BLKB_EN, 
        WENA => \U50_PATTERNS/ELINK_RWA[7]\, WENB => ELKS_RWB, 
        CLKA => CLK60MHZ, CLKB => CLK_40M_GL, RESET => 
        P_USB_MASTER_EN_c_0, DOUTA8 => OPEN, DOUTA7 => 
        \U50_PATTERNS/ELINK_DOUTA_7[7]\, DOUTA6 => 
        \U50_PATTERNS/ELINK_DOUTA_7[6]\, DOUTA5 => 
        \U50_PATTERNS/ELINK_DOUTA_7[5]\, DOUTA4 => 
        \U50_PATTERNS/ELINK_DOUTA_7[4]\, DOUTA3 => 
        \U50_PATTERNS/ELINK_DOUTA_7[3]\, DOUTA2 => 
        \U50_PATTERNS/ELINK_DOUTA_7[2]\, DOUTA1 => 
        \U50_PATTERNS/ELINK_DOUTA_7[1]\, DOUTA0 => 
        \U50_PATTERNS/ELINK_DOUTA_7[0]\, DOUTB8 => OPEN, DOUTB7
         => \PATT_ELK_DAT_7[7]\, DOUTB6 => \PATT_ELK_DAT_7[6]\, 
        DOUTB5 => \PATT_ELK_DAT_7[5]\, DOUTB4 => 
        \PATT_ELK_DAT_7[4]\, DOUTB3 => \PATT_ELK_DAT_7[3]\, 
        DOUTB2 => \PATT_ELK_DAT_7[2]\, DOUTB1 => 
        \PATT_ELK_DAT_7[1]\, DOUTB0 => \PATT_ELK_DAT_7[0]\);
    
    HIEFFPLA_INST_0_60429 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_9[3]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_10[3]\, S
         => \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_1[0]\, Y
         => HIEFFPLA_NET_0_116267);
    
    HIEFFPLA_INST_0_45538 : AO1A
      port map(A => HIEFFPLA_NET_0_119475, B => 
        \U50_PATTERNS/ELINKS_STOP_ADDR[3]\, C => 
        HIEFFPLA_NET_0_118809, Y => HIEFFPLA_NET_0_118894);
    
    HIEFFPLA_INST_0_44414 : NAND3C
      port map(A => HIEFFPLA_NET_0_119121, B => 
        HIEFFPLA_NET_0_119122, C => HIEFFPLA_NET_0_119123, Y => 
        HIEFFPLA_NET_0_119124);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_13[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116248, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_1, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_13[2]\);
    
    HIEFFPLA_INST_0_43044 : AND3B
      port map(A => \U50_PATTERNS/USB_TXE_B\, B => 
        \U50_PATTERNS/REG_STATE[3]_net_1\, C => 
        \U50_PATTERNS/REG_STATE[4]_net_1\, Y => 
        HIEFFPLA_NET_0_119393);
    
    HIEFFPLA_INST_0_60274 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_8[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_24[1]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_1[4]_net_1\, Y
         => HIEFFPLA_NET_0_116288);
    
    HIEFFPLA_INST_0_51242 : MX2
      port map(A => HIEFFPLA_NET_0_117822, B => 
        HIEFFPLA_NET_0_117818, S => \BIT_OS_SEL_4[0]\, Y => 
        \U_ELK9_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[2]\);
    
    HIEFFPLA_INST_0_54732 : NAND3B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[3]_net_1\, B => 
        HIEFFPLA_NET_0_117237, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[0]_net_1\, Y => 
        HIEFFPLA_NET_0_117214);
    
    HIEFFPLA_INST_0_47780 : MX2
      port map(A => HIEFFPLA_NET_0_118450, B => 
        HIEFFPLA_NET_0_118446, S => \BIT_OS_SEL_4[0]\, Y => 
        \U_ELK14_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[5]\);
    
    \U_ELK19_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL\ : DFN1C0
      port map(D => 
        \U_ELK19_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL_net_1\);
    
    HIEFFPLA_INST_0_43030 : AND3
      port map(A => HIEFFPLA_NET_0_119430, B => 
        HIEFFPLA_NET_0_119016, C => 
        \U50_PATTERNS/REG_STATE[1]_net_1\, Y => 
        HIEFFPLA_NET_0_119397);
    
    \U_ELK12_CH/U_ELK1_CMD_TX/SER_OUT_FI\ : DFN1C0
      port map(D => 
        \U_ELK12_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_10, Q
         => \U_ELK12_CH/U_ELK1_CMD_TX/SER_OUT_FI_net_1\);
    
    HIEFFPLA_INST_0_47194 : MX2
      port map(A => HIEFFPLA_NET_0_118539, B => 
        HIEFFPLA_NET_0_118535, S => \BIT_OS_SEL_4[1]\, Y => 
        HIEFFPLA_NET_0_118536);
    
    \U_ELK7_CH/U_ELK1_SERDAT_SOURCE/SERDAT[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117923, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_3, Q => 
        \U_ELK7_CH/ELK_TX_DAT[0]\);
    
    HIEFFPLA_INST_0_45176 : NAND3C
      port map(A => HIEFFPLA_NET_0_118799, B => 
        HIEFFPLA_NET_0_118877, C => HIEFFPLA_NET_0_118962, Y => 
        HIEFFPLA_NET_0_118971);
    
    HIEFFPLA_INST_0_53837 : MX2
      port map(A => HIEFFPLA_NET_0_117258, B => 
        HIEFFPLA_NET_0_117326, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[2]_net_1\, Y
         => HIEFFPLA_NET_0_117345);
    
    HIEFFPLA_INST_0_52344 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_BIT_OS_VAL[2]\, B
         => HIEFFPLA_NET_0_117574, S => HIEFFPLA_NET_0_117111, Y
         => HIEFFPLA_NET_0_117578);
    
    HIEFFPLA_INST_0_42392 : AO1A
      port map(A => HIEFFPLA_NET_0_119019, B => 
        \U50_PATTERNS/RD_USB_ADBUS[2]\, C => 
        HIEFFPLA_NET_0_119539, Y => HIEFFPLA_NET_0_119547);
    
    \U_EXEC_MASTER/DEV_RST_1B\ : DFI1C0
      port map(D => \U_EXEC_MASTER/DEV_RST_0B_net_1\, CLK => 
        CCC_160M_FXD, CLR => DEV_RST_B_c, QN => 
        \U_EXEC_MASTER/DEV_RST_1B_i\);
    
    \U_EXEC_MASTER/MPOR_B_0_0\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117787, CLK => CLK_40M_GL, CLR
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_2\, Q => 
        P_MASTER_POR_B_c_0_0);
    
    \U200A_TFC/RX_SER_WORD_2DEL[3]\ : DFN1C0
      port map(D => \U200A_TFC/RX_SER_WORD_1DEL[3]_net_1\, CLK
         => CLK_40M_GL, CLR => P_MASTER_POR_B_c, Q => 
        \U200A_TFC/RX_SER_WORD_2DEL[3]_net_1\);
    
    HIEFFPLA_INST_0_60597 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_13[4]\, B => 
        HIEFFPLA_NET_0_117166, S => HIEFFPLA_NET_0_117137, Y => 
        HIEFFPLA_NET_0_116246);
    
    \U_ELK18_CH/U_ELK1_CMD_TX/SER_OUT_RDEL\ : DFN1C0
      port map(D => \U_ELK18_CH/U_ELK1_CMD_TX/SER_OUT_RI_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_1, Q
         => \U_ELK18_CH/ELK_OUT_R\);
    
    HIEFFPLA_INST_0_49951 : MX2
      port map(A => HIEFFPLA_NET_0_118048, B => 
        HIEFFPLA_NET_0_118046, S => \BIT_OS_SEL_6[1]\, Y => 
        HIEFFPLA_NET_0_118038);
    
    HIEFFPLA_INST_0_46236 : NAND3C
      port map(A => HIEFFPLA_NET_0_118906, B => 
        HIEFFPLA_NET_0_118914, C => HIEFFPLA_NET_0_118917, Y => 
        HIEFFPLA_NET_0_118734);
    
    HIEFFPLA_INST_0_45769 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_9[5]\, C => 
        \U50_PATTERNS/SM_BANK_SEL[10]\, Y => 
        HIEFFPLA_NET_0_118848);
    
    HIEFFPLA_INST_0_43229 : AND3B
      port map(A => HIEFFPLA_NET_0_119367, B => 
        HIEFFPLA_NET_0_119369, C => HIEFFPLA_NET_0_119355, Y => 
        HIEFFPLA_NET_0_119342);
    
    \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[14]\ : DFN1C0
      port map(D => \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\, 
        CLK => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[14]_net_1\);
    
    HIEFFPLA_INST_0_58491 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_31[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_15[1]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_3[4]_net_1\, Y
         => HIEFFPLA_NET_0_116515);
    
    \U_TFC_CMD_TX/SER_CMD_WORD_F[2]\ : DFN1C0
      port map(D => \U_TFC_CMD_TX/N_SER_CMD_WORD_F[2]\, CLK => 
        CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_TFC_CMD_TX/SER_CMD_WORD_F[2]_net_1\);
    
    \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_2S_2\ : DFN1C0
      port map(D => 
        \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_1S_net_1\, CLK
         => CLK60MHZ, CLR => P_MASTER_POR_B_c_0_0, Q => 
        P_USB_MASTER_EN_c_2);
    
    HIEFFPLA_INST_0_43604 : NAND3C
      port map(A => HIEFFPLA_NET_0_119273, B => 
        HIEFFPLA_NET_0_119252, C => HIEFFPLA_NET_0_119266, Y => 
        HIEFFPLA_NET_0_119270);
    
    HIEFFPLA_INST_0_53656 : MX2
      port map(A => HIEFFPLA_NET_0_117332, B => 
        HIEFFPLA_NET_0_117266, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[1]_net_1\, Y
         => HIEFFPLA_NET_0_117376);
    
    HIEFFPLA_INST_0_45066 : NAND3C
      port map(A => HIEFFPLA_NET_0_118987, B => 
        HIEFFPLA_NET_0_119471, C => HIEFFPLA_NET_0_119452, Y => 
        HIEFFPLA_NET_0_118988);
    
    HIEFFPLA_INST_0_59606 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_13[0]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_29[0]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_5[4]_net_1\, Y
         => HIEFFPLA_NET_0_116371);
    
    HIEFFPLA_INST_0_58777 : MX2
      port map(A => HIEFFPLA_NET_0_116687, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_19[2]\, S => 
        HIEFFPLA_NET_0_117205, Y => HIEFFPLA_NET_0_116477);
    
    HIEFFPLA_INST_0_56380 : AO1
      port map(A => HIEFFPLA_NET_0_117431, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[8]_net_1\, C => 
        HIEFFPLA_NET_0_116858, Y => HIEFFPLA_NET_0_116882);
    
    \U_ELK4_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]\ : DFN1C0
      port map(D => \U_ELK4_CH/U_SLAVE_1ELK/Q[4]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]_net_1\);
    
    HIEFFPLA_INST_0_50668 : MX2
      port map(A => \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\, B
         => \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\, S => 
        \BIT_OS_SEL_4[2]\, Y => HIEFFPLA_NET_0_117908);
    
    HIEFFPLA_INST_0_47082 : AND2
      port map(A => \U_ELK12_CH/ELK_TX_DAT[0]\, B => 
        \U_ELK12_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118562);
    
    \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[10]\ : DFN1C0
      port map(D => 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]_net_1\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\);
    
    HIEFFPLA_INST_0_45917 : AND3A
      port map(A => HIEFFPLA_NET_0_119376, B => 
        \U50_PATTERNS/TFC_STRT_ADDR[1]\, C => 
        HIEFFPLA_NET_0_119431, Y => HIEFFPLA_NET_0_118811);
    
    HIEFFPLA_INST_0_45682 : NAND2A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_4[6]\, Y => 
        HIEFFPLA_NET_0_118865);
    
    \U50_PATTERNS/ELINK_DINA_17[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119806, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_19, Q => 
        \U50_PATTERNS/ELINK_DINA_17[1]\);
    
    HIEFFPLA_INST_0_40015 : MX2
      port map(A => HIEFFPLA_NET_0_119896, B => 
        \U50_PATTERNS/ELINK_BLKA[1]\, S => 
        \U50_PATTERNS/SM_BANK_SEL_0[20]\, Y => 
        HIEFFPLA_NET_0_119924);
    
    HIEFFPLA_INST_0_41786 : MX2
      port map(A => HIEFFPLA_NET_0_119672, B => 
        \U50_PATTERNS/ELINK_RWA[6]\, S => 
        \U50_PATTERNS/SM_BANK_SEL_0[20]\, Y => 
        HIEFFPLA_NET_0_119695);
    
    HIEFFPLA_INST_0_37700 : AND3C
      port map(A => \U200B_ELINKS/GP_PG_SM[4]_net_1\, B => 
        \U200B_ELINKS/GP_PG_SM[5]_net_1\, C => 
        HIEFFPLA_NET_0_120234, Y => HIEFFPLA_NET_0_120226);
    
    \U_ELK11_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U0\ : IOPADP_BI
      port map(N2PIN => 
        \U_ELK11_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2_N2P\, D => 
        \U_ELK11_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, E => 
        \U_ELK11_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET2\, PAD => 
        ELK11_DAT_P, Y => 
        \U_ELK11_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\);
    
    HIEFFPLA_INST_0_43572 : AND2B
      port map(A => \U50_PATTERNS/SM_BANK_SEL_0[21]\, B => 
        \U50_PATTERNS/SM_BANK_SEL[6]\, Y => HIEFFPLA_NET_0_119285);
    
    HIEFFPLA_INST_0_49333 : MX2
      port map(A => 
        \U_ELK2_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]_net_1\, B => 
        \U_ELK2_CH/ELK_TX_DAT[4]\, S => 
        \U_ELK2_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118155);
    
    \U_ELK5_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0\ : DFN1C0
      port map(D => CLK_40M_GL, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_9, Q => 
        \U_ELK5_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0_net_1\);
    
    \U_ELK1_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]\ : DFN1C0
      port map(D => \U_ELK1_CH/U_SLAVE_1ELK/Q[6]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]_net_1\);
    
    HIEFFPLA_INST_0_46895 : MX2
      port map(A => HIEFFPLA_NET_0_118587, B => 
        HIEFFPLA_NET_0_118584, S => \BIT_OS_SEL_5[1]\, Y => 
        HIEFFPLA_NET_0_118588);
    
    HIEFFPLA_INST_0_47891 : MX2
      port map(A => \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[3]_net_1\, 
        B => \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\, S => 
        \BIT_OS_SEL_1[2]\, Y => HIEFFPLA_NET_0_118408);
    
    HIEFFPLA_INST_0_38106 : MX2
      port map(A => ELKS_RWB, B => \U200B_ELINKS/N_232_li\, S => 
        \U200B_ELINKS/GP_PG_SM[10]_net_1\, Y => 
        HIEFFPLA_NET_0_120151);
    
    HIEFFPLA_INST_0_50348 : MX2
      port map(A => 
        \U_ELK6_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]_net_1\, B => 
        \U_ELK6_CH/ELK_TX_DAT[5]\, S => 
        \U_ELK6_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_117971);
    
    \U_ELK2_CH/ELK_IN_R\ : DFN1C0
      port map(D => \U_ELK2_CH/ELK_IN_DDR_R\, CLK => CCC_160M_ADJ, 
        CLR => DEV_RST_B_c, Q => \U_ELK2_CH/ELK_IN_R_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_0[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116570, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_15, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_0[2]\);
    
    \U_ELK15_CH/U_SLAVE_1ELK/Q[13]\ : DFN1C0
      port map(D => \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[13]_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/Q[13]_net_1\);
    
    HIEFFPLA_INST_0_53302 : AND2A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_0[8]_net_1\, B => 
        HIEFFPLA_NET_0_116957, Y => HIEFFPLA_NET_0_117437);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_4[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116327, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_21, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_4[2]\);
    
    HIEFFPLA_INST_0_53022 : MX2
      port map(A => HIEFFPLA_NET_0_117455, B => 
        HIEFFPLA_NET_0_117567, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[2]\, Y => 
        HIEFFPLA_NET_0_117475);
    
    HIEFFPLA_INST_0_62128 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_2[3]\, 
        B => HIEFFPLA_NET_0_117186, S => HIEFFPLA_NET_0_117176, Y
         => HIEFFPLA_NET_0_116032);
    
    HIEFFPLA_INST_0_40990 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_19[4]\, B => 
        HIEFFPLA_NET_0_119570, S => HIEFFPLA_NET_0_119293, Y => 
        HIEFFPLA_NET_0_119787);
    
    HIEFFPLA_INST_0_37805 : NAND3
      port map(A => HIEFFPLA_NET_0_120190, B => 
        \U200B_ELINKS/GP_PG_SM[2]_net_1\, C => \OP_MODE_c[6]\, Y
         => HIEFFPLA_NET_0_120204);
    
    \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM[3]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM_0[4]_net_1\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_22, Q => 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM[3]_net_1\);
    
    HIEFFPLA_INST_0_61661 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_25[0]\, B => 
        HIEFFPLA_NET_0_117190, S => HIEFFPLA_NET_0_117117, Y => 
        HIEFFPLA_NET_0_116095);
    
    HIEFFPLA_INST_0_49933 : MX2
      port map(A => \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\, B
         => \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\, S => 
        \BIT_OS_SEL_6[2]\, Y => HIEFFPLA_NET_0_118041);
    
    HIEFFPLA_INST_0_47092 : MX2
      port map(A => 
        \U_ELK12_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]_net_1\, B => 
        \U_ELK12_CH/ELK_TX_DAT[4]\, S => 
        \U_ELK12_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118560);
    
    \U_MASTER_DES/U13C_MASTER_DESER/ARB_WRD_40M_FIXED[14]\ : 
        DFN1C0
      port map(D => \U_MASTER_DES/U13C_MASTER_DESER/Q[14]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_28, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_WRD_40M_FIXED[14]_net_1\);
    
    \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[14]\ : DFN1C0
      port map(D => \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\, 
        CLK => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[14]_net_1\);
    
    \U_ELK0_SERDAT_SOURCE/SERDAT[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118660, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_10, Q => \ELK0_TX_DAT[0]\);
    
    HIEFFPLA_INST_0_54569 : AND2A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[2]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[4]_net_1\, Y => 
        HIEFFPLA_NET_0_117244);
    
    \U_ELK12_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118559, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_15, Q => 
        \U_ELK12_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]_net_1\);
    
    HIEFFPLA_INST_0_47449 : MX2
      port map(A => HIEFFPLA_NET_0_118500, B => 
        HIEFFPLA_NET_0_118497, S => \BIT_OS_SEL_3[1]\, Y => 
        HIEFFPLA_NET_0_118490);
    
    HIEFFPLA_INST_0_61538 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_7[3]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_23[3]\, S
         => \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[4]_net_1\, 
        Y => HIEFFPLA_NET_0_116113);
    
    HIEFFPLA_INST_0_41026 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_1[0]\, B => 
        HIEFFPLA_NET_0_119578, S => HIEFFPLA_NET_0_119243, Y => 
        HIEFFPLA_NET_0_119783);
    
    \U50_PATTERNS/SM_BANK_SEL[14]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119317, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_1_0, Q => 
        \U50_PATTERNS/SM_BANK_SEL[14]\);
    
    HIEFFPLA_INST_0_61586 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_24[0]\, B => 
        HIEFFPLA_NET_0_117190, S => HIEFFPLA_NET_0_117074, Y => 
        HIEFFPLA_NET_0_116105);
    
    HIEFFPLA_INST_0_37683 : AND3
      port map(A => HIEFFPLA_NET_0_120226, B => 
        HIEFFPLA_NET_0_120224, C => HIEFFPLA_NET_0_120225, Y => 
        HIEFFPLA_NET_0_120230);
    
    HIEFFPLA_INST_0_48122 : AND2A
      port map(A => \OP_MODE_c_2[1]\, B => \PATT_ELK_DAT_16[5]\, 
        Y => HIEFFPLA_NET_0_118368);
    
    \U_ELK5_CH/U_SLAVE_1ELK/Q[10]\ : DFN1C0
      port map(D => \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/Q[10]_net_1\);
    
    HIEFFPLA_INST_0_43449 : MX2
      port map(A => \U50_PATTERNS/SM_BANK_SEL[20]\, B => 
        HIEFFPLA_NET_0_119467, S => HIEFFPLA_NET_0_118691, Y => 
        HIEFFPLA_NET_0_119310);
    
    \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[7]\ : DFN1C0
      port map(D => \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\);
    
    HIEFFPLA_INST_0_37156 : XO1
      port map(A => \TFC_ADDRB[5]\, B => HIEFFPLA_NET_0_120260, C
         => \U200A_TFC/GP_PG_SM[10]_net_1\, Y => 
        HIEFFPLA_NET_0_120338);
    
    HIEFFPLA_INST_0_51673 : AND2B
      port map(A => \U_GEN_REF_CLK/GEN_40M_REFCNT[2]_net_1\, B
         => \U_GEN_REF_CLK/GEN_40M_REFCNT[1]_net_1\, Y => 
        HIEFFPLA_NET_0_117728);
    
    \U_ELK6_CH/U_SLAVE_1ELK/Q[2]\ : DFN1C0
      port map(D => \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/Q[2]_net_1\);
    
    HIEFFPLA_INST_0_58763 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_19[2]\, B => 
        HIEFFPLA_NET_0_116477, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_2[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116479);
    
    HIEFFPLA_INST_0_56375 : AO1
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[7]_net_1\, B => 
        HIEFFPLA_NET_0_117431, C => HIEFFPLA_NET_0_116859, Y => 
        HIEFFPLA_NET_0_116883);
    
    HIEFFPLA_INST_0_43566 : NAND2B
      port map(A => \U50_PATTERNS/SM_BANK_SEL[21]\, B => 
        \U50_PATTERNS/SM_BANK_SEL[12]\, Y => 
        HIEFFPLA_NET_0_119289);
    
    HIEFFPLA_INST_0_48848 : MX2
      port map(A => 
        \U_ELK19_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]_net_1\, B => 
        \U_ELK19_CH/ELK_TX_DAT[3]\, S => 
        \U_ELK19_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118242);
    
    HIEFFPLA_INST_0_45863 : AO1
      port map(A => HIEFFPLA_NET_0_119283, B => 
        \U50_PATTERNS/ELINK_DOUTA_13[3]\, C => 
        HIEFFPLA_NET_0_118778, Y => HIEFFPLA_NET_0_118825);
    
    HIEFFPLA_INST_0_41793 : MX2
      port map(A => HIEFFPLA_NET_0_119670, B => 
        \U50_PATTERNS/ELINK_RWA[7]\, S => 
        \U50_PATTERNS/SM_BANK_SEL_0[20]\, Y => 
        HIEFFPLA_NET_0_119694);
    
    \U_ELK11_CH/U_ELK1_SERDAT_SOURCE/SERDAT[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118597, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_0, Q => 
        \U_ELK11_CH/ELK_TX_DAT[1]\);
    
    HIEFFPLA_INST_0_57676 : AND3B
      port map(A => HIEFFPLA_NET_0_116633, B => 
        HIEFFPLA_NET_0_117179, C => HIEFFPLA_NET_0_116651, Y => 
        HIEFFPLA_NET_0_116637);
    
    HIEFFPLA_INST_0_46945 : MX2
      port map(A => \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\, 
        B => \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[12]_net_1\, S => 
        \BIT_OS_SEL_5[2]\, Y => HIEFFPLA_NET_0_118581);
    
    HIEFFPLA_INST_0_42002 : AO1A
      port map(A => \U50_PATTERNS/REG_STATE[5]_net_1\, B => 
        HIEFFPLA_NET_0_119380, C => HIEFFPLA_NET_0_119004, Y => 
        HIEFFPLA_NET_0_119634);
    
    HIEFFPLA_INST_0_58234 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_12[1]\, B => 
        HIEFFPLA_NET_0_116677, S => HIEFFPLA_NET_0_117089, Y => 
        HIEFFPLA_NET_0_116547);
    
    \U_EXEC_MASTER/MPOR_B_5\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117787, CLK => CLK_40M_GL, CLR
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_1\, Q => 
        P_MASTER_POR_B_c_5);
    
    HIEFFPLA_INST_0_60402 : MX2
      port map(A => HIEFFPLA_NET_0_117100, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_10[4]\, S => 
        HIEFFPLA_NET_0_117154, Y => HIEFFPLA_NET_0_116271);
    
    HIEFFPLA_INST_0_52232 : AND3A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[6]_net_1\, B => 
        HIEFFPLA_NET_0_117581, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[1]_net_1\, Y => 
        HIEFFPLA_NET_0_117604);
    
    \U_ELK4_CH/U_SLAVE_1ELK/RECD_SER_WORD[0]\ : DFN1C0
      port map(D => \U_ELK4_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[0]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_4[0]\);
    
    \U_ELK14_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]\ : DFN1C0
      port map(D => \U_ELK14_CH/U_SLAVE_1ELK/Q[4]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]_net_1\);
    
    HIEFFPLA_INST_0_37693 : AND2B
      port map(A => \U200B_ELINKS/GP_PG_SM[6]_net_1\, B => 
        \U200B_ELINKS/GP_PG_SM[7]_net_1\, Y => 
        HIEFFPLA_NET_0_120228);
    
    \U_ELK9_CH/U_SLAVE_1ELK/Q[13]\ : DFN1C0
      port map(D => \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[13]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/Q[13]_net_1\);
    
    HIEFFPLA_INST_0_52836 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_15[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_16[1]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_2[0]\, Y => 
        HIEFFPLA_NET_0_117503);
    
    HIEFFPLA_INST_0_41932 : NAND2
      port map(A => HIEFFPLA_NET_0_119389, B => 
        \U50_PATTERNS/SM_BANK_SEL[5]\, Y => HIEFFPLA_NET_0_119656);
    
    \U_MASTER_DES/U13C_MASTER_DESER/BEST_BIT_OS_VAL[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_117580, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_13, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_BIT_OS_VAL[0]\);
    
    \U50_PATTERNS/ELINK_DINA_11[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119850, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_11, Q => 
        \U50_PATTERNS/ELINK_DINA_11[5]\);
    
    HIEFFPLA_INST_0_49917 : MX2
      port map(A => HIEFFPLA_NET_0_118045, B => 
        HIEFFPLA_NET_0_118041, S => \BIT_OS_SEL_6[1]\, Y => 
        HIEFFPLA_NET_0_118043);
    
    HIEFFPLA_INST_0_45652 : NAND3C
      port map(A => HIEFFPLA_NET_0_118717, B => 
        HIEFFPLA_NET_0_118890, C => HIEFFPLA_NET_0_118705, Y => 
        HIEFFPLA_NET_0_118872);
    
    \U_ELK3_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]\ : DFN1C0
      port map(D => \U_ELK3_CH/U_SLAVE_1ELK/Q[4]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]_net_1\);
    
    HIEFFPLA_INST_0_61346 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_5[4]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_21[4]\, S
         => \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_1[4]_net_1\, 
        Y => HIEFFPLA_NET_0_116140);
    
    HIEFFPLA_INST_0_48337 : MX2
      port map(A => 
        \U_ELK17_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]_net_1\, B => 
        \U_ELK17_CH/ELK_TX_DAT[4]\, S => 
        \U_ELK17_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118335);
    
    \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[12]\ : DFN1C0
      port map(D => 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]_net_1\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[12]_net_1\);
    
    \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[4]\ : DFN1C0
      port map(D => 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\);
    
    \U_ELK10_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U1\ : IOBI_ID_OD_EB
      port map(DR => \U_ELK10_CH/ELK_OUT_R\, DF => 
        \U_ELK10_CH/ELK_OUT_F\, CLR => \GND\, E => 
        \AFLSDF_INV_14\, ICLK => CCC_160M_ADJ, OCLK => 
        CCC_160M_FXD, YIN => 
        \U_ELK10_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\, DOUT => 
        \U_ELK10_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, EOUT => 
        \U_ELK10_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET2\, YR => 
        \U_ELK10_CH/ELK_IN_DDR_R\, YF => 
        \U_ELK10_CH/ELK_IN_DDR_F\);
    
    HIEFFPLA_INST_0_53730 : MX2
      port map(A => HIEFFPLA_NET_0_117324, B => 
        HIEFFPLA_NET_0_117304, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[2]_net_1\, Y
         => HIEFFPLA_NET_0_117363);
    
    HIEFFPLA_INST_0_38056 : AOI1A
      port map(A => HIEFFPLA_NET_0_120229, B => 
        HIEFFPLA_NET_0_120220, C => HIEFFPLA_NET_0_120163, Y => 
        HIEFFPLA_NET_0_120164);
    
    \U_DDR_ELK0/BIBUF_LVDS_0/U0/U3\ : IOBI_ID_OD_EB
      port map(DR => ELK0_OUT_R_i_0, DF => ELK0_OUT_F_i_0, CLR
         => \GND\, E => \AFLSDF_INV_13\, ICLK => CCC_160M_ADJ, 
        OCLK => CCC_160M_FXD, YIN => 
        \U_DDR_ELK0/BIBUF_LVDS_0/U0/NET4\, DOUT => OPEN, EOUT => 
        \U_DDR_ELK0/BIBUF_LVDS_0/U0/NET3\, YR => OPEN, YF => OPEN);
    
    \U50_PATTERNS/TFC_STOP_ADDR[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119181, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_8, Q => 
        \U50_PATTERNS/TFC_STOP_ADDR[7]\);
    
    HIEFFPLA_INST_0_54998 : OA1A
      port map(A => HIEFFPLA_NET_0_117242, B => 
        HIEFFPLA_NET_0_117247, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_3[6]_net_1\, Y => 
        HIEFFPLA_NET_0_117145);
    
    \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[2]\ : DFN1C0
      port map(D => \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\);
    
    \U_ELK17_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]\ : DFN1C0
      port map(D => \U_ELK17_CH/U_SLAVE_1ELK/Q[2]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]_net_1\);
    
    \U200A_TFC/RX_SER_WORD_2DEL[0]\ : DFN1C0
      port map(D => \U200A_TFC/RX_SER_WORD_1DEL[0]_net_1\, CLK
         => CLK_40M_GL, CLR => P_MASTER_POR_B_c, Q => 
        \U200A_TFC/RX_SER_WORD_2DEL[0]_net_1\);
    
    \U_ELK4_CH/U_ELK1_SERDAT_SOURCE/SERDAT[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118058, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_16, Q => 
        \U_ELK4_CH/ELK_TX_DAT[0]\);
    
    HIEFFPLA_INST_0_39722 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_7[0]\, B => 
        HIEFFPLA_NET_0_119524, S => HIEFFPLA_NET_0_119289, Y => 
        HIEFFPLA_NET_0_119959);
    
    HIEFFPLA_INST_0_61121 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_1[0]\, 
        B => HIEFFPLA_NET_0_117190, S => HIEFFPLA_NET_0_117149, Y
         => HIEFFPLA_NET_0_116170);
    
    \U200A_TFC/RX_SER_WORD_1DEL[7]\ : DFN1C0
      port map(D => \TFC_RX_SER_WORD[7]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_31, Q => 
        \U200A_TFC/RX_SER_WORD_1DEL[7]_net_1\);
    
    HIEFFPLA_INST_0_62780 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/TUNE_CLKPHASE[1]\, B => 
        HIEFFPLA_NET_0_115957, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[1]_net_1\, Y => 
        HIEFFPLA_NET_0_115948);
    
    HIEFFPLA_INST_0_53541 : MX2
      port map(A => HIEFFPLA_NET_0_117333, B => 
        HIEFFPLA_NET_0_117311, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[0]_net_1\, Y
         => HIEFFPLA_NET_0_117391);
    
    \U60_TS_RD_BUF/_TRIBUFF_F_24U[0]_/U0/U1\ : IOTRI_OB_EB
      port map(D => USB_RD_BI, E => P_USB_MASTER_EN_c, DOUT => 
        \U60_TS_RD_BUF/\\\\TRIBUFF_F_24U[0]\\\\/U0/NET1\, EOUT
         => \U60_TS_RD_BUF/\\\\TRIBUFF_F_24U[0]\\\\/U0/NET2\);
    
    \U50_PATTERNS/ELINK_BLKA[2]/U1\ : DFN1P0
      port map(D => HIEFFPLA_NET_0_119923, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_19, Q => 
        \U50_PATTERNS/ELINK_BLKA[2]\);
    
    HIEFFPLA_INST_0_53198 : MX2
      port map(A => HIEFFPLA_NET_0_117529, B => 
        HIEFFPLA_NET_0_117521, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[3]\, Y => 
        HIEFFPLA_NET_0_117453);
    
    HIEFFPLA_INST_0_53134 : MX2
      port map(A => HIEFFPLA_NET_0_117545, B => 
        HIEFFPLA_NET_0_117541, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[3]\, Y => 
        HIEFFPLA_NET_0_117461);
    
    HIEFFPLA_INST_0_44880 : OA1A
      port map(A => \U50_PATTERNS/USB_RXF_B\, B => 
        HIEFFPLA_NET_0_119479, C => 
        \U50_PATTERNS/REG_STATE_0[4]_net_1\, Y => 
        HIEFFPLA_NET_0_119029);
    
    HIEFFPLA_INST_0_63156 : AX1C
      port map(A => HIEFFPLA_NET_0_115874, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[3]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[4]\, Y => 
        HIEFFPLA_NET_0_115873);
    
    HIEFFPLA_INST_0_60197 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_7[2]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_23[2]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_4[4]_net_1\, Y
         => HIEFFPLA_NET_0_116297);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_24[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116432, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_18, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_24[2]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_12[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116545, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_10, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_12[3]\);
    
    \U_EXEC_MASTER/USB_MASTER_EN/TEST_SM[0]\ : DFN1P0
      port map(D => \GND\, CLK => CLK_40M_GL, PRE => 
        P_MASTER_POR_B_c_24, Q => 
        \U_EXEC_MASTER/USB_MASTER_EN/TEST_SM[0]_net_1\);
    
    \U_EXEC_MASTER/DEL_CNT[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117791, CLK => CLK_40M_GL, CLR
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i\, Q => 
        \U_EXEC_MASTER/DEL_CNT[4]\);
    
    HIEFFPLA_INST_0_50937 : MX2
      port map(A => HIEFFPLA_NET_0_117862, B => 
        HIEFFPLA_NET_0_117858, S => \BIT_OS_SEL_3[1]\, Y => 
        HIEFFPLA_NET_0_117860);
    
    HIEFFPLA_INST_0_41823 : AOI1B
      port map(A => HIEFFPLA_NET_0_119389, B => 
        \U50_PATTERNS/SM_BANK_SEL[8]\, C => HIEFFPLA_NET_0_119661, 
        Y => HIEFFPLA_NET_0_119689);
    
    HIEFFPLA_INST_0_38073 : NAND3C
      port map(A => HIEFFPLA_NET_0_120161, B => 
        \U200B_ELINKS/RX_SER_WORD_2DEL[5]_net_1\, C => 
        HIEFFPLA_NET_0_120162, Y => HIEFFPLA_NET_0_120159);
    
    \U_ELK14_CH/U_SLAVE_1ELK/RECD_SER_WORD[0]\ : DFN1C0
      port map(D => \U_ELK14_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[0]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_14[0]\);
    
    \U_ELK10_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118646, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_3, Q => 
        \U_ELK10_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]_net_1\);
    
    HIEFFPLA_INST_0_51106 : NAND2B
      port map(A => \OP_MODE_c_3[1]\, B => \PATT_ELK_DAT_9[1]\, Y
         => HIEFFPLA_NET_0_117832);
    
    HIEFFPLA_INST_0_44384 : MX2
      port map(A => \TFC_STOP_ADDR[5]\, B => 
        \U50_PATTERNS/U4B_REGCROSS/SAMP_TWO[5]_net_1\, S => 
        HIEFFPLA_NET_0_119135, Y => HIEFFPLA_NET_0_119128);
    
    \U50_PATTERNS/OP_MODE_T[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119609, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_17, Q => 
        \U50_PATTERNS/OP_MODE_T[0]\);
    
    HIEFFPLA_INST_0_57328 : AOI1
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_3[0]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_3[1]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_3[2]\, Y => 
        HIEFFPLA_NET_0_116698);
    
    \U_ELK14_CH/U_SLAVE_1ELK/RECD_SER_WORD[1]\ : DFN1C0
      port map(D => \U_ELK14_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[1]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_14[1]\);
    
    HIEFFPLA_INST_0_55707 : MX2
      port map(A => HIEFFPLA_NET_0_115972, B => 
        HIEFFPLA_NET_0_116225, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_2[3]\, Y => 
        HIEFFPLA_NET_0_117001);
    
    \U_ELK4_CH/U_SLAVE_1ELK/Q[13]\ : DFN1C0
      port map(D => \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[13]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/Q[13]_net_1\);
    
    HIEFFPLA_INST_0_44718 : MX2
      port map(A => \OP_MODE_c_0[1]\, B => 
        \U50_PATTERNS/U4E_REGCROSS/SAMP_TWO[1]_net_1\, S => 
        HIEFFPLA_NET_0_119072, Y => HIEFFPLA_NET_0_119062);
    
    HIEFFPLA_INST_0_37722 : AND3C
      port map(A => \U200B_ELINKS/GP_PG_SM[2]_net_1\, B => 
        \U200B_ELINKS/GP_PG_SM[3]_net_1\, C => 
        \U200B_ELINKS/GP_PG_SM[0]_net_1\, Y => 
        HIEFFPLA_NET_0_120222);
    
    HIEFFPLA_INST_0_42677 : AND3A
      port map(A => HIEFFPLA_NET_0_118996, B => 
        HIEFFPLA_NET_0_119369, C => 
        \U50_PATTERNS/REG_STATE_0[5]_net_1\, Y => 
        HIEFFPLA_NET_0_119485);
    
    HIEFFPLA_INST_0_45523 : AO1A
      port map(A => HIEFFPLA_NET_0_119428, B => 
        \U50_PATTERNS/ELINKS_STRT_ADDR[0]\, C => 
        HIEFFPLA_NET_0_118794, Y => HIEFFPLA_NET_0_118897);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_16[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116509, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_16_0, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_16[3]\);
    
    HIEFFPLA_INST_0_37314 : NAND3A
      port map(A => \U200A_TFC/GP_PG_SM[4]_net_1\, B => 
        \U200A_TFC/GP_PG_SM[5]_net_1\, C => HIEFFPLA_NET_0_120326, 
        Y => HIEFFPLA_NET_0_120297);
    
    \U_ELK10_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118648, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_3, Q => 
        \U_ELK10_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]_net_1\);
    
    HIEFFPLA_INST_0_54924 : AO1C
      port map(A => HIEFFPLA_NET_0_117107, B => 
        HIEFFPLA_NET_0_117209, C => HIEFFPLA_NET_0_117180, Y => 
        HIEFFPLA_NET_0_117169);
    
    \U_ELK3_CH/U_ELK1_CMD_TX/SER_OUT_RI\ : DFI1C0
      port map(D => 
        \U_ELK3_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_14, QN
         => \U_ELK3_CH/U_ELK1_CMD_TX/SER_OUT_RI_i\);
    
    \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[7]\ : DFN1C0
      port map(D => \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\);
    
    HIEFFPLA_INST_0_55179 : AO1E
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[3]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[2]_net_1\, C => 
        \U_MASTER_DES/CCC_RX_CLK_LOCK\, Y => 
        HIEFFPLA_NET_0_117103);
    
    \U200B_ELINKS/ADDR_POINTER[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120169, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_31_0, Q => \ELKS_ADDRB[2]\);
    
    HIEFFPLA_INST_0_59954 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_4[0]\, B => 
        HIEFFPLA_NET_0_116680, S => HIEFFPLA_NET_0_117155, Y => 
        HIEFFPLA_NET_0_116329);
    
    \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[40]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117712, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_33, Q => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[40]_net_1\);
    
    \U_ELK8_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2\ : IOPADN_BI
      port map(DB => \U_ELK8_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, 
        E => \U_ELK8_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET3\, PAD => 
        ELK8_DAT_N, N2POUT => 
        \U_ELK8_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2_N2P\);
    
    \U_ELK7_CH/ELK_IN_R\ : DFN1C0
      port map(D => \U_ELK7_CH/ELK_IN_DDR_R\, CLK => CCC_160M_ADJ, 
        CLR => DEV_RST_B_c, Q => \U_ELK7_CH/ELK_IN_R_net_1\);
    
    \U_ELK3_CH/U_SLAVE_1ELK/RECD_SER_WORD[4]\ : DFN1C0
      port map(D => \U_ELK3_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[4]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_3[4]\);
    
    HIEFFPLA_INST_0_48660 : MX2
      port map(A => \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\, 
        B => \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\, S => 
        \BIT_OS_SEL_0[2]\, Y => HIEFFPLA_NET_0_118270);
    
    HIEFFPLA_INST_0_111787 : AND2B
      port map(A => HIEFFPLA_NET_0_115832, B => 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM[6]_net_1\, Y => 
        HIEFFPLA_NET_0_117670);
    
    HIEFFPLA_INST_0_43593 : NAND2B
      port map(A => \U50_PATTERNS/SM_BANK_SEL[9]\, B => 
        \U50_PATTERNS/SM_BANK_SEL[4]\, Y => HIEFFPLA_NET_0_119274);
    
    HIEFFPLA_INST_0_42881 : NAND2
      port map(A => \U50_PATTERNS/REG_STATE[4]_net_1\, B => 
        \U50_PATTERNS/REG_STATE[2]_net_1\, Y => 
        HIEFFPLA_NET_0_119437);
    
    \U_ELK8_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U3\ : IOBI_ID_OD_EB
      port map(DR => \U_ELK8_CH/ELK_OUT_R\, DF => 
        \U_ELK8_CH/ELK_OUT_F\, CLR => \GND\, E => \AFLSDF_INV_49\, 
        ICLK => CCC_160M_ADJ, OCLK => CCC_160M_FXD, YIN => 
        \U_ELK8_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\, DOUT => OPEN, 
        EOUT => \U_ELK8_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET3\, YR
         => OPEN, YF => OPEN);
    
    \U50_PATTERNS/U4E_REGCROSS/SAMP_ONE[7]\ : DFN1C0
      port map(D => \U50_PATTERNS/OP_MODE[7]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c, Q => 
        \U50_PATTERNS/U4E_REGCROSS/SAMP_ONE[7]_net_1\);
    
    \U50_PATTERNS/ELINK_ADDRA_9[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119936, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_10, Q => 
        \U50_PATTERNS/ELINK_ADDRA_9[7]\);
    
    \U50_PATTERNS/ELINK_DINA_3[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119766, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_11, Q => 
        \U50_PATTERNS/ELINK_DINA_3[1]\);
    
    \U50_PATTERNS/ELINK_DINA_3[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119765, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_11, Q => 
        \U50_PATTERNS/ELINK_DINA_3[2]\);
    
    HIEFFPLA_INST_0_39182 : MX2
      port map(A => HIEFFPLA_NET_0_119519, B => 
        \U50_PATTERNS/ELINK_ADDRA_18[4]\, S => 
        HIEFFPLA_NET_0_119264, Y => HIEFFPLA_NET_0_120019);
    
    HIEFFPLA_INST_0_54808 : MX2
      port map(A => HIEFFPLA_NET_0_117300, B => 
        HIEFFPLA_NET_0_117274, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[2]_net_1\, Y => 
        HIEFFPLA_NET_0_117197);
    
    \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_2S_0\ : DFN1C0
      port map(D => 
        \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_1S_net_1\, CLK
         => CLK60MHZ, CLR => P_MASTER_POR_B_c_0_0, Q => 
        P_USB_MASTER_EN_c_0);
    
    HIEFFPLA_INST_0_56029 : MX2
      port map(A => HIEFFPLA_NET_0_116980, B => 
        HIEFFPLA_NET_0_117002, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[2]\, Y => 
        HIEFFPLA_NET_0_116959);
    
    HIEFFPLA_INST_0_55890 : MX2
      port map(A => HIEFFPLA_NET_0_116990, B => 
        HIEFFPLA_NET_0_116963, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[1]\, Y => 
        HIEFFPLA_NET_0_116977);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_19[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116479, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_20, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_19[2]\);
    
    \U_ELK16_CH/ELK_IN_R\ : DFN1C0
      port map(D => \U_ELK16_CH/ELK_IN_DDR_R\, CLK => 
        CCC_160M_ADJ, CLR => DEV_RST_B_c, Q => 
        \U_ELK16_CH/ELK_IN_R_net_1\);
    
    \U_EXEC_MASTER/DEL_CNT[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117794, CLK => CLK_40M_GL, CLR
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i\, Q => 
        \U_EXEC_MASTER/DEL_CNT[1]\);
    
    HIEFFPLA_INST_0_53555 : NAND3C
      port map(A => HIEFFPLA_NET_0_117378, B => 
        HIEFFPLA_NET_0_117070, C => HIEFFPLA_NET_0_117127, Y => 
        HIEFFPLA_NET_0_117389);
    
    HIEFFPLA_INST_0_48117 : AND2A
      port map(A => \OP_MODE_c_2[1]\, B => \PATT_ELK_DAT_16[0]\, 
        Y => HIEFFPLA_NET_0_118373);
    
    HIEFFPLA_INST_0_47274 : MX2
      port map(A => HIEFFPLA_NET_0_118545, B => 
        HIEFFPLA_NET_0_118542, S => \BIT_OS_SEL_5[0]\, Y => 
        \U_ELK12_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[4]\);
    
    HIEFFPLA_INST_0_52416 : MX2
      port map(A => HIEFFPLA_NET_0_117518, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_29[2]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[3]\, Y => 
        HIEFFPLA_NET_0_117566);
    
    HIEFFPLA_INST_0_39011 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_16[1]\, B => 
        HIEFFPLA_NET_0_119523, S => HIEFFPLA_NET_0_119257, Y => 
        HIEFFPLA_NET_0_120038);
    
    HIEFFPLA_INST_0_49796 : MX2
      port map(A => HIEFFPLA_NET_0_118069, B => 
        HIEFFPLA_NET_0_118094, S => \BIT_OS_SEL_6[1]\, Y => 
        HIEFFPLA_NET_0_118071);
    
    HIEFFPLA_INST_0_38410 : MX2
      port map(A => \U50_PATTERNS/ELINKS_STRT_ADDR[5]\, B => 
        \U50_PATTERNS/ELINKS_STRT_ADDR_T[5]\, S => 
        HIEFFPLA_NET_0_119472, Y => HIEFFPLA_NET_0_120106);
    
    \U50_PATTERNS/ELINK_ADDRA_7[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119955, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_6, Q => 
        \U50_PATTERNS/ELINK_ADDRA_7[4]\);
    
    \U_ELK6_CH/U_SLAVE_1ELK/Q[11]\ : DFN1C0
      port map(D => \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/Q[11]_net_1\);
    
    \U_ELK12_CH/U_SLAVE_1ELK/Q[10]\ : DFN1C0
      port map(D => \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/Q[10]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[8]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_WRD_40M_FIXED[8]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_27, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[8]_net_1\);
    
    HIEFFPLA_INST_0_61898 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_11[2]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_27[2]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_2[4]_net_1\, Y
         => HIEFFPLA_NET_0_116063);
    
    \U50_PATTERNS/U4B_REGCROSS/LOCAL_REG_VAL[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119128, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_19, Q => \TFC_STOP_ADDR[5]\);
    
    HIEFFPLA_INST_0_55604 : MX2
      port map(A => HIEFFPLA_NET_0_116195, B => 
        HIEFFPLA_NET_0_116087, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_1[3]\, Y => 
        HIEFFPLA_NET_0_117015);
    
    HIEFFPLA_INST_0_44536 : XO1
      port map(A => \ELKS_STRT_ADDR[4]\, B => 
        \U50_PATTERNS/U4C_REGCROSS/SAMP_TWO[4]_net_1\, C => 
        HIEFFPLA_NET_0_119096, Y => HIEFFPLA_NET_0_119099);
    
    HIEFFPLA_INST_0_43033 : AO1
      port map(A => HIEFFPLA_NET_0_119430, B => 
        HIEFFPLA_NET_0_119414, C => HIEFFPLA_NET_0_119395, Y => 
        HIEFFPLA_NET_0_119396);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_25[4]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116091, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_10, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_25[4]\);
    
    \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_2S_22_0\ : DFN1C0
      port map(D => 
        \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_1S_0_net_1\, CLK
         => CLK60MHZ, CLR => P_MASTER_POR_B_c_0_0, Q => 
        P_USB_MASTER_EN_c_22_0);
    
    \U_ELK2_CH/U_ELK1_CMD_TX/SER_OUT_RI\ : DFN1C0
      port map(D => 
        \U_ELK2_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_5, Q => 
        \U_ELK2_CH/U_ELK1_CMD_TX/SER_OUT_RI_net_1\);
    
    HIEFFPLA_INST_0_43273 : AXOI4
      port map(A => HIEFFPLA_NET_0_119329, B => 
        HIEFFPLA_NET_0_119439, C => \U50_PATTERNS/SI_CNT[0]\, Y
         => HIEFFPLA_NET_0_119334);
    
    HIEFFPLA_INST_0_62298 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_3[3]\, 
        B => HIEFFPLA_NET_0_117075, S => HIEFFPLA_NET_0_117178, Y
         => HIEFFPLA_NET_0_116007);
    
    \U_ELK1_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118201, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_7, Q => 
        \U_ELK1_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]_net_1\);
    
    HIEFFPLA_INST_0_111899 : AOI1
      port map(A => HIEFFPLA_NET_0_115824, B => 
        \U50_PATTERNS/REG_STATE[2]_net_1\, C => 
        HIEFFPLA_NET_0_119473, Y => HIEFFPLA_NET_0_119018);
    
    \U_ELK0_CMD_TX/SER_CMD_WORD_R[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118662, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_14, Q => 
        \U_ELK0_CMD_TX/SER_CMD_WORD_R[3]_net_1\);
    
    \U50_PATTERNS/ELINK_DINA_15[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119817, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_16, Q => 
        \U50_PATTERNS/ELINK_DINA_15[6]\);
    
    HIEFFPLA_INST_0_52702 : MX2
      port map(A => HIEFFPLA_NET_0_117477, B => 
        HIEFFPLA_NET_0_117473, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[4]\, Y => 
        HIEFFPLA_NET_0_117525);
    
    HIEFFPLA_INST_0_45712 : NAND2A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_4[0]\, Y => 
        HIEFFPLA_NET_0_118860);
    
    \U200B_ELINKS/RX_SER_WORD_2DEL[4]\ : DFN1C0
      port map(D => \U200B_ELINKS/RX_SER_WORD_1DEL[4]_net_1\, CLK
         => CLK_40M_GL, CLR => P_MASTER_POR_B_c_25, Q => 
        \U200B_ELINKS/RX_SER_WORD_2DEL[4]_net_1\);
    
    \U50_PATTERNS/CHKSUM[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120139, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_3, Q => \U50_PATTERNS/CHKSUM[4]\);
    
    HIEFFPLA_INST_0_42791 : AND3A
      port map(A => HIEFFPLA_NET_0_119432, B => 
        HIEFFPLA_NET_0_119466, C => 
        \U50_PATTERNS/REG_STATE_0[4]_net_1\, Y => 
        HIEFFPLA_NET_0_119462);
    
    HIEFFPLA_INST_0_53829 : MX2
      port map(A => HIEFFPLA_NET_0_116124, B => 
        HIEFFPLA_NET_0_116022, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[3]_net_1\, Y
         => HIEFFPLA_NET_0_117346);
    
    \U50_PATTERNS/ELINK_ADDRA_12[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120069, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_2_0, Q => 
        \U50_PATTERNS/ELINK_ADDRA_12[2]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_15[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116229, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_4, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_15[1]\);
    
    HIEFFPLA_INST_0_49407 : MX2
      port map(A => \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\, B
         => \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\, S => 
        \BIT_OS_SEL_7[2]\, Y => HIEFFPLA_NET_0_118135);
    
    HIEFFPLA_INST_0_41017 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_19[7]\, B => 
        HIEFFPLA_NET_0_119560, S => HIEFFPLA_NET_0_119293, Y => 
        HIEFFPLA_NET_0_119784);
    
    \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[7]\ : DFN1C0
      port map(D => \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\);
    
    \U50_PATTERNS/TFC_STOP_ADDR_T[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119177, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_15, Q => 
        \U50_PATTERNS/TFC_STOP_ADDR_T[3]\);
    
    \U50_PATTERNS/RD_XFER_TYPE[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119548, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c, Q => 
        \U50_PATTERNS/RD_XFER_TYPE[1]_net_1\);
    
    HIEFFPLA_INST_0_48744 : MX2
      port map(A => HIEFFPLA_NET_0_118264, B => 
        HIEFFPLA_NET_0_118260, S => \BIT_OS_SEL_2[0]\, Y => 
        \U_ELK18_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[1]\);
    
    HIEFFPLA_INST_0_47381 : MX2
      port map(A => \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[2]_net_1\, 
        B => \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\, S => 
        \BIT_OS_SEL_2[2]\, Y => HIEFFPLA_NET_0_118500);
    
    HIEFFPLA_INST_0_46600 : MX2
      port map(A => 
        \U_ELK10_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]_net_1\, B => 
        \U_ELK10_CH/ELK_TX_DAT[6]\, S => 
        \U_ELK10_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118649);
    
    HIEFFPLA_INST_0_60093 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_6[3]\, B => 
        HIEFFPLA_NET_0_116307, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_0[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116311);
    
    HIEFFPLA_INST_0_49607 : MX2
      port map(A => 
        \U_ELK3_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]_net_1\, B => 
        \U_ELK3_CH/ELK_TX_DAT[7]\, S => 
        \U_ELK3_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118105);
    
    HIEFFPLA_INST_0_38040 : AND3B
      port map(A => \U200B_ELINKS/LOC_STRT_ADDR[2]\, B => 
        HIEFFPLA_NET_0_120190, C => HIEFFPLA_NET_0_120234, Y => 
        HIEFFPLA_NET_0_120167);
    
    HIEFFPLA_INST_0_50342 : MX2
      port map(A => 
        \U_ELK6_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]_net_1\, B => 
        \U_ELK6_CH/ELK_TX_DAT[3]\, S => 
        \U_ELK6_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_117972);
    
    AFLSDF_INV_38 : INV
      port map(A => DCB_SALT_SEL_c, Y => \AFLSDF_INV_38\);
    
    \U_ELK8_CH/U_ELK1_SERDAT_SOURCE/SERDAT[6]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117872, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_5, Q => 
        \U_ELK8_CH/ELK_TX_DAT[6]\);
    
    HIEFFPLA_INST_0_57981 : NAND3A
      port map(A => HIEFFPLA_NET_0_116590, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_7[6]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_7[5]\, Y => 
        HIEFFPLA_NET_0_116585);
    
    HIEFFPLA_INST_0_42616 : AOI1A
      port map(A => HIEFFPLA_NET_0_119514, B => 
        \U50_PATTERNS/REG_ADDR[3]\, C => 
        \U50_PATTERNS/REG_ADDR[4]\, Y => HIEFFPLA_NET_0_119499);
    
    \U_ELK14_CH/U_SLAVE_1ELK/Q[4]\ : DFN1C0
      port map(D => \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/Q[4]_net_1\);
    
    HIEFFPLA_INST_0_45797 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_12[6]\, C => 
        \U50_PATTERNS/SM_BANK_SEL[7]\, Y => HIEFFPLA_NET_0_118839);
    
    HIEFFPLA_INST_0_41779 : MX2
      port map(A => HIEFFPLA_NET_0_119674, B => 
        \U50_PATTERNS/ELINK_RWA[5]\, S => 
        \U50_PATTERNS/SM_BANK_SEL_0[20]\, Y => 
        HIEFFPLA_NET_0_119696);
    
    \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[2]\ : DFN1C0
      port map(D => 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[2]_net_1\);
    
    \U_ELK14_CH/U_ELK1_SERDAT_SOURCE/SERDAT[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118461, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_6, Q => 
        \U_ELK14_CH/ELK_TX_DAT[2]\);
    
    HIEFFPLA_INST_0_45513 : AO1A
      port map(A => HIEFFPLA_NET_0_119428, B => 
        \U50_PATTERNS/ELINKS_STRT_ADDR[6]\, C => 
        HIEFFPLA_NET_0_118806, Y => HIEFFPLA_NET_0_118899);
    
    \U_MASTER_DES/U13C_MASTER_DESER/MAX_CNT[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_116947, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_16, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/MAX_CNT[7]\);
    
    \U_ELK17_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0\ : DFN1C0
      port map(D => CLK_40M_GL, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_9, Q => 
        \U_ELK17_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0_net_1\);
    
    \U50_PATTERNS/ELINK_DINA_9[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119715, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_20, Q => 
        \U50_PATTERNS/ELINK_DINA_9[4]\);
    
    HIEFFPLA_INST_0_44651 : AND2
      port map(A => \U50_PATTERNS/U4E_REGCROSS/DELCNT[0]_net_1\, 
        B => \U50_PATTERNS/U4E_REGCROSS/DELCNT[1]_net_1\, Y => 
        HIEFFPLA_NET_0_119072);
    
    \U50_PATTERNS/ELINK_ADDRA_4[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119982, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_2, Q => 
        \U50_PATTERNS/ELINK_ADDRA_4[1]\);
    
    HIEFFPLA_INST_0_49622 : MX2
      port map(A => \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[1]_net_1\, B
         => \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\, S => 
        \BIT_OS_SEL_7[2]\, Y => HIEFFPLA_NET_0_118095);
    
    \U_ELK13_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]\ : DFN1C0
      port map(D => \U_ELK13_CH/U_SLAVE_1ELK/Q[0]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]_net_1\);
    
    \U_ELK10_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]\ : DFN1C0
      port map(D => \U_ELK10_CH/U_SLAVE_1ELK/Q[6]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]_net_1\);
    
    \U50_PATTERNS/OP_MODE_T[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119603, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_17, Q => 
        \U50_PATTERNS/OP_MODE_T[6]\);
    
    HIEFFPLA_INST_0_40306 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_10[0]\, B => 
        HIEFFPLA_NET_0_119578, S => HIEFFPLA_NET_0_119239, Y => 
        HIEFFPLA_NET_0_119863);
    
    HIEFFPLA_INST_0_58175 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_11[0]\, B => 
        HIEFFPLA_NET_0_116680, S => HIEFFPLA_NET_0_117163, Y => 
        HIEFFPLA_NET_0_116554);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_2[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116754, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_5, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_2[1]\);
    
    \U50_PATTERNS/OP_MODE_T[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119602, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_17, Q => 
        \U50_PATTERNS/OP_MODE_T[7]\);
    
    AFLSDF_INV_49 : INV
      port map(A => DCB_SALT_SEL_c, Y => \AFLSDF_INV_49\);
    
    \U50_PATTERNS/ELINK_DINA_15[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119822, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_16, Q => 
        \U50_PATTERNS/ELINK_DINA_15[1]\);
    
    HIEFFPLA_INST_0_48343 : MX2
      port map(A => 
        \U_ELK17_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]_net_1\, B => 
        \U_ELK17_CH/ELK_TX_DAT[6]\, S => 
        \U_ELK17_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118334);
    
    \U50_PATTERNS/ELINK_DINA_10[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119862, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_9, Q => 
        \U50_PATTERNS/ELINK_DINA_10[1]\);
    
    HIEFFPLA_INST_0_37970 : MX2
      port map(A => \U200B_ELINKS/LOC_STOP_ADDR[6]\, B => 
        \ELKS_STOP_ADDR[6]\, S => 
        \U200B_ELINKS/GP_PG_SM_0[10]_net_1\, Y => 
        HIEFFPLA_NET_0_120181);
    
    \U_ELK19_CH/U_ELK1_SERDAT_SOURCE/SERDAT[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118236, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_15, Q => 
        \U_ELK19_CH/ELK_TX_DAT[2]\);
    
    HIEFFPLA_INST_0_53310 : AND2A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[8]_net_1\, B => 
        HIEFFPLA_NET_0_116982, Y => HIEFFPLA_NET_0_117433);
    
    \U_ELK2_CH/U_ELK1_SERDAT_SOURCE/SERDAT[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118148, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_13, Q => 
        \U_ELK2_CH/ELK_TX_DAT[0]\);
    
    HIEFFPLA_INST_0_61463 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_6[3]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_22[3]\, S
         => \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_5[4]_net_1\, 
        Y => HIEFFPLA_NET_0_116123);
    
    HIEFFPLA_INST_0_47208 : MX2
      port map(A => HIEFFPLA_NET_0_118544, B => 
        HIEFFPLA_NET_0_118541, S => \BIT_OS_SEL_4[1]\, Y => 
        HIEFFPLA_NET_0_118534);
    
    HIEFFPLA_INST_0_63080 : XA1B
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[1]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[0]\, C => 
        HIEFFPLA_NET_0_117078, Y => HIEFFPLA_NET_0_115893);
    
    HIEFFPLA_INST_0_45793 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_7[5]\, C => 
        \U50_PATTERNS/SM_BANK_SEL[12]\, Y => 
        HIEFFPLA_NET_0_118840);
    
    HIEFFPLA_INST_0_115779 : AO18
      port map(A => HIEFFPLA_NET_0_115805, B => 
        \U200A_TFC/LOC_STOP_ADDR[1]\, C => \TFC_ADDRB[1]\, Y => 
        HIEFFPLA_NET_0_115807);
    
    \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[1]\ : DFN1C0
      port map(D => 
        \U_ELK6_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\);
    
    HIEFFPLA_INST_0_46477 : AO1A
      port map(A => HIEFFPLA_NET_0_119571, B => 
        HIEFFPLA_NET_0_119556, C => 
        \U50_PATTERNS/WR_XFER_TYPE[7]_net_1\, Y => 
        HIEFFPLA_NET_0_118682);
    
    \U50_PATTERNS/ELINKS_STRT_ADDR_T[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120102, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_21, Q => 
        \U50_PATTERNS/ELINKS_STRT_ADDR_T[1]\);
    
    HIEFFPLA_INST_0_62280 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_3[1]\, 
        B => HIEFFPLA_NET_0_117114, S => HIEFFPLA_NET_0_117178, Y
         => HIEFFPLA_NET_0_116009);
    
    \U_MASTER_DES/U13C_MASTER_DESER/RECD_SER_WORD[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_116902, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_29, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/RECD_SER_WORD[2]_net_1\);
    
    \U_ELK16_CH/U_ELK1_CMD_TX/SER_OUT_RI\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118375, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_10, Q => 
        \U_ELK16_CH/U_ELK1_CMD_TX/SER_OUT_RI_net_1\);
    
    HIEFFPLA_INST_0_43901 : MX2
      port map(A => HIEFFPLA_NET_0_119578, B => 
        \U50_PATTERNS/TFC_DINA[0]\, S => HIEFFPLA_NET_0_119294, Y
         => HIEFFPLA_NET_0_119197);
    
    HIEFFPLA_INST_0_59516 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_28[2]\, B => 
        HIEFFPLA_NET_0_116687, S => HIEFFPLA_NET_0_117094, Y => 
        HIEFFPLA_NET_0_116384);
    
    HIEFFPLA_INST_0_53680 : MX2
      port map(A => HIEFFPLA_NET_0_117383, B => 
        HIEFFPLA_NET_0_117234, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[1]_net_1\, Y
         => HIEFFPLA_NET_0_117373);
    
    HIEFFPLA_INST_0_50618 : MX2
      port map(A => HIEFFPLA_NET_0_117904, B => 
        HIEFFPLA_NET_0_117902, S => \BIT_OS_SEL_4[1]\, Y => 
        HIEFFPLA_NET_0_117915);
    
    HIEFFPLA_INST_0_47622 : NAND2B
      port map(A => \OP_MODE_c_2[1]\, B => \PATT_ELK_DAT_14[3]\, 
        Y => HIEFFPLA_NET_0_118460);
    
    AFLSDF_INV_47 : INV
      port map(A => DCB_SALT_SEL_c, Y => \AFLSDF_INV_47\);
    
    HIEFFPLA_INST_0_41206 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_3[4]\, B => 
        HIEFFPLA_NET_0_119570, S => HIEFFPLA_NET_0_119247, Y => 
        HIEFFPLA_NET_0_119763);
    
    HIEFFPLA_INST_0_54626 : AO1E
      port map(A => HIEFFPLA_NET_0_116678, B => 
        HIEFFPLA_NET_0_116593, C => HIEFFPLA_NET_0_117204, Y => 
        HIEFFPLA_NET_0_117231);
    
    HIEFFPLA_INST_0_44206 : MX2
      port map(A => \U50_PATTERNS/TFC_STRT_ADDR_T[4]\, B => 
        \U50_PATTERNS/RD_USB_ADBUS[4]\, S => 
        HIEFFPLA_NET_0_119491, Y => HIEFFPLA_NET_0_119160);
    
    \U_ELK16_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]\ : DFN1C0
      port map(D => \U_ELK16_CH/U_SLAVE_1ELK/Q[10]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]_net_1\);
    
    \U50_PATTERNS/WR_USB_ADBUS[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118984, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_15, Q => 
        \U50_PATTERNS/WR_USB_ADBUS[1]\);
    
    \U200A_TFC/RX_SER_WORD_2DEL[4]\ : DFN1C0
      port map(D => \U200A_TFC/RX_SER_WORD_1DEL[4]_net_1\, CLK
         => CLK_40M_GL, CLR => P_MASTER_POR_B_c, Q => 
        \U200A_TFC/RX_SER_WORD_2DEL[4]_net_1\);
    
    HIEFFPLA_INST_0_59118 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_24[1]\, B => 
        HIEFFPLA_NET_0_116429, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_2[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116433);
    
    \U_ELK11_CH/U_SLAVE_1ELK/RECD_SER_WORD[4]\ : DFN1C0
      port map(D => \U_ELK11_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[4]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_11[4]\);
    
    HIEFFPLA_INST_0_56534 : AND3A
      port map(A => HIEFFPLA_NET_0_117430, B => \BIT_OS_SEL_1[2]\, 
        C => \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[10]_net_1\, 
        Y => HIEFFPLA_NET_0_116844);
    
    \U_EXEC_MASTER/SYNC_BRD_RST_BI_1\ : DFI1P0
      port map(D => \U_EXEC_MASTER/DEV_RST_1B_i\, CLK => 
        CCC_160M_FXD, PRE => DEV_RST_B_c, QN => 
        \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_1\);
    
    \U50_PATTERNS/U4D_REGCROSS/SAMP_ONE[6]\ : DFN1C0
      port map(D => \U50_PATTERNS/ELINKS_STOP_ADDR[6]\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_25, Q => 
        \U50_PATTERNS/U4D_REGCROSS/SAMP_ONE[6]_net_1\);
    
    HIEFFPLA_INST_0_38081 : NAND3C
      port map(A => \U200B_ELINKS/RX_SER_WORD_3DEL_i_0[1]\, B => 
        \U200B_ELINKS/RX_SER_WORD_3DEL[0]_net_1\, C => 
        HIEFFPLA_NET_0_120156, Y => HIEFFPLA_NET_0_120157);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_13[4]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116246, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_1, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_13[4]\);
    
    \U50_PATTERNS/ELINK_ADDRA_19[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120010, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_13, Q => 
        \U50_PATTERNS/ELINK_ADDRA_19[5]\);
    
    \U_ELK19_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]\ : DFN1C0
      port map(D => \U_ELK19_CH/U_SLAVE_1ELK/Q[1]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]_net_1\);
    
    \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[3]\ : DFN1C0
      port map(D => \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\);
    
    \U50_PATTERNS/U4E_REGCROSS/LOCAL_REG_VAL_3[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119059, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_1, Q => \OP_MODE_c_3[1]\);
    
    HIEFFPLA_INST_0_42382 : AO1A
      port map(A => HIEFFPLA_NET_0_119019, B => 
        \U50_PATTERNS/RD_USB_ADBUS[0]\, C => 
        HIEFFPLA_NET_0_119541, Y => HIEFFPLA_NET_0_119549);
    
    \U_ELK8_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0\ : DFN1C0
      port map(D => CLK_40M_GL, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_12, Q => 
        \U_ELK8_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0_net_1\);
    
    \ALL_PLL_LOCK_pad/U0/U1\ : IOTRI_OB_EB
      port map(D => ALL_PLL_LOCK_c, E => \VCC\, DOUT => 
        \ALL_PLL_LOCK_pad/U0/NET1\, EOUT => 
        \ALL_PLL_LOCK_pad/U0/NET2\);
    
    \U_ELK5_CH/U_ELK1_CMD_TX/SER_OUT_FI\ : DFN1C0
      port map(D => 
        \U_ELK5_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_14, Q
         => \U_ELK5_CH/U_ELK1_CMD_TX/SER_OUT_FI_net_1\);
    
    \U_ELK17_CH/U_SLAVE_1ELK/Q[6]\ : DFN1C0
      port map(D => \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/Q[6]_net_1\);
    
    HIEFFPLA_INST_0_53672 : MX2
      port map(A => HIEFFPLA_NET_0_116121, B => 
        HIEFFPLA_NET_0_116024, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[3]_net_1\, Y
         => HIEFFPLA_NET_0_117374);
    
    HIEFFPLA_INST_0_41395 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_6[1]\, B => 
        HIEFFPLA_NET_0_119576, S => HIEFFPLA_NET_0_119258, Y => 
        HIEFFPLA_NET_0_119742);
    
    HIEFFPLA_INST_0_51290 : MX2
      port map(A => HIEFFPLA_NET_0_117799, B => 
        HIEFFPLA_NET_0_117819, S => \BIT_OS_SEL_2[1]\, Y => 
        HIEFFPLA_NET_0_117801);
    
    HIEFFPLA_INST_0_46993 : MX2
      port map(A => HIEFFPLA_NET_0_118566, B => 
        HIEFFPLA_NET_0_118586, S => \BIT_OS_SEL[0]\, Y => 
        \U_ELK11_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[0]\);
    
    HIEFFPLA_INST_0_57131 : XA1B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_2[0]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_2[1]\, C => 
        HIEFFPLA_NET_0_117179, Y => HIEFFPLA_NET_0_116734);
    
    HIEFFPLA_INST_0_54442 : MX2
      port map(A => HIEFFPLA_NET_0_116182, B => 
        HIEFFPLA_NET_0_116071, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[3]_net_1\, Y => 
        HIEFFPLA_NET_0_117265);
    
    HIEFFPLA_INST_0_54325 : MX2
      port map(A => HIEFFPLA_NET_0_116147, B => 
        HIEFFPLA_NET_0_116048, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_2[3]_net_1\, Y
         => HIEFFPLA_NET_0_117280);
    
    HIEFFPLA_INST_0_52782 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_11[0]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_12[0]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_1[0]\, Y => 
        HIEFFPLA_NET_0_117512);
    
    HIEFFPLA_INST_0_47477 : MX2
      port map(A => HIEFFPLA_NET_0_118499, B => 
        HIEFFPLA_NET_0_118496, S => \BIT_OS_SEL_3[1]\, Y => 
        HIEFFPLA_NET_0_118486);
    
    \U_ELK1_CH/U_ELK1_CMD_TX/SER_OUT_FI\ : DFI1C0
      port map(D => 
        \U_ELK1_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_14, QN
         => \U_ELK1_CH/U_ELK1_CMD_TX/SER_OUT_FI_i\);
    
    HIEFFPLA_INST_0_37797 : AND3
      port map(A => HIEFFPLA_NET_0_120223, B => 
        HIEFFPLA_NET_0_120233, C => HIEFFPLA_NET_0_120198, Y => 
        HIEFFPLA_NET_0_120205);
    
    HIEFFPLA_INST_0_47624 : AND2A
      port map(A => \OP_MODE_c_2[1]\, B => \PATT_ELK_DAT_14[5]\, 
        Y => HIEFFPLA_NET_0_118458);
    
    HIEFFPLA_INST_0_53460 : MX2
      port map(A => HIEFFPLA_NET_0_116220, B => 
        HIEFFPLA_NET_0_116113, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[3]_net_1\, Y
         => HIEFFPLA_NET_0_117405);
    
    HIEFFPLA_INST_0_45420 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_14[0]\, C => 
        \U50_PATTERNS/SM_BANK_SEL[5]\, Y => HIEFFPLA_NET_0_118916);
    
    \U_ELK14_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118465, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_2, Q => 
        \U_ELK14_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]_net_1\);
    
    HIEFFPLA_INST_0_42301 : AND2A
      port map(A => HIEFFPLA_NET_0_119275, B => 
        \U50_PATTERNS/RD_USB_ADBUS[0]\, Y => 
        HIEFFPLA_NET_0_119578);
    
    HIEFFPLA_INST_0_41422 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_6[4]\, B => 
        HIEFFPLA_NET_0_119570, S => HIEFFPLA_NET_0_119258, Y => 
        HIEFFPLA_NET_0_119739);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_10[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116562, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_6, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_10[0]\);
    
    \U_ELK15_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118424, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_9, Q => 
        \U_ELK15_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]_net_1\);
    
    HIEFFPLA_INST_0_60268 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_8[0]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_24[0]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_1[4]_net_1\, Y
         => HIEFFPLA_NET_0_116289);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_30[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116354, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_18, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_30[2]\);
    
    HIEFFPLA_INST_0_58207 : MX2
      port map(A => HIEFFPLA_NET_0_116687, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_11[2]\, S => 
        HIEFFPLA_NET_0_117329, Y => HIEFFPLA_NET_0_116550);
    
    HIEFFPLA_INST_0_54610 : MX2
      port map(A => HIEFFPLA_NET_0_117287, B => 
        HIEFFPLA_NET_0_117280, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[2]_net_1\, Y => 
        HIEFFPLA_NET_0_117233);
    
    \U_ELK17_CH/U_SLAVE_1ELK/Q[11]\ : DFN1C0
      port map(D => \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/Q[11]_net_1\);
    
    \U_ELK13_CH/U_ELK1_SERDAT_SOURCE/SERDAT[7]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118501, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_4, Q => 
        \U_ELK13_CH/ELK_TX_DAT[7]\);
    
    HIEFFPLA_INST_0_41873 : AOI1B
      port map(A => HIEFFPLA_NET_0_119389, B => 
        \U50_PATTERNS/SM_BANK_SEL[17]\, C => 
        HIEFFPLA_NET_0_119647, Y => HIEFFPLA_NET_0_119678);
    
    \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[7]\ : DFN1C0
      port map(D => \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\);
    
    \U_EXEC_MASTER/DEL_CNT[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117789, CLK => CLK_40M_GL, CLR
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i\, Q => 
        \U_EXEC_MASTER/DEL_CNT[6]\);
    
    HIEFFPLA_INST_0_57949 : NAND2B
      port map(A => HIEFFPLA_NET_0_116649, B => 
        HIEFFPLA_NET_0_116589, Y => HIEFFPLA_NET_0_116594);
    
    HIEFFPLA_INST_0_48270 : MX2
      port map(A => HIEFFPLA_NET_0_118361, B => 
        HIEFFPLA_NET_0_118359, S => \BIT_OS_SEL_3[0]\, Y => 
        \U_ELK16_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[4]\);
    
    \U200A_TFC/ADDR_POINTER[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120368, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_30, Q => \TFC_ADDRB[0]\);
    
    HIEFFPLA_INST_0_45236 : NAND3C
      port map(A => HIEFFPLA_NET_0_118736, B => 
        HIEFFPLA_NET_0_118747, C => HIEFFPLA_NET_0_118756, Y => 
        HIEFFPLA_NET_0_118960);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_27[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116393, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_2, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_27[1]\);
    
    \U_ELK2_CH/U_SLAVE_1ELK/Q[11]\ : DFN1C0
      port map(D => \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/Q[11]_net_1\);
    
    HIEFFPLA_INST_0_44328 : XO1
      port map(A => \TFC_STRT_ADDR[4]\, B => 
        \U50_PATTERNS/U4A_REGCROSS/SAMP_TWO[4]_net_1\, C => 
        HIEFFPLA_NET_0_119138, Y => HIEFFPLA_NET_0_119141);
    
    \U_DDR_TFC/BIBUF_LVDS_0/U0/U1\ : IOBI_ID_OD_EB
      port map(DR => TFC_OUT_R, DF => TFC_OUT_F, CLR => \GND\, E
         => DCB_SALT_SEL_c, ICLK => CCC_160M_ADJ, OCLK => 
        CCC_160M_FXD, YIN => \U_DDR_TFC/BIBUF_LVDS_0/U0/NET4\, 
        DOUT => \U_DDR_TFC/BIBUF_LVDS_0/U0/NET1\, EOUT => 
        \U_DDR_TFC/BIBUF_LVDS_0/U0/NET2\, YR => TFC_IN_DDR_R, YF
         => TFC_IN_DDR_F);
    
    \U50_PATTERNS/ELINK_DINA_15[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119816, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_17, Q => 
        \U50_PATTERNS/ELINK_DINA_15[7]\);
    
    \U_ELK11_CH/U_ELK1_SERDAT_SOURCE/SERDAT[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118598, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_0, Q => 
        \U_ELK11_CH/ELK_TX_DAT[0]\);
    
    HIEFFPLA_INST_0_60435 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_9[4]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_10[4]\, S
         => \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_1[0]\, Y
         => HIEFFPLA_NET_0_116266);
    
    \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[11]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117719, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_33, Q => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[11]_net_1\);
    
    HIEFFPLA_INST_0_51130 : MX2
      port map(A => HIEFFPLA_NET_0_117812, B => 
        HIEFFPLA_NET_0_117810, S => \BIT_OS_SEL_3[1]\, Y => 
        HIEFFPLA_NET_0_117823);
    
    HIEFFPLA_INST_0_49358 : MX2
      port map(A => 
        \U_ELK2_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]_net_1\, B => 
        \U_ELK2_CH/ELK_TX_DAT[7]\, S => 
        \U_ELK2_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118150);
    
    HIEFFPLA_INST_0_61400 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_21[4]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_22[4]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_3[0]\, Y => 
        HIEFFPLA_NET_0_116131);
    
    HIEFFPLA_INST_0_55770 : MX2
      port map(A => HIEFFPLA_NET_0_117017, B => 
        HIEFFPLA_NET_0_116040, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[2]\, Y => 
        HIEFFPLA_NET_0_116992);
    
    \U0_200M_BUF/_INBUF_LVDS[0]_/U0/U1\ : IOIN_IB
      port map(YIN => \U0_200M_BUF/\\\\INBUF_LVDS[0]\\\\/U0/NET1\, 
        Y => Y);
    
    HIEFFPLA_INST_0_60579 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_13[2]\, B => 
        HIEFFPLA_NET_0_117181, S => HIEFFPLA_NET_0_117137, Y => 
        HIEFFPLA_NET_0_116248);
    
    HIEFFPLA_INST_0_57027 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_2[2]\, B => 
        HIEFFPLA_NET_0_116733, S => HIEFFPLA_NET_0_117601, Y => 
        HIEFFPLA_NET_0_116753);
    
    HIEFFPLA_INST_0_56310 : AO1
      port map(A => HIEFFPLA_NET_0_117429, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[1]_net_1\, C => 
        HIEFFPLA_NET_0_116872, Y => HIEFFPLA_NET_0_116896);
    
    \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[9]\ : DFN1C0
      port map(D => \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\);
    
    HIEFFPLA_INST_0_53519 : NAND3A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[4]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[2]_net_1\, C => 
        HIEFFPLA_NET_0_117318, Y => HIEFFPLA_NET_0_117396);
    
    HIEFFPLA_INST_0_43056 : AOI1D
      port map(A => HIEFFPLA_NET_0_119434, B => 
        HIEFFPLA_NET_0_119365, C => HIEFFPLA_NET_0_119014, Y => 
        HIEFFPLA_NET_0_119390);
    
    \U50_PATTERNS/U4C_REGCROSS/SAMP_TWO[7]\ : DFN1C0
      port map(D => \U50_PATTERNS/U4C_REGCROSS/SAMP_ONE[7]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_22_0, Q => 
        \U50_PATTERNS/U4C_REGCROSS/SAMP_TWO[7]_net_1\);
    
    HIEFFPLA_INST_0_46058 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_14[5]\, C => 
        \U50_PATTERNS/SM_BANK_SEL[5]\, Y => HIEFFPLA_NET_0_118776);
    
    HIEFFPLA_INST_0_43651 : AND2A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/SM_BANK_SEL[13]\, Y => 
        HIEFFPLA_NET_0_119254);
    
    HIEFFPLA_INST_0_49601 : MX2
      port map(A => 
        \U_ELK3_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]_net_1\, B => 
        \U_ELK3_CH/ELK_TX_DAT[5]\, S => 
        \U_ELK3_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118106);
    
    HIEFFPLA_INST_0_46333 : NAND3C
      port map(A => HIEFFPLA_NET_0_118859, B => 
        HIEFFPLA_NET_0_118864, C => HIEFFPLA_NET_0_118870, Y => 
        HIEFFPLA_NET_0_118714);
    
    HIEFFPLA_INST_0_48714 : MX2
      port map(A => \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\, 
        B => \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[13]_net_1\, S => 
        \BIT_OS_SEL_0[2]\, Y => HIEFFPLA_NET_0_118262);
    
    HIEFFPLA_INST_0_51437 : XA1A
      port map(A => HIEFFPLA_NET_0_117782, B => 
        \U_EXEC_MASTER/DEL_CNT[4]\, C => 
        \U_EXEC_MASTER/CCC_1_LOCK_STAT_1D_net_1\, Y => 
        HIEFFPLA_NET_0_117774);
    
    HIEFFPLA_INST_0_49615 : AND2A
      port map(A => \OP_MODE_c_5[1]\, B => \PATT_ELK_DAT_3[4]\, Y
         => HIEFFPLA_NET_0_118099);
    
    \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[1]\ : DFN1C0
      port map(D => 
        \U_ELK8_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\);
    
    \U_ELK1_CH/U_SLAVE_1ELK/RECD_SER_WORD[3]\ : DFN1C0
      port map(D => \U_ELK1_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[3]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_1[3]\);
    
    \U50_PATTERNS/ELINK_DINA_17[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119804, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_19, Q => 
        \U50_PATTERNS/ELINK_DINA_17[3]\);
    
    \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[5]\ : DFN1C0
      port map(D => \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\);
    
    \U_MASTER_DES/U13A_ADJ_160M/SDIN/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117670, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_6, Q => \U_MASTER_DES/AUX_SDIN\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_SEL_6[2]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_BIT_OS_VAL[2]\, CLK
         => CLK_40M_GL, CLR => P_MASTER_POR_B_c_27_0, Q => 
        \BIT_OS_SEL_6[2]\);
    
    \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[14]\ : DFN1C0
      port map(D => 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]_net_1\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[14]_net_1\);
    
    HIEFFPLA_INST_0_37818 : AOI1B
      port map(A => HIEFFPLA_NET_0_120158, B => 
        HIEFFPLA_NET_0_120160, C => 
        \U200B_ELINKS/GP_PG_SM[7]_net_1\, Y => 
        HIEFFPLA_NET_0_120200);
    
    \U_ELK2_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]\ : DFN1C0
      port map(D => \U_ELK2_CH/U_SLAVE_1ELK/Q[12]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]_net_1\);
    
    HIEFFPLA_INST_0_59257 : AO1C
      port map(A => HIEFFPLA_NET_0_117394, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_25[2]\, C => 
        HIEFFPLA_NET_0_117366, Y => HIEFFPLA_NET_0_116414);
    
    HIEFFPLA_INST_0_52283 : AND3A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[0]_net_1\, B => 
        HIEFFPLA_NET_0_117593, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[3]_net_1\, Y => 
        HIEFFPLA_NET_0_117591);
    
    HIEFFPLA_INST_0_43025 : OR3A
      port map(A => \U50_PATTERNS/REG_STATE[4]_net_1\, B => 
        HIEFFPLA_NET_0_119415, C => HIEFFPLA_NET_0_119398, Y => 
        HIEFFPLA_NET_0_119399);
    
    \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117721, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_31, Q => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[0]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_31[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116341, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_20, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_31[2]\);
    
    \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[1]\ : DFN1C0
      port map(D => 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[1]_net_1\);
    
    HIEFFPLA_INST_0_55949 : MX2
      port map(A => HIEFFPLA_NET_0_117014, B => 
        HIEFFPLA_NET_0_116038, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[2]\, Y => 
        HIEFFPLA_NET_0_116969);
    
    \U_EXEC_MASTER/MPOR_B_17_0\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117787, CLK => CLK_40M_GL, CLR
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_0\, Q => 
        P_MASTER_POR_B_c_17_0);
    
    \U_ELK5_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]\ : DFN1C0
      port map(D => \U_ELK5_CH/U_SLAVE_1ELK/Q[6]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]_net_1\);
    
    \U50_PATTERNS/ELINK_DINA_14[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119824, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_16, Q => 
        \U50_PATTERNS/ELINK_DINA_14[7]\);
    
    \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[2]\ : DFN1C0
      port map(D => 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[2]_net_1\);
    
    \U_ELK4_CH/U_SLAVE_1ELK/Q[2]\ : DFN1C0
      port map(D => \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/Q[2]_net_1\);
    
    HIEFFPLA_INST_0_51274 : MX2
      port map(A => HIEFFPLA_NET_0_117823, B => 
        HIEFFPLA_NET_0_117820, S => \BIT_OS_SEL_4[0]\, Y => 
        \U_ELK9_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[6]\);
    
    HIEFFPLA_INST_0_47596 : MX2
      port map(A => 
        \U_ELK14_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]_net_1\, B => 
        \U_ELK14_CH/ELK_TX_DAT[6]\, S => 
        \U_ELK14_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118469);
    
    HIEFFPLA_INST_0_42521 : OA1A
      port map(A => HIEFFPLA_NET_0_119433, B => 
        HIEFFPLA_NET_0_119010, C => \U50_PATTERNS/REG_ADDR[1]\, Y
         => HIEFFPLA_NET_0_119523);
    
    HIEFFPLA_INST_0_52274 : AND2A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[2]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[7]_net_1\, Y => 
        HIEFFPLA_NET_0_117594);
    
    \U_MASTER_DES/U13C_MASTER_DESER/BEST_BIT_OS_VAL[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_117577, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_14, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_BIT_OS_VAL[3]\);
    
    \U50_PATTERNS/TFC_DINA[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119192, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_4, Q => \U50_PATTERNS/TFC_DINA[5]\);
    
    HIEFFPLA_INST_0_58586 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_17[0]\, B => 
        HIEFFPLA_NET_0_116680, S => HIEFFPLA_NET_0_117161, Y => 
        HIEFFPLA_NET_0_116501);
    
    HIEFFPLA_INST_0_46654 : MX2
      port map(A => HIEFFPLA_NET_0_118623, B => 
        HIEFFPLA_NET_0_118620, S => \BIT_OS_SEL_5[1]\, Y => 
        HIEFFPLA_NET_0_118632);
    
    HIEFFPLA_INST_0_42866 : AO1D
      port map(A => HIEFFPLA_NET_0_119380, B => 
        HIEFFPLA_NET_0_119432, C => HIEFFPLA_NET_0_119447, Y => 
        HIEFFPLA_NET_0_119443);
    
    \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[5]\ : DFN1C0
      port map(D => 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\);
    
    HIEFFPLA_INST_0_63015 : NAND3
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[5]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[6]\, C => 
        HIEFFPLA_NET_0_115908, Y => HIEFFPLA_NET_0_115914);
    
    \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[7]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117701, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_31, Q => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[7]_net_1\);
    
    HIEFFPLA_INST_0_46076 : AND3A
      port map(A => HIEFFPLA_NET_0_119376, B => 
        \U50_PATTERNS/TFC_STRT_ADDR[2]\, C => 
        HIEFFPLA_NET_0_119431, Y => HIEFFPLA_NET_0_118772);
    
    HIEFFPLA_INST_0_45824 : NAND2A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_14[6]\, Y => 
        HIEFFPLA_NET_0_118831);
    
    HIEFFPLA_INST_0_58025 : XA1C
      port map(A => HIEFFPLA_NET_0_116573, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_7[8]\, C => 
        HIEFFPLA_NET_0_117179, Y => HIEFFPLA_NET_0_116576);
    
    HIEFFPLA_INST_0_47298 : MX2
      port map(A => HIEFFPLA_NET_0_118532, B => 
        HIEFFPLA_NET_0_118520, S => \BIT_OS_SEL_5[0]\, Y => 
        \U_ELK12_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[7]\);
    
    HIEFFPLA_INST_0_41377 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_5[7]\, B => 
        HIEFFPLA_NET_0_119560, S => HIEFFPLA_NET_0_119251, Y => 
        HIEFFPLA_NET_0_119744);
    
    \U_ELK6_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL\ : DFN1C0
      port map(D => 
        \U_ELK6_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL_net_1\);
    
    HIEFFPLA_INST_0_53787 : MX2
      port map(A => HIEFFPLA_NET_0_117265, B => 
        HIEFFPLA_NET_0_117316, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[2]_net_1\, Y
         => HIEFFPLA_NET_0_117352);
    
    \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[9]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[7]_net_1\, CLK => 
        CCC_160M_ADJ, CLR => P_MASTER_POR_B_c_34_0, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[9]_net_1\);
    
    \U_ELK4_CH/U_ELK1_CMD_TX/START_RISE\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118059, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_13, Q => 
        \U_ELK4_CH/U_ELK1_CMD_TX/START_RISE_net_1\);
    
    \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[8]\ : DFN1C0
      port map(D => 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\);
    
    HIEFFPLA_INST_0_45544 : NOR2A
      port map(A => \U50_PATTERNS/ELINKS_STRT_ADDR[4]\, B => 
        HIEFFPLA_NET_0_119428, Y => HIEFFPLA_NET_0_118893);
    
    HIEFFPLA_INST_0_42377 : NAND3B
      port map(A => \U50_PATTERNS/RD_XFER_TYPE[6]_net_1\, B => 
        \U50_PATTERNS/RD_XFER_TYPE[3]_net_1\, C => 
        HIEFFPLA_NET_0_119550, Y => HIEFFPLA_NET_0_119551);
    
    HIEFFPLA_INST_0_50136 : MX2
      port map(A => \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[1]_net_1\, B
         => \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\, S => 
        \BIT_OS_SEL_6[2]\, Y => HIEFFPLA_NET_0_118003);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_28[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116383, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_2, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_28[3]\);
    
    AFLSDF_INV_23 : INV
      port map(A => DCB_SALT_SEL_c, Y => \AFLSDF_INV_23\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_115939, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_24_0, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[2]_net_1\);
    
    HIEFFPLA_INST_0_63028 : AND2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[11]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[13]\, Y => 
        HIEFFPLA_NET_0_115909);
    
    HIEFFPLA_INST_0_55122 : AO1C
      port map(A => HIEFFPLA_NET_0_117107, B => 
        HIEFFPLA_NET_0_117394, C => HIEFFPLA_NET_0_117086, Y => 
        HIEFFPLA_NET_0_117117);
    
    HIEFFPLA_INST_0_41937 : AND3C
      port map(A => HIEFFPLA_NET_0_119253, B => 
        HIEFFPLA_NET_0_119262, C => \U50_PATTERNS/SM_BANK_SEL[9]\, 
        Y => HIEFFPLA_NET_0_119654);
    
    \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[11]\ : DFN1C0
      port map(D => \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\);
    
    \U_ELK12_CH/U_ELK1_SERDAT_SOURCE/SERDAT[7]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118546, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_2, Q => 
        \U_ELK12_CH/ELK_TX_DAT[7]\);
    
    HIEFFPLA_INST_0_63151 : AND2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[3]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[2]_net_1\, Y => 
        HIEFFPLA_NET_0_115875);
    
    \U_ELK9_CH/U_SLAVE_1ELK/Q[12]\ : DFN1C0
      port map(D => \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/Q[12]_net_1\);
    
    \U_ELK3_CH/U_SLAVE_1ELK/Q[3]\ : DFN1C0
      port map(D => \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/Q[3]_net_1\);
    
    HIEFFPLA_INST_0_51433 : XA1A
      port map(A => HIEFFPLA_NET_0_117778, B => 
        \U_EXEC_MASTER/DEL_CNT[3]\, C => 
        \U_EXEC_MASTER/CCC_1_LOCK_STAT_1D_net_1\, Y => 
        HIEFFPLA_NET_0_117775);
    
    HIEFFPLA_INST_0_41751 : MX2
      port map(A => HIEFFPLA_NET_0_119679, B => 
        \U50_PATTERNS/ELINK_RWA[1]\, S => 
        \U50_PATTERNS/SM_BANK_SEL_0[20]\, Y => 
        HIEFFPLA_NET_0_119700);
    
    \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[10]\ : DFN1C0
      port map(D => 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\);
    
    \U50_PATTERNS/U4D_REGCROSS/SAMP_ONE[3]\ : DFN1C0
      port map(D => \U50_PATTERNS/ELINKS_STOP_ADDR[3]\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_25, Q => 
        \U50_PATTERNS/U4D_REGCROSS/SAMP_ONE[3]_net_1\);
    
    HIEFFPLA_INST_0_38088 : NAND2B
      port map(A => \U200B_ELINKS/RX_SER_WORD_3DEL_i_0[7]\, B => 
        \U200B_ELINKS/RX_SER_WORD_3DEL[6]_net_1\, Y => 
        HIEFFPLA_NET_0_120155);
    
    HIEFFPLA_INST_0_43853 : MX2
      port map(A => HIEFFPLA_NET_0_119519, B => 
        \U50_PATTERNS/TFC_ADDRA[4]\, S => HIEFFPLA_NET_0_119294, 
        Y => HIEFFPLA_NET_0_119203);
    
    \U50_PATTERNS/ELINK_DINA_7[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119735, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_17, Q => 
        \U50_PATTERNS/ELINK_DINA_7[0]\);
    
    HIEFFPLA_INST_0_58530 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_16[3]\, B => 
        HIEFFPLA_NET_0_116505, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_1[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116509);
    
    HIEFFPLA_INST_0_57943 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_7[8]\, B => 
        HIEFFPLA_NET_0_116576, S => HIEFFPLA_NET_0_117113, Y => 
        HIEFFPLA_NET_0_116595);
    
    \U_ELK3_CH/U_SLAVE_1ELK/Q[8]\ : DFN1C0
      port map(D => \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/Q[8]_net_1\);
    
    \U_ELK16_CH/U_SLAVE_1ELK/RECD_SER_WORD[2]\ : DFN1C0
      port map(D => \U_ELK16_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[2]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_16[2]\);
    
    HIEFFPLA_INST_0_54854 : AND3A
      port map(A => HIEFFPLA_NET_0_117369, B => 
        HIEFFPLA_NET_0_117361, C => HIEFFPLA_NET_0_117179, Y => 
        HIEFFPLA_NET_0_117189);
    
    HIEFFPLA_INST_0_44441 : XOR2
      port map(A => \TFC_STOP_ADDR[7]\, B => 
        \U50_PATTERNS/U4B_REGCROSS/SAMP_TWO[7]_net_1\, Y => 
        HIEFFPLA_NET_0_119116);
    
    HIEFFPLA_INST_0_56519 : AND3A
      port map(A => HIEFFPLA_NET_0_117430, B => \BIT_OS_SEL_1[2]\, 
        C => \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[7]_net_1\, 
        Y => HIEFFPLA_NET_0_116847);
    
    HIEFFPLA_INST_0_46537 : AND2
      port map(A => \ELK0_TX_DAT[0]\, B => 
        \U_ELK0_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118669);
    
    HIEFFPLA_INST_0_45835 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_14[2]\, C => 
        \U50_PATTERNS/SM_BANK_SEL[5]\, Y => HIEFFPLA_NET_0_118829);
    
    \U50_PATTERNS/ELINK_ADDRA_7[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119953, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_6, Q => 
        \U50_PATTERNS/ELINK_ADDRA_7[6]\);
    
    HIEFFPLA_INST_0_41152 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_2[6]\, B => 
        HIEFFPLA_NET_0_119566, S => HIEFFPLA_NET_0_119278, Y => 
        HIEFFPLA_NET_0_119769);
    
    HIEFFPLA_INST_0_51458 : NAND2
      port map(A => DCB_SALT_SEL_c, B => HIEFFPLA_NET_0_117787, Y
         => HIEFFPLA_NET_0_117769);
    
    HIEFFPLA_INST_0_45073 : AO1D
      port map(A => \U50_PATTERNS/REG_STATE[1]_net_1\, B => 
        HIEFFPLA_NET_0_119432, C => HIEFFPLA_NET_0_118986, Y => 
        HIEFFPLA_NET_0_118987);
    
    HIEFFPLA_INST_0_43973 : MX2
      port map(A => HIEFFPLA_NET_0_119275, B => 
        \U50_PATTERNS/TFC_RWA\, S => HIEFFPLA_NET_0_119294, Y => 
        HIEFFPLA_NET_0_119189);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_6[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116629, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_12, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_6[3]\);
    
    HIEFFPLA_INST_0_62511 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_7[0]\, 
        B => HIEFFPLA_NET_0_117096, S => HIEFFPLA_NET_0_117174, Y
         => HIEFFPLA_NET_0_115980);
    
    HIEFFPLA_INST_0_50190 : MX2
      port map(A => \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\, B
         => \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\, S => 
        \BIT_OS_SEL_6[2]\, Y => HIEFFPLA_NET_0_117995);
    
    HIEFFPLA_INST_0_43570 : NAND2B
      port map(A => \U50_PATTERNS/SM_BANK_SEL[12]\, B => 
        \U50_PATTERNS/SM_BANK_SEL[13]\, Y => 
        HIEFFPLA_NET_0_119286);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_1[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116169, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_8, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_1[1]\);
    
    HIEFFPLA_INST_0_43733 : AND3B
      port map(A => HIEFFPLA_NET_0_119580, B => 
        HIEFFPLA_NET_0_119590, C => 
        \U50_PATTERNS/RD_USB_ADBUS[4]\, Y => 
        HIEFFPLA_NET_0_119228);
    
    HIEFFPLA_INST_0_45992 : NAND3C
      port map(A => HIEFFPLA_NET_0_118938, B => 
        HIEFFPLA_NET_0_118830, C => HIEFFPLA_NET_0_118951, Y => 
        HIEFFPLA_NET_0_118795);
    
    HIEFFPLA_INST_0_43639 : NAND2B
      port map(A => \U50_PATTERNS/SM_BANK_SEL_0[21]\, B => 
        \U50_PATTERNS/SM_BANK_SEL[13]\, Y => 
        HIEFFPLA_NET_0_119258);
    
    HIEFFPLA_INST_0_41107 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_2[1]\, B => 
        HIEFFPLA_NET_0_119576, S => HIEFFPLA_NET_0_119278, Y => 
        HIEFFPLA_NET_0_119774);
    
    HIEFFPLA_INST_0_60054 : MX2
      port map(A => HIEFFPLA_NET_0_116687, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_5[2]\, S => 
        HIEFFPLA_NET_0_117218, Y => HIEFFPLA_NET_0_116316);
    
    HIEFFPLA_INST_0_54949 : AND3
      port map(A => HIEFFPLA_NET_0_117244, B => 
        HIEFFPLA_NET_0_117240, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_3[6]_net_1\, Y => 
        HIEFFPLA_NET_0_117161);
    
    \U_EXEC_MASTER/DEL_CNT[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117792, CLK => CLK_40M_GL, CLR
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i\, Q => 
        \U_EXEC_MASTER/DEL_CNT[3]\);
    
    AFLSDF_INV_14 : INV
      port map(A => DCB_SALT_SEL_c, Y => \AFLSDF_INV_14\);
    
    HIEFFPLA_INST_0_44916 : NAND2B
      port map(A => HIEFFPLA_NET_0_119019, B => 
        \U50_PATTERNS/USB_RXF_B\, Y => HIEFFPLA_NET_0_119020);
    
    HIEFFPLA_INST_0_111645 : AO18
      port map(A => HIEFFPLA_NET_0_115950, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_SEQCNT[1]\, C => 
        HIEFFPLA_NET_0_116976, Y => HIEFFPLA_NET_0_115836);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_21[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116145, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_3, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_21[0]\);
    
    \U50_PATTERNS/ELINK_RWA[7]/U1\ : DFN1P0
      port map(D => HIEFFPLA_NET_0_119694, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_6, Q => \U50_PATTERNS/ELINK_RWA[7]\);
    
    HIEFFPLA_INST_0_56467 : AOI1D
      port map(A => HIEFFPLA_NET_0_117432, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_SEL[3]_net_1\, C
         => \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[7]_net_1\, Y
         => HIEFFPLA_NET_0_116857);
    
    HIEFFPLA_INST_0_59653 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_2[1]\, B => 
        HIEFFPLA_NET_0_116677, S => HIEFFPLA_NET_0_117090, Y => 
        HIEFFPLA_NET_0_116366);
    
    HIEFFPLA_INST_0_49866 : AND2A
      port map(A => \OP_MODE_c_1[1]\, B => \PATT_ELK_DAT_4[6]\, Y
         => HIEFFPLA_NET_0_118052);
    
    \U_ELK9_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]\ : DFN1C0
      port map(D => \U_ELK9_CH/U_SLAVE_1ELK/Q[2]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]_net_1\);
    
    HIEFFPLA_INST_0_44808 : AOI1A
      port map(A => \U50_PATTERNS/USB_RXF_B\, B => 
        HIEFFPLA_NET_0_119452, C => HIEFFPLA_NET_0_119042, Y => 
        HIEFFPLA_NET_0_119044);
    
    \U200B_ELINKS/RX_SER_WORD_1DEL[5]\ : DFN1C0
      port map(D => \ELK_RX_SER_WORD_0[5]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_23, Q => 
        \U200B_ELINKS/RX_SER_WORD_1DEL[5]_net_1\);
    
    HIEFFPLA_INST_0_54937 : AND2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_3[6]_net_1\, B => 
        HIEFFPLA_NET_0_117341, Y => HIEFFPLA_NET_0_117165);
    
    \U_MASTER_DES/U13C_MASTER_DESER/Q[11]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[11]_net_1\, CLK => 
        CCC_160M_FXD, CLR => P_MASTER_POR_B_c_23, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/Q[11]_net_1\);
    
    \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[0]\ : DFN1C0
      port map(D => 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[0]_net_1\);
    
    \U_ELK19_CH/U_SLAVE_1ELK/Q[9]\ : DFN1C0
      port map(D => \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/Q[9]_net_1\);
    
    HIEFFPLA_INST_0_61637 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_8[1]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_24[1]\, S
         => \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_4[4]_net_1\, 
        Y => HIEFFPLA_NET_0_116099);
    
    \U_ELK4_CH/U_SLAVE_1ELK/Q[12]\ : DFN1C0
      port map(D => \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/Q[12]_net_1\);
    
    HIEFFPLA_INST_0_46135 : AO1
      port map(A => HIEFFPLA_NET_0_119277, B => 
        \U50_PATTERNS/ELINK_DOUTA_11[4]\, C => 
        HIEFFPLA_NET_0_118933, Y => HIEFFPLA_NET_0_118758);
    
    HIEFFPLA_INST_0_45200 : NAND3C
      port map(A => HIEFFPLA_NET_0_118745, B => 
        HIEFFPLA_NET_0_118754, C => HIEFFPLA_NET_0_118762, Y => 
        HIEFFPLA_NET_0_118966);
    
    HIEFFPLA_INST_0_62869 : AXOI3
      port map(A => HIEFFPLA_NET_0_117078, B => 
        HIEFFPLA_NET_0_117073, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[0]\, Y => 
        HIEFFPLA_NET_0_115934);
    
    HIEFFPLA_INST_0_61283 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_19[0]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_20[0]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_4[0]\, Y => 
        HIEFFPLA_NET_0_116148);
    
    \U_ELK8_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]\ : DFN1C0
      port map(D => \U_ELK8_CH/U_SLAVE_1ELK/Q[3]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]_net_1\);
    
    \U_ELK3_CH/U_ELK1_SERDAT_SOURCE/SERDAT[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118100, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_15, Q => 
        \U_ELK3_CH/ELK_TX_DAT[3]\);
    
    HIEFFPLA_INST_0_41765 : MX2
      port map(A => HIEFFPLA_NET_0_119677, B => 
        \U50_PATTERNS/ELINK_RWA[3]\, S => 
        \U50_PATTERNS/SM_BANK_SEL_0[20]\, Y => 
        HIEFFPLA_NET_0_119698);
    
    \U_ELK6_CH/ELK_IN_F\ : DFN1C0
      port map(D => \U_ELK6_CH/ELK_IN_DDR_F\, CLK => CCC_160M_ADJ, 
        CLR => DEV_RST_B_c, Q => \U_ELK6_CH/ELK_IN_F_net_1\);
    
    HIEFFPLA_INST_0_51821 : AOI1D
      port map(A => \U_MASTER_DES/U13A_ADJ_160M/BITCNT[5]\, B => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[4]\, C => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[6]\, Y => 
        HIEFFPLA_NET_0_117687);
    
    \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[73]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117706, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_33, Q => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[73]_net_1\);
    
    \U50_PATTERNS/TFC_ADDRA[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119204, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_9, Q => \U50_PATTERNS/TFC_ADDRA[3]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[7]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_WRD_40M_FIXED[7]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_27, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[7]_net_1\);
    
    \U_ELK16_CH/U_SLAVE_1ELK/RECD_SER_WORD[4]\ : DFN1C0
      port map(D => \U_ELK16_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[4]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_16[4]\);
    
    HIEFFPLA_INST_0_46873 : NAND2B
      port map(A => \OP_MODE_c[1]\, B => \PATT_ELK_DAT_11[1]\, Y
         => HIEFFPLA_NET_0_118597);
    
    HIEFFPLA_INST_0_45965 : NAND3C
      port map(A => HIEFFPLA_NET_0_118946, B => 
        HIEFFPLA_NET_0_118955, C => HIEFFPLA_NET_0_118700, Y => 
        HIEFFPLA_NET_0_118800);
    
    \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_115941, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_24_0, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[1]_net_1\);
    
    \U50_PATTERNS/TFC_STRT_ADDR[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119168, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_13, Q => 
        \U50_PATTERNS/TFC_STRT_ADDR[4]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_7[8]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116595, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_14, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_7[8]\);
    
    \U_ELK14_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0\ : DFN1C0
      port map(D => CLK_40M_GL, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_7, Q => 
        \U_ELK14_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0_net_1\);
    
    HIEFFPLA_INST_0_57008 : AXOI4
      port map(A => HIEFFPLA_NET_0_117085, B => 
        HIEFFPLA_NET_0_117601, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_2[0]\, Y => 
        HIEFFPLA_NET_0_116755);
    
    HIEFFPLA_INST_0_42364 : XOR2
      port map(A => \U50_PATTERNS/RD_XFER_TYPE[1]_net_1\, B => 
        \U50_PATTERNS/RD_XFER_TYPE[0]_net_1\, Y => 
        HIEFFPLA_NET_0_119555);
    
    AFLSDF_INV_26 : INV
      port map(A => DCB_SALT_SEL_c, Y => \AFLSDF_INV_26\);
    
    \U_ELK15_CH/U_ELK1_SERDAT_SOURCE/SERDAT[7]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118411, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_8, Q => 
        \U_ELK15_CH/ELK_TX_DAT[7]\);
    
    \U50_PATTERNS/ELINK_DINA_7[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119731, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_17, Q => 
        \U50_PATTERNS/ELINK_DINA_7[4]\);
    
    \U200B_ELINKS/RX_SER_WORD_1DEL[3]\ : DFN1C0
      port map(D => \ELK_RX_SER_WORD_0[3]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_23, Q => 
        \U200B_ELINKS/RX_SER_WORD_1DEL[3]_net_1\);
    
    HIEFFPLA_INST_0_60684 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_14[2]\, B => 
        HIEFFPLA_NET_0_117181, S => HIEFFPLA_NET_0_117228, Y => 
        HIEFFPLA_NET_0_116233);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_10[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116561, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_6, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_10[1]\);
    
    \U_ELK1_CH/U_ELK1_CMD_TX/SER_OUT_FDEL\ : DFN1P0
      port map(D => \U_ELK1_CH/U_ELK1_CMD_TX/SER_OUT_FI_i\, CLK
         => CCC_160M_FXD, PRE => MASTER_SALT_POR_B_i_0_i_1, Q => 
        \U_ELK1_CH/ELK_OUT_F_i_0\);
    
    \U200B_ELINKS/RX_SER_WORD_1DEL[1]\ : DFN1C0
      port map(D => \ELK_RX_SER_WORD_0[1]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_23, Q => 
        \U200B_ELINKS/RX_SER_WORD_1DEL[1]_net_1\);
    
    HIEFFPLA_INST_0_53254 : XA1B
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[3]\, 
        B => HIEFFPLA_NET_0_115870, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[8]_net_1\, Y => 
        HIEFFPLA_NET_0_117444);
    
    \U_ELK16_CH/U_SLAVE_1ELK/Q[14]\ : DFN1C0
      port map(D => \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[14]_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/Q[14]_net_1\);
    
    HIEFFPLA_INST_0_48648 : MX2
      port map(A => \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[2]_net_1\, 
        B => \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\, S => 
        \BIT_OS_SEL_0[2]\, Y => HIEFFPLA_NET_0_118272);
    
    HIEFFPLA_INST_0_60959 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_1[0]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_17[0]\, S
         => \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_3[4]_net_1\, 
        Y => HIEFFPLA_NET_0_116192);
    
    HIEFFPLA_INST_0_48551 : MX2
      port map(A => HIEFFPLA_NET_0_118294, B => 
        HIEFFPLA_NET_0_118318, S => \BIT_OS_SEL_1[1]\, Y => 
        HIEFFPLA_NET_0_118296);
    
    \U_ELK4_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118062, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_17, Q => 
        \U_ELK4_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]_net_1\);
    
    \U_EXEC_MASTER/MPOR_B_8\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117787, CLK => CLK_40M_GL, CLR
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_1\, Q => 
        P_MASTER_POR_B_c_8);
    
    HIEFFPLA_INST_0_45269 : AO1
      port map(A => HIEFFPLA_NET_0_119236, B => 
        \U50_PATTERNS/ELINK_DOUTA_0[4]\, C => 
        HIEFFPLA_NET_0_118833, Y => HIEFFPLA_NET_0_118954);
    
    \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[4]\ : DFN1C0
      port map(D => \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\);
    
    HIEFFPLA_INST_0_63241 : AND2A
      port map(A => \OP_MODE_c_0[1]\, B => \PATT_TFC_DAT[4]\, Y
         => \U_TFC_SERDAT_SOURCE/N_SERDAT[4]\);
    
    HIEFFPLA_INST_0_49840 : AND2
      port map(A => \U_ELK4_CH/ELK_TX_DAT[1]\, B => 
        \U_ELK4_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118063);
    
    HIEFFPLA_INST_0_47873 : AND2A
      port map(A => \OP_MODE_c_6[1]\, B => \PATT_ELK_DAT_15[5]\, 
        Y => HIEFFPLA_NET_0_118413);
    
    HIEFFPLA_INST_0_47457 : MX2
      port map(A => \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\, 
        B => \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[12]_net_1\, S => 
        \BIT_OS_SEL_3[2]\, Y => HIEFFPLA_NET_0_118489);
    
    HIEFFPLA_INST_0_47146 : MX2
      port map(A => \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\, 
        B => \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\, S => 
        \BIT_OS_SEL_3[2]\, Y => HIEFFPLA_NET_0_118543);
    
    HIEFFPLA_INST_0_45814 : NAND2A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_12[3]\, Y => 
        HIEFFPLA_NET_0_118834);
    
    \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[14]\ : DFN1C0
      port map(D => 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]_net_1\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[14]_net_1\);
    
    HIEFFPLA_INST_0_46967 : MX2
      port map(A => \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\, 
        B => \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[13]_net_1\, S => 
        \BIT_OS_SEL_5[2]\, Y => HIEFFPLA_NET_0_118578);
    
    HIEFFPLA_INST_0_60423 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_9[2]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_10[2]\, S
         => \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_1[0]\, Y
         => HIEFFPLA_NET_0_116268);
    
    \U_ELK6_CH/U_ELK1_CMD_TX/SER_OUT_RI\ : DFN1C0
      port map(D => 
        \U_ELK6_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_3, Q => 
        \U_ELK6_CH/U_ELK1_CMD_TX/SER_OUT_RI_net_1\);
    
    HIEFFPLA_INST_0_52321 : AND3A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[3]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[0]_net_1\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[7]_net_1\, Y => 
        HIEFFPLA_NET_0_117581);
    
    HIEFFPLA_INST_0_48694 : MX2
      port map(A => \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\, 
        B => \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[11]_net_1\, S => 
        \BIT_OS_SEL_0[2]\, Y => HIEFFPLA_NET_0_118265);
    
    HIEFFPLA_INST_0_46698 : MX2
      port map(A => \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\, 
        B => \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[12]_net_1\, S => 
        \BIT_OS_SEL_6[2]\, Y => HIEFFPLA_NET_0_118626);
    
    HIEFFPLA_INST_0_58020 : XA1C
      port map(A => HIEFFPLA_NET_0_116585, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_7[7]\, C => 
        HIEFFPLA_NET_0_117179, Y => HIEFFPLA_NET_0_116577);
    
    HIEFFPLA_INST_0_47623 : AND2A
      port map(A => \OP_MODE_c_2[1]\, B => \PATT_ELK_DAT_14[4]\, 
        Y => HIEFFPLA_NET_0_118459);
    
    HIEFFPLA_INST_0_38525 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_0[3]\, B => 
        HIEFFPLA_NET_0_119520, S => HIEFFPLA_NET_0_119272, Y => 
        HIEFFPLA_NET_0_120092);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_8[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_115968, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_19, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_8[2]\);
    
    \U_ELK13_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL\ : DFN1C0
      port map(D => 
        \U_ELK13_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL_net_1\);
    
    HIEFFPLA_INST_0_57907 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_7[4]\, B => 
        HIEFFPLA_NET_0_116580, S => HIEFFPLA_NET_0_117113, Y => 
        HIEFFPLA_NET_0_116599);
    
    HIEFFPLA_INST_0_56463 : AOI1D
      port map(A => HIEFFPLA_NET_0_117432, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_SEL[3]_net_1\, C
         => \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[5]_net_1\, Y
         => HIEFFPLA_NET_0_116859);
    
    HIEFFPLA_INST_0_40459 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_12[1]\, B => 
        HIEFFPLA_NET_0_119576, S => HIEFFPLA_NET_0_119295, Y => 
        HIEFFPLA_NET_0_119846);
    
    \U_EXEC_MASTER/MPOR_B_14\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117787, CLK => CLK_40M_GL, CLR
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_1\, Q => 
        P_MASTER_POR_B_c_14);
    
    HIEFFPLA_INST_0_52014 : MX2
      port map(A => HIEFFPLA_NET_0_117642, B => 
        HIEFFPLA_NET_0_117640, S => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[1]\, Y => 
        HIEFFPLA_NET_0_117652);
    
    \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_115940, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_24_0, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[0]_net_1\);
    
    \U_EXEC_MASTER/PRESCALE[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117765, CLK => CLK_40M_GL, CLR
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i\, Q => 
        \U_EXEC_MASTER/PRESCALE[3]\);
    
    \U_ELK7_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2\ : IOPADN_BI
      port map(DB => \U_ELK7_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, 
        E => \U_ELK7_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET3\, PAD => 
        ELK7_DAT_N, N2POUT => 
        \U_ELK7_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2_N2P\);
    
    HIEFFPLA_INST_0_50182 : MX2
      port map(A => HIEFFPLA_NET_0_117998, B => 
        HIEFFPLA_NET_0_117994, S => \BIT_OS_SEL_6[1]\, Y => 
        HIEFFPLA_NET_0_117996);
    
    \U50_PATTERNS/U4B_REGCROSS/SAMP_ONE[5]\ : DFN1C0
      port map(D => \U50_PATTERNS/TFC_STOP_ADDR[5]\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_25, Q => 
        \U50_PATTERNS/U4B_REGCROSS/SAMP_ONE[5]_net_1\);
    
    HIEFFPLA_INST_0_52746 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_21[2]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_22[2]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[0]\, Y => 
        HIEFFPLA_NET_0_117518);
    
    HIEFFPLA_INST_0_52027 : AND2A
      port map(A => \U_MASTER_DES/U13A_ADJ_160M/BITCNT[0]\, B => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[42]_net_1\, Y => 
        HIEFFPLA_NET_0_117649);
    
    HIEFFPLA_INST_0_112188 : AOI1C
      port map(A => \U200A_TFC/GP_PG_SM[4]_net_1\, B => 
        \U200A_TFC/GP_PG_SM[5]_net_1\, C => HIEFFPLA_NET_0_120293, 
        Y => HIEFFPLA_NET_0_115816);
    
    \U50_PATTERNS/TFC_STRT_ADDR[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119166, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_13, Q => 
        \U50_PATTERNS/TFC_STRT_ADDR[6]\);
    
    HIEFFPLA_INST_0_61934 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_27[3]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_28[3]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[0]\, Y => 
        HIEFFPLA_NET_0_116057);
    
    HIEFFPLA_INST_0_51708 : NAND2B
      port map(A => 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM[4]_net_1\, B => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[1]_net_1\, Y => 
        HIEFFPLA_NET_0_117718);
    
    HIEFFPLA_INST_0_54708 : MX2
      port map(A => HIEFFPLA_NET_0_117308, B => 
        HIEFFPLA_NET_0_117229, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[0]_net_1\, Y => 
        HIEFFPLA_NET_0_117220);
    
    \U_ELK7_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U3\ : IOBI_ID_OD_EB
      port map(DR => \U_ELK7_CH/ELK_OUT_R\, DF => 
        \U_ELK7_CH/ELK_OUT_F\, CLR => \GND\, E => \AFLSDF_INV_47\, 
        ICLK => CCC_160M_ADJ, OCLK => CCC_160M_FXD, YIN => 
        \U_ELK7_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\, DOUT => OPEN, 
        EOUT => \U_ELK7_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET3\, YR
         => OPEN, YF => OPEN);
    
    \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[1]\ : DFN1C0
      port map(D => 
        \U_ELK19_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\);
    
    HIEFFPLA_INST_0_54381 : MX2
      port map(A => HIEFFPLA_NET_0_116153, B => 
        HIEFFPLA_NET_0_116046, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_2[3]_net_1\, Y
         => HIEFFPLA_NET_0_117273);
    
    HIEFFPLA_INST_0_49860 : AND2A
      port map(A => \OP_MODE_c_1[1]\, B => \PATT_ELK_DAT_4[0]\, Y
         => HIEFFPLA_NET_0_118058);
    
    HIEFFPLA_INST_0_48403 : MX2
      port map(A => \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\, 
        B => \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\, S => 
        \BIT_OS_SEL_0[2]\, Y => HIEFFPLA_NET_0_118316);
    
    \U_ELK16_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL\ : DFN1C0
      port map(D => 
        \U_ELK16_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL_net_1\);
    
    \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[3]\ : DFN1C0
      port map(D => \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\);
    
    \U_ELK9_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117835, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_0, Q => 
        \U_ELK9_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]_net_1\);
    
    \U50_PATTERNS/ELINK_DINA_19[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119789, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_0, Q => 
        \U50_PATTERNS/ELINK_DINA_19[2]\);
    
    HIEFFPLA_INST_0_54602 : MX2
      port map(A => HIEFFPLA_NET_0_117301, B => 
        HIEFFPLA_NET_0_117283, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[2]_net_1\, Y => 
        HIEFFPLA_NET_0_117234);
    
    \U50_PATTERNS/ELINK_DINA_18[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119794, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_21, Q => 
        \U50_PATTERNS/ELINK_DINA_18[5]\);
    
    HIEFFPLA_INST_0_63137 : AX1C
      port map(A => HIEFFPLA_NET_0_117125, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[0]_net_1\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[1]_net_1\, Y => 
        HIEFFPLA_NET_0_115879);
    
    HIEFFPLA_INST_0_42781 : AOI1D
      port map(A => HIEFFPLA_NET_0_118992, B => 
        HIEFFPLA_NET_0_119006, C => 
        \U50_PATTERNS/REG_STATE_0[5]_net_1\, Y => 
        HIEFFPLA_NET_0_119464);
    
    HIEFFPLA_INST_0_41716 : MX2
      port map(A => HIEFFPLA_NET_0_119685, B => 
        \U50_PATTERNS/ELINK_RWA[15]\, S => 
        \U50_PATTERNS/SM_BANK_SEL_0[20]\, Y => 
        HIEFFPLA_NET_0_119705);
    
    HIEFFPLA_INST_0_53854 : MX2
      port map(A => HIEFFPLA_NET_0_117282, B => 
        HIEFFPLA_NET_0_117198, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[2]_net_1\, Y
         => HIEFFPLA_NET_0_117342);
    
    HIEFFPLA_INST_0_44538 : XOR2
      port map(A => \ELKS_STRT_ADDR[1]\, B => 
        \U50_PATTERNS/U4C_REGCROSS/SAMP_TWO[1]_net_1\, Y => 
        HIEFFPLA_NET_0_119097);
    
    HIEFFPLA_INST_0_49364 : NAND2B
      port map(A => \OP_MODE_c_1[1]\, B => \PATT_ELK_DAT_2[2]\, Y
         => HIEFFPLA_NET_0_118146);
    
    HIEFFPLA_INST_0_60618 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_13[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_29[1]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_2[4]_net_1\, Y
         => HIEFFPLA_NET_0_116243);
    
    HIEFFPLA_INST_0_38085 : NAND3C
      port map(A => HIEFFPLA_NET_0_120155, B => 
        \U200B_ELINKS/RX_SER_WORD_3DEL[4]_net_1\, C => 
        \U200B_ELINKS/RX_SER_WORD_3DEL[5]_net_1\, Y => 
        HIEFFPLA_NET_0_120156);
    
    HIEFFPLA_INST_0_42288 : NAND3C
      port map(A => \U50_PATTERNS/RD_USB_ADBUS[3]\, B => 
        \U50_PATTERNS/RD_USB_ADBUS[2]\, C => 
        \U50_PATTERNS/RD_USB_ADBUS[4]\, Y => 
        HIEFFPLA_NET_0_119581);
    
    HIEFFPLA_INST_0_58097 : MX2
      port map(A => HIEFFPLA_NET_0_116687, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_0[2]\, S => 
        HIEFFPLA_NET_0_117201, Y => HIEFFPLA_NET_0_116564);
    
    \U_REFCLKBUF/_BIBUF_LVDS[0]_/U0/U3\ : IOBI_IB_OB_EB
      port map(D => CLK_40M_GL, E => DCB_SALT_SEL_c, YIN => 
        \U_REFCLKBUF/\\\\BIBUF_LVDS[0]\\\\/U0/NET4\, DOUT => OPEN, 
        EOUT => \U_REFCLKBUF/\\\\BIBUF_LVDS[0]\\\\/U0/NET3\, Y
         => OPEN);
    
    HIEFFPLA_INST_0_43783 : AND3A
      port map(A => HIEFFPLA_NET_0_119585, B => 
        HIEFFPLA_NET_0_119562, C => HIEFFPLA_NET_0_119597, Y => 
        HIEFFPLA_NET_0_119215);
    
    \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[3]\ : DFN1C0
      port map(D => 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[3]_net_1\);
    
    \U_ELK6_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]\ : DFN1C0
      port map(D => \U_ELK6_CH/U_SLAVE_1ELK/Q[7]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]_net_1\);
    
    HIEFFPLA_INST_0_54741 : NAND3B
      port map(A => HIEFFPLA_NET_0_117246, B => 
        HIEFFPLA_NET_0_117252, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[1]_net_1\, Y => 
        HIEFFPLA_NET_0_117211);
    
    HIEFFPLA_INST_0_51411 : NAND2A
      port map(A => DCB_SALT_SEL_c, B => HIEFFPLA_NET_0_117787, Y
         => HIEFFPLA_NET_0_117781);
    
    \U_ELK2_CH/U_SLAVE_1ELK/Q[2]\ : DFN1C0
      port map(D => \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/Q[2]_net_1\);
    
    \U_ELK13_CH/U_ELK1_CMD_TX/SER_OUT_RDEL\ : DFN1C0
      port map(D => \U_ELK13_CH/U_ELK1_CMD_TX/SER_OUT_RI_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_1, Q
         => \U_ELK13_CH/ELK_OUT_R\);
    
    \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[2]\ : DFN1C0
      port map(D => 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[2]_net_1\);
    
    \U_ELK2_CH/U_SLAVE_1ELK/RECD_SER_WORD[4]\ : DFN1C0
      port map(D => \U_ELK2_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[4]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_2[4]\);
    
    \U_ELK1_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]\ : DFN1C0
      port map(D => \U_ELK1_CH/U_SLAVE_1ELK/Q[1]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]_net_1\);
    
    ELK0_IN_F : DFN1C0
      port map(D => \AFLSDF_INV_57\, CLK => CCC_160M_ADJ, CLR => 
        DEV_RST_B_c, Q => \ELK0_IN_F\);
    
    \U200B_ELINKS/RX_SER_WORD_3DEL[7]\ : DFN1P0
      port map(D => \AFLSDF_INV_58\, CLK => CLK_40M_GL, PRE => 
        P_MASTER_POR_B_c_31_0, Q => 
        \U200B_ELINKS/RX_SER_WORD_3DEL_i_0[7]\);
    
    \U50_PATTERNS/ELINK_DINA_12[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119846, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_12, Q => 
        \U50_PATTERNS/ELINK_DINA_12[1]\);
    
    \U200A_TFC/ADDR_POINTER[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120364, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_30, Q => \TFC_ADDRB[2]\);
    
    HIEFFPLA_INST_0_44158 : MX2
      port map(A => \U50_PATTERNS/TFC_STRT_ADDR[6]\, B => 
        \U50_PATTERNS/TFC_STRT_ADDR_T[6]\, S => 
        HIEFFPLA_NET_0_119472, Y => HIEFFPLA_NET_0_119166);
    
    \U50_PATTERNS/SM_BANK_SEL[19]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119312, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_1_0, Q => 
        \U50_PATTERNS/SM_BANK_SEL[19]\);
    
    HIEFFPLA_INST_0_57274 : NAND3A
      port map(A => HIEFFPLA_NET_0_116712, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_3[7]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_3[6]\, Y => 
        HIEFFPLA_NET_0_116709);
    
    HIEFFPLA_INST_0_50551 : MX2
      port map(A => HIEFFPLA_NET_0_117947, B => 
        HIEFFPLA_NET_0_117933, S => \BIT_OS_SEL_6[1]\, Y => 
        HIEFFPLA_NET_0_117935);
    
    \U_EXEC_MASTER/MPOR_B_0\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117787, CLK => CLK_40M_GL, CLR
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_2\, Q => 
        \U_EXEC_MASTER/P_MASTER_POR_B_c_0\);
    
    \U50_PATTERNS/ELINK_DINA_8[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119723, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_18, Q => 
        \U50_PATTERNS/ELINK_DINA_8[4]\);
    
    HIEFFPLA_INST_0_37610 : AO1A
      port map(A => HIEFFPLA_NET_0_120239, B => 
        HIEFFPLA_NET_0_120234, C => HIEFFPLA_NET_0_120236, Y => 
        HIEFFPLA_NET_0_120247);
    
    \U50_PATTERNS/ELINK_ADDRA_9[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119939, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_10, Q => 
        \U50_PATTERNS/ELINK_ADDRA_9[4]\);
    
    \U200B_ELINKS/LOC_STRT_ADDR[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120173, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_12, Q => 
        \U200B_ELINKS/LOC_STRT_ADDR[6]\);
    
    HIEFFPLA_INST_0_55738 : MX2
      port map(A => HIEFFPLA_NET_0_117019, B => 
        HIEFFPLA_NET_0_117007, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[2]\, Y => 
        HIEFFPLA_NET_0_116996);
    
    HIEFFPLA_INST_0_50369 : MX2
      port map(A => HIEFFPLA_NET_0_117949, B => 
        HIEFFPLA_NET_0_117947, S => \BIT_OS_SEL_5[1]\, Y => 
        HIEFFPLA_NET_0_117960);
    
    HIEFFPLA_INST_0_43998 : MX2
      port map(A => \U50_PATTERNS/TFC_STOP_ADDR[2]\, B => 
        \U50_PATTERNS/TFC_STOP_ADDR_T[2]\, S => 
        HIEFFPLA_NET_0_119472, Y => HIEFFPLA_NET_0_119186);
    
    \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[7]\ : DFN1C0
      port map(D => \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\);
    
    HIEFFPLA_INST_0_47515 : MX2
      port map(A => HIEFFPLA_NET_0_118486, B => 
        HIEFFPLA_NET_0_118498, S => \BIT_OS_SEL_4[0]\, Y => 
        \U_ELK13_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[3]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_24[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116102, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_8, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_24[3]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_SEL_4[0]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_BIT_OS_VAL[0]\, CLK
         => CLK_40M_GL, CLR => P_MASTER_POR_B_c_27_0, Q => 
        \BIT_OS_SEL_4[0]\);
    
    \U50_PATTERNS/ELINK_ADDRA_17[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120025, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_11, Q => 
        \U50_PATTERNS/ELINK_ADDRA_17[6]\);
    
    HIEFFPLA_INST_0_54504 : MX2
      port map(A => HIEFFPLA_NET_0_116332, B => 
        HIEFFPLA_NET_0_116387, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[3]_net_1\, Y => 
        HIEFFPLA_NET_0_117257);
    
    HIEFFPLA_INST_0_47377 : NAND2B
      port map(A => \OP_MODE_c[1]\, B => \PATT_ELK_DAT_13[7]\, Y
         => HIEFFPLA_NET_0_118501);
    
    HIEFFPLA_INST_0_58033 : AOI1A
      port map(A => HIEFFPLA_NET_0_116590, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_7[5]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_7[6]\, Y => 
        HIEFFPLA_NET_0_116574);
    
    HIEFFPLA_INST_0_51449 : AX1A
      port map(A => HIEFFPLA_NET_0_117785, B => 
        \U_EXEC_MASTER/DEL_CNT[5]\, C => 
        \U_EXEC_MASTER/DEL_CNT[6]\, Y => HIEFFPLA_NET_0_117771);
    
    HIEFFPLA_INST_0_44859 : NAND3C
      port map(A => HIEFFPLA_NET_0_119027, B => 
        HIEFFPLA_NET_0_119421, C => HIEFFPLA_NET_0_119588, Y => 
        HIEFFPLA_NET_0_119033);
    
    \U_ELK19_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]\ : DFN1C0
      port map(D => \U_ELK19_CH/U_SLAVE_1ELK/Q[4]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]_net_1\);
    
    \U50_PATTERNS/ELINK_BLKA[3]/U1\ : DFN1P0
      port map(D => HIEFFPLA_NET_0_119922, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_19, Q => 
        \U50_PATTERNS/ELINK_BLKA[3]\);
    
    HIEFFPLA_INST_0_41879 : AND2
      port map(A => HIEFFPLA_NET_0_119389, B => 
        \U50_PATTERNS/SM_BANK_SEL[16]\, Y => 
        HIEFFPLA_NET_0_119676);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_1[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116167, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_8, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_1[3]\);
    
    \U_ELK8_CH/U_ELK1_SERDAT_SOURCE/SERDAT[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117878, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_5, Q => 
        \U_ELK8_CH/ELK_TX_DAT[0]\);
    
    \U_ELK14_CH/U_SLAVE_1ELK/Q[3]\ : DFN1C0
      port map(D => \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/Q[3]_net_1\);
    
    HIEFFPLA_INST_0_61205 : MX2
      port map(A => HIEFFPLA_NET_0_117167, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_20[1]\, S => 
        HIEFFPLA_NET_0_117141, Y => HIEFFPLA_NET_0_116159);
    
    HIEFFPLA_INST_0_48654 : MX2
      port map(A => \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[3]_net_1\, 
        B => \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\, S => 
        \BIT_OS_SEL_0[2]\, Y => HIEFFPLA_NET_0_118271);
    
    \U_ELK9_CH/U_SLAVE_1ELK/Q[9]\ : DFN1C0
      port map(D => \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/Q[9]_net_1\);
    
    HIEFFPLA_INST_0_51536 : AO1C
      port map(A => 
        \U_EXEC_MASTER/USB_MASTER_EN/TEST_SM[1]_net_1\, B => 
        \U_EXEC_MASTER/USB_MASTER_EN/TEST_SM_i_0[2]\, C => 
        \U_EXEC_MASTER/USB_MASTER_EN/TERMCNT_FG40M2S_net_1\, Y
         => HIEFFPLA_NET_0_117751);
    
    \U50_PATTERNS/ELINK_ADDRA_15[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120047, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_6, Q => 
        \U50_PATTERNS/ELINK_ADDRA_15[0]\);
    
    HIEFFPLA_INST_0_57389 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_4[5]\, B => 
        HIEFFPLA_NET_0_116666, S => HIEFFPLA_NET_0_117122, Y => 
        HIEFFPLA_NET_0_116691);
    
    HIEFFPLA_INST_0_51532 : MX2B
      port map(A => 
        \U_EXEC_MASTER/USB_MASTER_EN/TEST_SM[0]_net_1\, B => 
        \U_EXEC_MASTER/USB_MASTER_EN/TERMCNT_FG40M2S_net_1\, S
         => \U_EXEC_MASTER/USB_MASTER_EN/TEST_SM[1]_net_1\, Y => 
        HIEFFPLA_NET_0_117752);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_15[4]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116226, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_4, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_15[4]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_SEL[2]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_BIT_OS_VAL[2]\, CLK
         => CLK_40M_GL, CLR => P_MASTER_POR_B_c_27_1, Q => 
        \BIT_OS_SEL[2]\);
    
    \U_ELK4_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118063, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_16, Q => 
        \U_ELK4_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]_net_1\);
    
    \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[9]\ : DFN1C0
      port map(D => 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\);
    
    HIEFFPLA_INST_0_111823 : AX1E
      port map(A => HIEFFPLA_NET_0_117747, B => 
        \U_EXEC_MASTER/USB_MASTER_EN/T_CNT60M[4]_net_1\, C => 
        \U_EXEC_MASTER/USB_MASTER_EN/T_CNT60M[5]_net_1\, Y => 
        HIEFFPLA_NET_0_115828);
    
    \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_3[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_116999, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_16_0, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_3[0]\);
    
    \U_ELK1_CH/U_SLAVE_1ELK/Q[0]\ : DFN1C0
      port map(D => \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/Q[0]_net_1\);
    
    HIEFFPLA_INST_0_51138 : MX2
      port map(A => HIEFFPLA_NET_0_117819, B => 
        HIEFFPLA_NET_0_117816, S => \BIT_OS_SEL_3[1]\, Y => 
        HIEFFPLA_NET_0_117822);
    
    \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[0]\ : DFN1C0
      port map(D => 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[0]_net_1\);
    
    \U_ELK7_CH/U_SLAVE_1ELK/Q[11]\ : DFN1C0
      port map(D => \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/Q[11]_net_1\);
    
    HIEFFPLA_INST_0_61697 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_25[4]\, B => 
        HIEFFPLA_NET_0_117166, S => HIEFFPLA_NET_0_117117, Y => 
        HIEFFPLA_NET_0_116091);
    
    HIEFFPLA_INST_0_37946 : MX2
      port map(A => \U200B_ELINKS/LOC_STOP_ADDR[2]\, B => 
        \ELKS_STOP_ADDR[2]\, S => 
        \U200B_ELINKS/GP_PG_SM_0[10]_net_1\, Y => 
        HIEFFPLA_NET_0_120185);
    
    HIEFFPLA_INST_0_40801 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_16[7]\, B => 
        HIEFFPLA_NET_0_119560, S => HIEFFPLA_NET_0_119257, Y => 
        HIEFFPLA_NET_0_119808);
    
    HIEFFPLA_INST_0_57098 : NAND2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_2[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_2[2]\, Y => 
        HIEFFPLA_NET_0_116745);
    
    HIEFFPLA_INST_0_40711 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_15[5]\, B => 
        HIEFFPLA_NET_0_119567, S => HIEFFPLA_NET_0_119297, Y => 
        HIEFFPLA_NET_0_119818);
    
    HIEFFPLA_INST_0_53166 : MX2
      port map(A => HIEFFPLA_NET_0_117537, B => 
        HIEFFPLA_NET_0_117533, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_1[3]\, Y => 
        HIEFFPLA_NET_0_117457);
    
    HIEFFPLA_INST_0_48618 : NAND2B
      port map(A => \OP_MODE_c_1[1]\, B => \PATT_ELK_DAT_18[3]\, 
        Y => HIEFFPLA_NET_0_118280);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_5[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116661, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_11, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_5[0]\);
    
    HIEFFPLA_INST_0_56197 : XA1C
      port map(A => HIEFFPLA_NET_0_116945, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/MAX_CNT[7]\, C => 
        HIEFFPLA_NET_0_117112, Y => HIEFFPLA_NET_0_116932);
    
    HIEFFPLA_INST_0_49591 : AND2
      port map(A => \U_ELK3_CH/ELK_TX_DAT[1]\, B => 
        \U_ELK3_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118108);
    
    HIEFFPLA_INST_0_54573 : AND2A
      port map(A => HIEFFPLA_NET_0_116620, B => 
        HIEFFPLA_NET_0_117208, Y => HIEFFPLA_NET_0_117243);
    
    \U_ELK7_CH/U_ELK1_CMD_TX/SER_OUT_RI\ : DFN1C0
      port map(D => 
        \U_ELK7_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_13, Q
         => \U_ELK7_CH/U_ELK1_CMD_TX/SER_OUT_RI_net_1\);
    
    \U_ELK2_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]\ : DFN1C0
      port map(D => \U_ELK2_CH/U_SLAVE_1ELK/Q[5]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]_net_1\);
    
    \U50_PATTERNS/U4A_REGCROSS/SAMP_TWO[5]\ : DFN1C0
      port map(D => \U50_PATTERNS/U4A_REGCROSS/SAMP_ONE[5]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_22, Q => 
        \U50_PATTERNS/U4A_REGCROSS/SAMP_TWO[5]_net_1\);
    
    HIEFFPLA_INST_0_39497 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_3[7]\, B => 
        HIEFFPLA_NET_0_119516, S => HIEFFPLA_NET_0_119247, Y => 
        HIEFFPLA_NET_0_119984);
    
    HIEFFPLA_INST_0_62239 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_31[2]\, B => 
        HIEFFPLA_NET_0_117181, S => HIEFFPLA_NET_0_117319, Y => 
        HIEFFPLA_NET_0_116018);
    
    HIEFFPLA_INST_0_40112 : AOI1C
      port map(A => \U50_PATTERNS/ELINK_BLKA[16]\, B => 
        HIEFFPLA_NET_0_119653, C => HIEFFPLA_NET_0_119901, Y => 
        HIEFFPLA_NET_0_119902);
    
    HIEFFPLA_INST_0_50354 : MX2
      port map(A => 
        \U_ELK6_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]_net_1\, B => 
        \U_ELK6_CH/ELK_TX_DAT[7]\, S => 
        \U_ELK6_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_117970);
    
    \U_ELK10_CH/U_ELK1_CMD_TX/SER_OUT_RDEL\ : DFN1C0
      port map(D => \U_ELK10_CH/U_ELK1_CMD_TX/SER_OUT_RI_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_5, Q
         => \U_ELK10_CH/ELK_OUT_R\);
    
    \U50_PATTERNS/ELINK_DINA_19[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119785, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_1, Q => 
        \U50_PATTERNS/ELINK_DINA_19[6]\);
    
    \U_MASTER_DES/U13A_ADJ_160M/BITCNT[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117697, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_14, Q => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[1]\);
    
    HIEFFPLA_INST_0_57490 : XA1B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_4[0]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_4[1]\, C => 
        HIEFFPLA_NET_0_117179, Y => HIEFFPLA_NET_0_116670);
    
    HIEFFPLA_INST_0_58813 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_1[2]\, B => 
        HIEFFPLA_NET_0_116469, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_1[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116473);
    
    \U_ELK8_CH/U_SLAVE_1ELK/Q[3]\ : DFN1C0
      port map(D => \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/Q[3]_net_1\);
    
    \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[4]\ : DFN1C0
      port map(D => \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\);
    
    \U_ELK4_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]\ : DFN1C0
      port map(D => \U_ELK4_CH/U_SLAVE_1ELK/Q[10]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]_net_1\);
    
    HIEFFPLA_INST_0_57399 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_4[6]\, B => 
        HIEFFPLA_NET_0_116665, S => HIEFFPLA_NET_0_117122, Y => 
        HIEFFPLA_NET_0_116690);
    
    HIEFFPLA_INST_0_55385 : AO1
      port map(A => HIEFFPLA_NET_0_117087, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[0]\, C => 
        HIEFFPLA_NET_0_116997, Y => HIEFFPLA_NET_0_117045);
    
    \U50_PATTERNS/U119_PATT_ELINK_BLK/DPRT_512X9_SRAM_R0C0\ : 
        RAM4K9
      generic map(MEMORYFILE => "DPRT_512X9_SRAM_R0C0.mem")

      port map(ADDRA11 => AFLSDF_GND, ADDRA10 => AFLSDF_GND, 
        ADDRA9 => AFLSDF_GND, ADDRA8 => \GND\, ADDRA7 => 
        \U50_PATTERNS/ELINK_ADDRA_19[7]\, ADDRA6 => 
        \U50_PATTERNS/ELINK_ADDRA_19[6]\, ADDRA5 => 
        \U50_PATTERNS/ELINK_ADDRA_19[5]\, ADDRA4 => 
        \U50_PATTERNS/ELINK_ADDRA_19[4]\, ADDRA3 => 
        \U50_PATTERNS/ELINK_ADDRA_19[3]\, ADDRA2 => 
        \U50_PATTERNS/ELINK_ADDRA_19[2]\, ADDRA1 => 
        \U50_PATTERNS/ELINK_ADDRA_19[1]\, ADDRA0 => 
        \U50_PATTERNS/ELINK_ADDRA_19[0]\, ADDRB11 => AFLSDF_GND, 
        ADDRB10 => AFLSDF_GND, ADDRB9 => AFLSDF_GND, ADDRB8 => 
        \GND\, ADDRB7 => \ELKS_ADDRB[7]\, ADDRB6 => 
        \ELKS_ADDRB[6]\, ADDRB5 => \ELKS_ADDRB[5]\, ADDRB4 => 
        \ELKS_ADDRB[4]\, ADDRB3 => \ELKS_ADDRB[3]\, ADDRB2 => 
        \ELKS_ADDRB[2]\, ADDRB1 => \ELKS_ADDRB[1]\, ADDRB0 => 
        \ELKS_ADDRB[0]\, DINA8 => \GND\, DINA7 => 
        \U50_PATTERNS/ELINK_DINA_19[7]\, DINA6 => 
        \U50_PATTERNS/ELINK_DINA_19[6]\, DINA5 => 
        \U50_PATTERNS/ELINK_DINA_19[5]\, DINA4 => 
        \U50_PATTERNS/ELINK_DINA_19[4]\, DINA3 => 
        \U50_PATTERNS/ELINK_DINA_19[3]\, DINA2 => 
        \U50_PATTERNS/ELINK_DINA_19[2]\, DINA1 => 
        \U50_PATTERNS/ELINK_DINA_19[1]\, DINA0 => 
        \U50_PATTERNS/ELINK_DINA_19[0]\, DINB8 => \GND\, DINB7
         => \ELK_RX_SER_WORD_19[7]\, DINB6 => 
        \ELK_RX_SER_WORD_19[6]\, DINB5 => \ELK_RX_SER_WORD_19[5]\, 
        DINB4 => \ELK_RX_SER_WORD_19[4]\, DINB3 => 
        \ELK_RX_SER_WORD_19[3]\, DINB2 => \ELK_RX_SER_WORD_19[2]\, 
        DINB1 => \ELK_RX_SER_WORD_19[1]\, DINB0 => 
        \ELK_RX_SER_WORD_19[0]\, WIDTHA0 => \VCC\, WIDTHA1 => 
        \VCC\, WIDTHB0 => \VCC\, WIDTHB1 => \VCC\, PIPEA => \VCC\, 
        PIPEB => \VCC\, WMODEA => \GND\, WMODEB => \GND\, BLKA
         => \U50_PATTERNS/ELINK_BLKA[19]\, BLKB => 
        ELKS_RAM_BLKB_EN, WENA => \U50_PATTERNS/ELINK_RWA[19]\, 
        WENB => ELKS_RWB, CLKA => CLK60MHZ, CLKB => CLK_40M_GL, 
        RESET => P_USB_MASTER_EN_c_0, DOUTA8 => OPEN, DOUTA7 => 
        \U50_PATTERNS/ELINK_DOUTA_19[7]\, DOUTA6 => 
        \U50_PATTERNS/ELINK_DOUTA_19[6]\, DOUTA5 => 
        \U50_PATTERNS/ELINK_DOUTA_19[5]\, DOUTA4 => 
        \U50_PATTERNS/ELINK_DOUTA_19[4]\, DOUTA3 => 
        \U50_PATTERNS/ELINK_DOUTA_19[3]\, DOUTA2 => 
        \U50_PATTERNS/ELINK_DOUTA_19[2]\, DOUTA1 => 
        \U50_PATTERNS/ELINK_DOUTA_19[1]\, DOUTA0 => 
        \U50_PATTERNS/ELINK_DOUTA_19[0]\, DOUTB8 => OPEN, DOUTB7
         => \PATT_ELK_DAT_19[7]\, DOUTB6 => \PATT_ELK_DAT_19[6]\, 
        DOUTB5 => \PATT_ELK_DAT_19[5]\, DOUTB4 => 
        \PATT_ELK_DAT_19[4]\, DOUTB3 => \PATT_ELK_DAT_19[3]\, 
        DOUTB2 => \PATT_ELK_DAT_19[2]\, DOUTB1 => 
        \PATT_ELK_DAT_19[1]\, DOUTB0 => \PATT_ELK_DAT_19[0]\);
    
    \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[42]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117710, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_33, Q => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[42]_net_1\);
    
    \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[9]\ : DFN1C0
      port map(D => 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\);
    
    \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[7]\ : DFN1C0
      port map(D => 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\);
    
    HIEFFPLA_INST_0_37132 : AND3B
      port map(A => \U200A_TFC/LOC_STRT_ADDR[7]\, B => 
        HIEFFPLA_NET_0_120293, C => HIEFFPLA_NET_0_120328, Y => 
        HIEFFPLA_NET_0_120341);
    
    \U_ELK19_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2\ : IOPADN_BI
      port map(DB => \U_ELK19_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, 
        E => \U_ELK19_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET3\, PAD
         => ELK19_DAT_N, N2POUT => 
        \U_ELK19_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2_N2P\);
    
    \U_ELK16_CH/U_SLAVE_1ELK/Q[3]\ : DFN1C0
      port map(D => \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/Q[3]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_21[4]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116141, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_3, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_21[4]\);
    
    \U_EXEC_MASTER/USB_MASTER_EN/T_CNT60M[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117742, CLK => CLK60MHZ, CLR
         => P_MASTER_POR_B_c_28, Q => 
        \U_EXEC_MASTER/USB_MASTER_EN/T_CNT60M[1]_net_1\);
    
    \U50_PATTERNS/ELINK_ADDRA_1[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120001, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_20, Q => 
        \U50_PATTERNS/ELINK_ADDRA_1[6]\);
    
    HIEFFPLA_INST_0_43678 : NAND3C
      port map(A => HIEFFPLA_NET_0_119273, B => 
        HIEFFPLA_NET_0_119252, C => HIEFFPLA_NET_0_119274, Y => 
        HIEFFPLA_NET_0_119245);
    
    HIEFFPLA_INST_0_45777 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_18[0]\, C => 
        \U50_PATTERNS/SM_BANK_SEL[1]\, Y => HIEFFPLA_NET_0_118845);
    
    \U_ELK17_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118333, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_14, Q => 
        \U_ELK17_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]_net_1\);
    
    HIEFFPLA_INST_0_63033 : AND2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[7]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[3]\, Y => 
        HIEFFPLA_NET_0_115908);
    
    HIEFFPLA_INST_0_50608 : NAND2B
      port map(A => \OP_MODE_c_4[1]\, B => \PATT_ELK_DAT_7[1]\, Y
         => HIEFFPLA_NET_0_117922);
    
    \P_OP_MODE5_AAE_pad/U0/U1\ : IOTRI_OB_EB
      port map(D => \OP_MODE_c[5]\, E => \VCC\, DOUT => 
        \P_OP_MODE5_AAE_pad/U0/NET1\, EOUT => 
        \P_OP_MODE5_AAE_pad/U0/NET2\);
    
    HIEFFPLA_INST_0_47662 : MX2
      port map(A => HIEFFPLA_NET_0_118449, B => 
        HIEFFPLA_NET_0_118445, S => \BIT_OS_SEL_2[1]\, Y => 
        HIEFFPLA_NET_0_118450);
    
    HIEFFPLA_INST_0_63120 : NOR2A
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[12]\, 
        B => HIEFFPLA_NET_0_115912, Y => HIEFFPLA_NET_0_115883);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_27[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116068, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_13, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_27[2]\);
    
    HIEFFPLA_INST_0_45388 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/SM_BANK_SEL[9]\, C => 
        \U50_PATTERNS/ELINK_DOUTA_10[7]\, Y => 
        HIEFFPLA_NET_0_118923);
    
    HIEFFPLA_INST_0_41903 : AOI1B
      port map(A => HIEFFPLA_NET_0_119389, B => 
        \U50_PATTERNS/SM_BANK_SEL[11]\, C => 
        HIEFFPLA_NET_0_119639, Y => HIEFFPLA_NET_0_119668);
    
    \U_ELK12_CH/U_SLAVE_1ELK/Q[1]\ : DFN1C0
      port map(D => \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/Q[1]_net_1\);
    
    HIEFFPLA_INST_0_62119 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_2[2]\, 
        B => HIEFFPLA_NET_0_117181, S => HIEFFPLA_NET_0_117176, Y
         => HIEFFPLA_NET_0_116033);
    
    HIEFFPLA_INST_0_46472 : AO1A
      port map(A => HIEFFPLA_NET_0_119571, B => 
        HIEFFPLA_NET_0_119579, C => HIEFFPLA_NET_0_118683, Y => 
        HIEFFPLA_NET_0_118684);
    
    HIEFFPLA_INST_0_51957 : MX2A
      port map(A => HIEFFPLA_NET_0_117650, B => 
        HIEFFPLA_NET_0_117649, S => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[1]\, Y => 
        HIEFFPLA_NET_0_117659);
    
    HIEFFPLA_INST_0_46951 : MX2
      port map(A => HIEFFPLA_NET_0_118584, B => 
        HIEFFPLA_NET_0_118578, S => \BIT_OS_SEL_5[1]\, Y => 
        HIEFFPLA_NET_0_118580);
    
    \U50_PATTERNS/ELINK_ADDRA_14[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120049, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_5, Q => 
        \U50_PATTERNS/ELINK_ADDRA_14[6]\);
    
    HIEFFPLA_INST_0_40324 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_10[2]\, B => 
        HIEFFPLA_NET_0_119575, S => HIEFFPLA_NET_0_119239, Y => 
        HIEFFPLA_NET_0_119861);
    
    \U_ELK6_CH/U_SLAVE_1ELK/RECD_SER_WORD[4]\ : DFN1C0
      port map(D => \U_ELK6_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[4]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_6[4]\);
    
    \U_ELK17_CH/U_SLAVE_1ELK/RECD_SER_WORD[4]\ : DFN1C0
      port map(D => \U_ELK17_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[4]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_17[4]\);
    
    HIEFFPLA_INST_0_58839 : MX2
      port map(A => HIEFFPLA_NET_0_116687, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_1[2]\, S => 
        HIEFFPLA_NET_0_117216, Y => HIEFFPLA_NET_0_116469);
    
    HIEFFPLA_INST_0_45773 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/SM_BANK_SEL[6]\, C => 
        \U50_PATTERNS/ELINK_DOUTA_13[6]\, Y => 
        HIEFFPLA_NET_0_118847);
    
    HIEFFPLA_INST_0_113074 : AO18
      port map(A => HIEFFPLA_NET_0_115810, B => 
        \U200A_TFC/LOC_STOP_ADDR[6]\, C => \TFC_ADDRB[6]\, Y => 
        HIEFFPLA_NET_0_115817);
    
    \U50_PATTERNS/WR_USB_ADBUS[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118981, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_15, Q => 
        \U50_PATTERNS/WR_USB_ADBUS[4]\);
    
    \U_ELK8_CH/U_SLAVE_1ELK/Q[5]\ : DFN1C0
      port map(D => \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/Q[5]_net_1\);
    
    \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[6]\ : DFN1C0
      port map(D => \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\);
    
    HIEFFPLA_INST_0_63242 : AND2A
      port map(A => \OP_MODE_c_0[1]\, B => \PATT_TFC_DAT[5]\, Y
         => \U_TFC_SERDAT_SOURCE/N_SERDAT[5]\);
    
    HIEFFPLA_INST_0_41314 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_5[0]\, B => 
        HIEFFPLA_NET_0_119578, S => HIEFFPLA_NET_0_119251, Y => 
        HIEFFPLA_NET_0_119751);
    
    AFLSDF_INV_59 : INV
      port map(A => \U200A_TFC/RX_SER_WORD_2DEL[7]_net_1\, Y => 
        \AFLSDF_INV_59\);
    
    \U50_PATTERNS/TFC_ADDRA[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119202, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_10, Q => 
        \U50_PATTERNS/TFC_ADDRA[5]\);
    
    \U50_PATTERNS/ELINKS_STRT_ADDR[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120110, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_17, Q => 
        \U50_PATTERNS/ELINKS_STRT_ADDR[1]\);
    
    HIEFFPLA_INST_0_52740 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_21[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_22[1]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[0]\, Y => 
        HIEFFPLA_NET_0_117519);
    
    \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[14]\ : DFN1C0
      port map(D => 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[14]_net_1\);
    
    \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[14]\ : DFN1C0
      port map(D => \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\, 
        CLK => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[14]_net_1\);
    
    HIEFFPLA_INST_0_39425 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_2[7]\, B => 
        HIEFFPLA_NET_0_119516, S => HIEFFPLA_NET_0_119278, Y => 
        HIEFFPLA_NET_0_119992);
    
    \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[9]\ : DFN1C0
      port map(D => \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\);
    
    \U_ELK7_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117932, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_14, Q => 
        \U_ELK7_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]_net_1\);
    
    HIEFFPLA_INST_0_56566 : AND3
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[8]_net_1\, B => 
        HIEFFPLA_NET_0_117426, C => HIEFFPLA_NET_0_117425, Y => 
        HIEFFPLA_NET_0_116837);
    
    HIEFFPLA_INST_0_54890 : NAND2A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_0[6]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_0[8]_net_1\, Y => 
        HIEFFPLA_NET_0_117180);
    
    HIEFFPLA_INST_0_44444 : AND2A
      port map(A => \U50_PATTERNS/U4C_REGCROSS/DELCNT[0]_net_1\, 
        B => \U50_PATTERNS/U4C_REGCROSS/SYNC_SM[0]_net_1\, Y => 
        HIEFFPLA_NET_0_119113);
    
    \U_ELK16_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]\ : DFN1C0
      port map(D => \U_ELK16_CH/U_SLAVE_1ELK/Q[8]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]_net_1\);
    
    \U50_PATTERNS/ELINK_RWA[17]/U1\ : DFN1P0
      port map(D => HIEFFPLA_NET_0_119703, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_12, Q => 
        \U50_PATTERNS/ELINK_RWA[17]\);
    
    \U50_PATTERNS/ELINK_BLKA[18]/U1\ : DFN1P0
      port map(D => HIEFFPLA_NET_0_119926, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_20, Q => 
        \U50_PATTERNS/ELINK_BLKA[18]\);
    
    HIEFFPLA_INST_0_52144 : NAND3B
      port map(A => HIEFFPLA_NET_0_117683, B => 
        HIEFFPLA_NET_0_117688, C => 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM[0]_net_1\, Y => 
        HIEFFPLA_NET_0_117626);
    
    \U50_PATTERNS/ELINK_DINA_13[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119837, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_14, Q => 
        \U50_PATTERNS/ELINK_DINA_13[2]\);
    
    \U_EXEC_MASTER/MPOR_SALT_B_9\ : DFI1P0
      port map(D => HIEFFPLA_NET_0_117781, CLK => CLK_40M_GL, PRE
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_2\, QN => 
        MASTER_SALT_POR_B_i_0_i_9);
    
    \U50_PATTERNS/U4C_REGCROSS/LOCAL_REG_VAL[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119105, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_21, Q => \ELKS_STRT_ADDR[7]\);
    
    HIEFFPLA_INST_0_52212 : MX2
      port map(A => HIEFFPLA_NET_0_161297, B => 
        HIEFFPLA_NET_0_161296, S => HIEFFPLA_NET_0_161295, Y => 
        HIEFFPLA_NET_0_117610);
    
    AFLSDF_INV_57 : INV
      port map(A => \U_DDR_ELK0/ELK0_IN_DDR_F\, Y => 
        \AFLSDF_INV_57\);
    
    \U50_PATTERNS/ELINK_DINA_12[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119841, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_12, Q => 
        \U50_PATTERNS/ELINK_DINA_12[6]\);
    
    HIEFFPLA_INST_0_44823 : NAND2B
      port map(A => HIEFFPLA_NET_0_119038, B => 
        HIEFFPLA_NET_0_119040, Y => HIEFFPLA_NET_0_119041);
    
    \U_ELK2_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL\ : DFN1C0
      port map(D => \U_ELK2_CH/ELK_IN_F_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL_net_1\);
    
    HIEFFPLA_INST_0_62631 : MX2
      port map(A => HIEFFPLA_NET_0_117096, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_9[0]\, S => 
        HIEFFPLA_NET_0_117183, Y => HIEFFPLA_NET_0_115965);
    
    HIEFFPLA_INST_0_53746 : AND2A
      port map(A => HIEFFPLA_NET_0_117391, B => 
        HIEFFPLA_NET_0_117392, Y => HIEFFPLA_NET_0_117360);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_4[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116329, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_20, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_4[0]\);
    
    HIEFFPLA_INST_0_60086 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_6[2]\, B => 
        HIEFFPLA_NET_0_116308, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_0[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116312);
    
    HIEFFPLA_INST_0_49694 : MX2
      port map(A => HIEFFPLA_NET_0_118095, B => 
        HIEFFPLA_NET_0_118092, S => \BIT_OS_SEL_6[1]\, Y => 
        HIEFFPLA_NET_0_118084);
    
    HIEFFPLA_INST_0_46401 : AO1
      port map(A => HIEFFPLA_NET_0_119276, B => 
        \U50_PATTERNS/ELINK_DOUTA_10[5]\, C => 
        HIEFFPLA_NET_0_118848, Y => HIEFFPLA_NET_0_118698);
    
    HIEFFPLA_INST_0_43982 : MX2
      port map(A => \U50_PATTERNS/TFC_STOP_ADDR[0]\, B => 
        \U50_PATTERNS/TFC_STOP_ADDR_T[0]\, S => 
        HIEFFPLA_NET_0_119472, Y => HIEFFPLA_NET_0_119188);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_22[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116448, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_15, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_22[2]\);
    
    HIEFFPLA_INST_0_45091 : MX2
      port map(A => HIEFFPLA_NET_0_118976, B => 
        \U50_PATTERNS/WR_USB_ADBUS[1]\, S => 
        HIEFFPLA_NET_0_119486, Y => HIEFFPLA_NET_0_118984);
    
    HIEFFPLA_INST_0_40792 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_16[6]\, B => 
        HIEFFPLA_NET_0_119566, S => HIEFFPLA_NET_0_119257, Y => 
        HIEFFPLA_NET_0_119809);
    
    HIEFFPLA_INST_0_37290 : AND2
      port map(A => \U200A_TFC/N_232_li\, B => 
        \U200A_TFC/GP_PG_SM[9]_net_1\, Y => HIEFFPLA_NET_0_120303);
    
    HIEFFPLA_INST_0_57067 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_2[6]\, B => 
        HIEFFPLA_NET_0_116729, S => HIEFFPLA_NET_0_117601, Y => 
        HIEFFPLA_NET_0_116749);
    
    HIEFFPLA_INST_0_45284 : AO1
      port map(A => HIEFFPLA_NET_0_119236, B => 
        \U50_PATTERNS/ELINK_DOUTA_0[7]\, C => 
        HIEFFPLA_NET_0_118838, Y => HIEFFPLA_NET_0_118951);
    
    HIEFFPLA_INST_0_59924 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_3[2]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_19[2]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_5[4]_net_1\, Y
         => HIEFFPLA_NET_0_116333);
    
    HIEFFPLA_INST_0_38071 : OR3B
      port map(A => \U200B_ELINKS/RX_SER_WORD_2DEL[3]_net_1\, B
         => \U200B_ELINKS/RX_SER_WORD_2DEL[2]_net_1\, C => 
        HIEFFPLA_NET_0_120159, Y => HIEFFPLA_NET_0_120160);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_23[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116119, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_6, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_23[1]\);
    
    HIEFFPLA_INST_0_54550 : MX2
      port map(A => HIEFFPLA_NET_0_117270, B => 
        HIEFFPLA_NET_0_117284, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[2]_net_1\, Y => 
        HIEFFPLA_NET_0_117250);
    
    HIEFFPLA_INST_0_62744 : AND2A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_SEQCNT[0]\, B => 
        HIEFFPLA_NET_0_116957, Y => HIEFFPLA_NET_0_115950);
    
    HIEFFPLA_INST_0_56909 : NAND3A
      port map(A => HIEFFPLA_NET_0_116777, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_1[7]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_1[6]\, Y => 
        HIEFFPLA_NET_0_116778);
    
    HIEFFPLA_INST_0_46690 : MX2
      port map(A => HIEFFPLA_NET_0_118628, B => 
        HIEFFPLA_NET_0_118624, S => \BIT_OS_SEL_5[1]\, Y => 
        HIEFFPLA_NET_0_118627);
    
    HIEFFPLA_INST_0_42975 : AO1
      port map(A => HIEFFPLA_NET_0_119014, B => 
        HIEFFPLA_NET_0_119377, C => HIEFFPLA_NET_0_119445, Y => 
        HIEFFPLA_NET_0_119412);
    
    \U_MASTER_DES/U13A_ADJ_160M/SSHIFT/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117615, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_13, Q => \U_MASTER_DES/AUX_SSHIFT\);
    
    HIEFFPLA_INST_0_37505 : NAND3B
      port map(A => \U200A_TFC/RX_SER_WORD_2DEL[0]_net_1\, B => 
        HIEFFPLA_NET_0_120271, C => 
        \U200A_TFC/RX_SER_WORD_2DEL[1]_net_1\, Y => 
        HIEFFPLA_NET_0_120272);
    
    \U_ELK1_CH/U_SLAVE_1ELK/RECD_SER_WORD[7]\ : DFN1C0
      port map(D => \U_ELK1_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[7]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_1[7]\);
    
    \U50_PATTERNS/TFC_DINA[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119191, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_4, Q => \U50_PATTERNS/TFC_DINA[6]\);
    
    HIEFFPLA_INST_0_52570 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_1[2]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_2[2]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[0]\, Y => 
        HIEFFPLA_NET_0_117546);
    
    HIEFFPLA_INST_0_46879 : NAND2B
      port map(A => \OP_MODE_c[1]\, B => \PATT_ELK_DAT_11[7]\, Y
         => HIEFFPLA_NET_0_118591);
    
    HIEFFPLA_INST_0_45212 : NAND3C
      port map(A => HIEFFPLA_NET_0_118743, B => 
        HIEFFPLA_NET_0_118752, C => HIEFFPLA_NET_0_118760, Y => 
        HIEFFPLA_NET_0_118964);
    
    AFLSDF_INV_63 : INV
      port map(A => \U_ELK1_CH/U_DDR_ELK1/ELK_IN_DDR_R\, Y => 
        \AFLSDF_INV_63\);
    
    \U50_PATTERNS/ELINK_DINA_12[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119847, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_12, Q => 
        \U50_PATTERNS/ELINK_DINA_12[0]\);
    
    HIEFFPLA_INST_0_43562 : NAND2B
      port map(A => \U50_PATTERNS/SM_BANK_SEL[21]\, B => 
        \U50_PATTERNS/SM_BANK_SEL[10]\, Y => 
        HIEFFPLA_NET_0_119292);
    
    HIEFFPLA_INST_0_38822 : MX2
      port map(A => HIEFFPLA_NET_0_119519, B => 
        \U50_PATTERNS/ELINK_ADDRA_13[4]\, S => 
        HIEFFPLA_NET_0_119285, Y => HIEFFPLA_NET_0_120059);
    
    \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[7]\ : DFN1C0
      port map(D => 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\);
    
    HIEFFPLA_INST_0_44339 : AND2
      port map(A => \U50_PATTERNS/U4B_REGCROSS/DELCNT[0]_net_1\, 
        B => \U50_PATTERNS/U4B_REGCROSS/DELCNT[1]_net_1\, Y => 
        HIEFFPLA_NET_0_119135);
    
    HIEFFPLA_INST_0_112187 : AO1A
      port map(A => HIEFFPLA_NET_0_120328, B => 
        HIEFFPLA_NET_0_115816, C => HIEFFPLA_NET_0_120323, Y => 
        HIEFFPLA_NET_0_120349);
    
    \U_ELK14_CH/U_SLAVE_1ELK/Q[0]\ : DFN1C0
      port map(D => \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/Q[0]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_9[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116283, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_6, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_9[2]\);
    
    \U_EXEC_MASTER/MPOR_B_32\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117787, CLK => CLK_40M_GL, CLR
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_0\, Q => 
        P_MASTER_POR_B_c_32);
    
    \U_ELK7_CH/U_SLAVE_1ELK/RECD_SER_WORD[2]\ : DFN1C0
      port map(D => \U_ELK7_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[2]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_7[2]\);
    
    HIEFFPLA_INST_0_55746 : MX2
      port map(A => HIEFFPLA_NET_0_116975, B => 
        HIEFFPLA_NET_0_117001, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[2]\, Y => 
        HIEFFPLA_NET_0_116995);
    
    \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[1]\ : DFN1C0
      port map(D => 
        \U_ELK14_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\);
    
    HIEFFPLA_INST_0_54956 : AND2A
      port map(A => HIEFFPLA_NET_0_117212, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_3[6]_net_1\, Y => 
        HIEFFPLA_NET_0_117157);
    
    HIEFFPLA_INST_0_47748 : MX2
      port map(A => HIEFFPLA_NET_0_118447, B => 
        HIEFFPLA_NET_0_118443, S => \BIT_OS_SEL_4[0]\, Y => 
        \U_ELK14_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[1]\);
    
    HIEFFPLA_INST_0_60441 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_11[0]\, B => 
        HIEFFPLA_NET_0_117096, S => HIEFFPLA_NET_0_117348, Y => 
        HIEFFPLA_NET_0_116265);
    
    HIEFFPLA_INST_0_46228 : AO1
      port map(A => HIEFFPLA_NET_0_119246, B => 
        \U50_PATTERNS/ELINK_DOUTA_3[5]\, C => 
        HIEFFPLA_NET_0_118908, Y => HIEFFPLA_NET_0_118737);
    
    \U_ELK3_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2\ : IOPADN_BI
      port map(DB => \U_ELK3_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, 
        E => \U_ELK3_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET3\, PAD => 
        ELK3_DAT_N, N2POUT => 
        \U_ELK3_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2_N2P\);
    
    \U_ELK16_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118376, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_10, Q => 
        \U_ELK16_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]_net_1\);
    
    \U_ELK12_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2\ : IOPADN_BI
      port map(DB => \U_ELK12_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, 
        E => \U_ELK12_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET3\, PAD
         => ELK12_DAT_N, N2POUT => 
        \U_ELK12_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2_N2P\);
    
    HIEFFPLA_INST_0_45358 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_18[6]\, C => 
        \U50_PATTERNS/SM_BANK_SEL[1]\, Y => HIEFFPLA_NET_0_118931);
    
    HIEFFPLA_INST_0_57095 : AND3
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_2[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_2[0]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_2[2]\, Y => 
        HIEFFPLA_NET_0_116746);
    
    HIEFFPLA_INST_0_50702 : MX2
      port map(A => \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\, B
         => \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[11]_net_1\, S => 
        \BIT_OS_SEL_4[2]\, Y => HIEFFPLA_NET_0_117903);
    
    HIEFFPLA_INST_0_45366 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_9[0]\, C => 
        \U50_PATTERNS/SM_BANK_SEL[10]\, Y => 
        HIEFFPLA_NET_0_118929);
    
    \U200B_ELINKS/ADDR_POINTER[5]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120250, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_32, Q => \ELKS_ADDRB[5]\);
    
    HIEFFPLA_INST_0_56428 : AND3
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[6]_net_1\, B => 
        HIEFFPLA_NET_0_117427, C => HIEFFPLA_NET_0_117423, Y => 
        HIEFFPLA_NET_0_116869);
    
    HIEFFPLA_INST_0_37507 : NAND3C
      port map(A => HIEFFPLA_NET_0_120274, B => 
        \U200A_TFC/RX_SER_WORD_2DEL[4]_net_1\, C => 
        \U200A_TFC/RX_SER_WORD_2DEL[5]_net_1\, Y => 
        HIEFFPLA_NET_0_120271);
    
    \U_ELK3_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U3\ : IOBI_ID_OD_EB
      port map(DR => \U_ELK3_CH/ELK_OUT_R_i_0\, DF => 
        \U_ELK3_CH/ELK_OUT_F_i_0\, CLR => \GND\, E => 
        \AFLSDF_INV_39\, ICLK => CCC_160M_ADJ, OCLK => 
        CCC_160M_FXD, YIN => 
        \U_ELK3_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\, DOUT => OPEN, 
        EOUT => \U_ELK3_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET3\, YR
         => OPEN, YF => OPEN);
    
    \U50_PATTERNS/OP_MODE[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119612, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_15, Q => \U50_PATTERNS/OP_MODE[5]\);
    
    HIEFFPLA_INST_0_45997 : AND3B
      port map(A => HIEFFPLA_NET_0_119426, B => 
        HIEFFPLA_NET_0_119379, C => \U50_PATTERNS/OP_MODE[1]\, Y
         => HIEFFPLA_NET_0_118793);
    
    HIEFFPLA_INST_0_45907 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_9[6]\, C => 
        \U50_PATTERNS/SM_BANK_SEL[10]\, Y => 
        HIEFFPLA_NET_0_118814);
    
    \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[0]\ : DFN1C0
      port map(D => 
        \U_ELK6_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\);
    
    HIEFFPLA_INST_0_47879 : MX2
      port map(A => \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[1]_net_1\, 
        B => \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\, S => 
        \BIT_OS_SEL_1[2]\, Y => HIEFFPLA_NET_0_118410);
    
    HIEFFPLA_INST_0_60884 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_17[2]\, B => 
        HIEFFPLA_NET_0_117181, S => HIEFFPLA_NET_0_117169, Y => 
        HIEFFPLA_NET_0_116203);
    
    HIEFFPLA_INST_0_52291 : AND3
      port map(A => HIEFFPLA_NET_0_117603, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[4]_net_1\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[5]_net_1\, Y => 
        HIEFFPLA_NET_0_117589);
    
    HIEFFPLA_INST_0_42921 : AND3A
      port map(A => \U50_PATTERNS/REG_STATE[5]_net_1\, B => 
        \U50_PATTERNS/REG_STATE[2]_net_1\, C => 
        \U50_PATTERNS/REG_STATE[3]_net_1\, Y => 
        HIEFFPLA_NET_0_119424);
    
    \U_ELK1_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0\ : DFN1C0
      port map(D => CLK_40M_GL, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_7, Q => 
        \U_ELK1_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_115939, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_24_0, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[2]_net_1\);
    
    \U50_PATTERNS/WR_USB_ADBUS[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118978, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_15, Q => 
        \U50_PATTERNS/WR_USB_ADBUS[7]\);
    
    HIEFFPLA_INST_0_111897 : XO1
      port map(A => \U50_PATTERNS/U4E_REGCROSS/SAMP_TWO[3]_net_1\, 
        B => \U50_PATTERNS/U4E_REGCROSS/LOCAL_REG_VAL[3]\, C => 
        HIEFFPLA_NET_0_115825, Y => HIEFFPLA_NET_0_119052);
    
    \U_ELK13_CH/U_SLAVE_1ELK/Q[12]\ : DFN1C0
      port map(D => \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/Q[12]_net_1\);
    
    \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_2S_11\ : DFN1C0
      port map(D => 
        \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_1S_net_1\, CLK
         => CLK60MHZ, CLR => \U_EXEC_MASTER/P_MASTER_POR_B_c_0\, 
        Q => P_USB_MASTER_EN_c_11);
    
    \U_ELK8_CH/U_ELK1_CMD_TX/START_RISE\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117879, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_12, Q => 
        \U_ELK8_CH/U_ELK1_CMD_TX/START_RISE_net_1\);
    
    HIEFFPLA_INST_0_58804 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_1[1]\, B => 
        HIEFFPLA_NET_0_116677, S => HIEFFPLA_NET_0_117158, Y => 
        HIEFFPLA_NET_0_116474);
    
    \U_ELK5_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118016, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_2, Q => 
        \U_ELK5_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]_net_1\);
    
    HIEFFPLA_INST_0_51829 : AOI1D
      port map(A => HIEFFPLA_NET_0_117684, B => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[2]\, C => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[3]\, Y => 
        HIEFFPLA_NET_0_117683);
    
    HIEFFPLA_INST_0_43559 : NAND2B
      port map(A => \U50_PATTERNS/SM_BANK_SEL_0[21]\, B => 
        \U50_PATTERNS/SM_BANK_SEL[7]\, Y => HIEFFPLA_NET_0_119295);
    
    \U_EXEC_MASTER/MPOR_SALT_B\ : DFI1P0
      port map(D => HIEFFPLA_NET_0_117781, CLK => CLK_40M_GL, PRE
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i\, QN => 
        MASTER_SALT_POR_B_i_0_i);
    
    \U_ELK14_CH/U_ELK1_SERDAT_SOURCE/SERDAT[5]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118458, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_6, Q => 
        \U_ELK14_CH/ELK_TX_DAT[5]\);
    
    HIEFFPLA_INST_0_55683 : MX2
      port map(A => HIEFFPLA_NET_0_115975, B => 
        HIEFFPLA_NET_0_116218, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_2[3]\, Y => 
        HIEFFPLA_NET_0_117004);
    
    HIEFFPLA_INST_0_39254 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_19[4]\, B => 
        HIEFFPLA_NET_0_119519, S => HIEFFPLA_NET_0_119293, Y => 
        HIEFFPLA_NET_0_120011);
    
    HIEFFPLA_INST_0_62263 : AND2A
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[0]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_31[0]\, Y
         => HIEFFPLA_NET_0_116015);
    
    AFLSDF_INV_30 : INV
      port map(A => DCB_SALT_SEL_c, Y => \AFLSDF_INV_30\);
    
    \U_ELK14_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]\ : DFN1C0
      port map(D => \U_ELK14_CH/U_SLAVE_1ELK/Q[12]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]_net_1\);
    
    \U200A_TFC/RX_SER_WORD_2DEL[6]\ : DFN1C0
      port map(D => \U200A_TFC/RX_SER_WORD_1DEL[6]_net_1\, CLK
         => CLK_40M_GL, CLR => P_MASTER_POR_B_c, Q => 
        \U200A_TFC/RX_SER_WORD_2DEL[6]_net_1\);
    
    \U_ELK2_CH/U_SLAVE_1ELK/RECD_SER_WORD[3]\ : DFN1C0
      port map(D => \U_ELK2_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[3]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_2[3]\);
    
    HIEFFPLA_INST_0_54149 : MX2
      port map(A => HIEFFPLA_NET_0_116175, B => 
        HIEFFPLA_NET_0_116064, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_1[3]_net_1\, Y
         => HIEFFPLA_NET_0_117302);
    
    HIEFFPLA_INST_0_55215 : NAND2A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[6]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[8]_net_1\, Y => 
        HIEFFPLA_NET_0_117086);
    
    \U_ELK11_CH/U_ELK1_SERDAT_SOURCE/SERDAT[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118595, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_0, Q => 
        \U_ELK11_CH/ELK_TX_DAT[3]\);
    
    HIEFFPLA_INST_0_55922 : MX2
      port map(A => HIEFFPLA_NET_0_117016, B => 
        HIEFFPLA_NET_0_117005, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[2]\, Y => 
        HIEFFPLA_NET_0_116973);
    
    \U_EXEC_MASTER/USB_MASTER_EN/T_CNT60M[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117743, CLK => CLK60MHZ, CLR
         => P_MASTER_POR_B_c_28, Q => 
        \U_EXEC_MASTER/USB_MASTER_EN/T_CNT60M[0]_net_1\);
    
    HIEFFPLA_INST_0_54815 : AO1B
      port map(A => HIEFFPLA_NET_0_117147, B => 
        HIEFFPLA_NET_0_117217, C => HIEFFPLA_NET_0_117086, Y => 
        HIEFFPLA_NET_0_117196);
    
    HIEFFPLA_INST_0_44793 : XOR2
      port map(A => \OP_MODE_c[6]\, B => 
        \U50_PATTERNS/U4E_REGCROSS/SAMP_TWO[6]_net_1\, Y => 
        HIEFFPLA_NET_0_119048);
    
    \U_ELK12_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]\ : DFN1C0
      port map(D => \U_ELK12_CH/U_SLAVE_1ELK/Q[9]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]_net_1\);
    
    \U_ELK19_CH/U_ELK1_SERDAT_SOURCE/SERDAT[5]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118233, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_15, Q => 
        \U_ELK19_CH/ELK_TX_DAT[5]\);
    
    HIEFFPLA_INST_0_50959 : MX2
      port map(A => \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\, B
         => \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[11]_net_1\, S => 
        \BIT_OS_SEL_3[2]\, Y => HIEFFPLA_NET_0_117857);
    
    HIEFFPLA_INST_0_41593 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_8[7]\, B => 
        HIEFFPLA_NET_0_119560, S => HIEFFPLA_NET_0_119291, Y => 
        HIEFFPLA_NET_0_119720);
    
    HIEFFPLA_INST_0_46630 : NAND2B
      port map(A => \OP_MODE_c_3[1]\, B => \PATT_ELK_DAT_10[7]\, 
        Y => HIEFFPLA_NET_0_118636);
    
    \U50_PATTERNS/ELINK_DINA_11[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119853, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_11, Q => 
        \U50_PATTERNS/ELINK_DINA_11[2]\);
    
    HIEFFPLA_INST_0_61928 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_27[2]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_28[2]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[0]\, Y => 
        HIEFFPLA_NET_0_116058);
    
    HIEFFPLA_INST_0_38759 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_12[5]\, B => 
        HIEFFPLA_NET_0_119518, S => HIEFFPLA_NET_0_119295, Y => 
        HIEFFPLA_NET_0_120066);
    
    AFLSDF_INV_66 : INV
      port map(A => \U_ELK3_CH/U_DDR_ELK1/ELK_IN_DDR_F\, Y => 
        \AFLSDF_INV_66\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_25[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116092, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_10, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_25[3]\);
    
    \U_ELK9_CH/U_ELK1_CMD_TX/SER_OUT_FI\ : DFN1C0
      port map(D => 
        \U_ELK9_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_12, Q
         => \U_ELK9_CH/U_ELK1_CMD_TX/SER_OUT_FI_net_1\);
    
    HIEFFPLA_INST_0_48180 : MX2
      port map(A => \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\, 
        B => \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[11]_net_1\, S => 
        \BIT_OS_SEL_1[2]\, Y => HIEFFPLA_NET_0_118357);
    
    HIEFFPLA_INST_0_45254 : AO1
      port map(A => HIEFFPLA_NET_0_119276, B => 
        \U50_PATTERNS/ELINK_DOUTA_10[1]\, C => 
        HIEFFPLA_NET_0_118844, Y => HIEFFPLA_NET_0_118957);
    
    HIEFFPLA_INST_0_51414 : AND3
      port map(A => HIEFFPLA_NET_0_117783, B => 
        \U_EXEC_MASTER/DEL_CNT[7]\, C => 
        \U_EXEC_MASTER/DEL_CNT[1]\, Y => HIEFFPLA_NET_0_117780);
    
    \U_ELK9_CH/U_ELK1_SERDAT_SOURCE/SERDAT[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117831, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_7, Q => 
        \U_ELK9_CH/ELK_TX_DAT[2]\);
    
    \U50_PATTERNS/U4E_REGCROSS/SAMP_ONE[6]\ : DFN1C0
      port map(D => \U50_PATTERNS/OP_MODE[6]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c, Q => 
        \U50_PATTERNS/U4E_REGCROSS/SAMP_ONE[6]_net_1\);
    
    HIEFFPLA_INST_0_45616 : NAND3C
      port map(A => HIEFFPLA_NET_0_118724, B => 
        HIEFFPLA_NET_0_118896, C => HIEFFPLA_NET_0_118714, Y => 
        HIEFFPLA_NET_0_118880);
    
    \U50_PATTERNS/ELINK_DINA_17[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119802, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_19, Q => 
        \U50_PATTERNS/ELINK_DINA_17[5]\);
    
    \U200B_ELINKS/LOC_STOP_ADDR[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120181, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_7, Q => 
        \U200B_ELINKS/LOC_STOP_ADDR[6]\);
    
    HIEFFPLA_INST_0_45310 : AO1
      port map(A => HIEFFPLA_NET_0_119277, B => 
        \U50_PATTERNS/ELINK_DOUTA_11[3]\, C => 
        HIEFFPLA_NET_0_118825, Y => HIEFFPLA_NET_0_118945);
    
    \U_ELK14_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U1\ : IOBI_ID_OD_EB
      port map(DR => \U_ELK14_CH/ELK_OUT_R\, DF => 
        \U_ELK14_CH/ELK_OUT_F\, CLR => \GND\, E => 
        \AFLSDF_INV_22\, ICLK => CCC_160M_ADJ, OCLK => 
        CCC_160M_FXD, YIN => 
        \U_ELK14_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\, DOUT => 
        \U_ELK14_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, EOUT => 
        \U_ELK14_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET2\, YR => 
        \U_ELK14_CH/ELK_IN_DDR_R\, YF => 
        \U_ELK14_CH/ELK_IN_DDR_F\);
    
    \U0B_TX40M_REFCLK/\\\\OUTBUF_LVDS[0]\\\\/U0/U0\ : IOPADP_TRI
      port map(D => 
        \U0B_TX40M_REFCLK/\\\\OUTBUF_LVDS[0]\\\\/U0/NET1\, E => 
        \U0B_TX40M_REFCLK/\\\\OUTBUF_LVDS[0]\\\\/U0/NET2\, PAD
         => TX_CLK40M_P);
    
    HIEFFPLA_INST_0_62039 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_29[2]\, B => 
        HIEFFPLA_NET_0_117131, S => HIEFFPLA_NET_0_117072, Y => 
        HIEFFPLA_NET_0_116043);
    
    HIEFFPLA_INST_0_53248 : AND2B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[8]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[0]\, Y => 
        HIEFFPLA_NET_0_117447);
    
    HIEFFPLA_INST_0_49212 : MX2
      port map(A => HIEFFPLA_NET_0_118182, B => 
        HIEFFPLA_NET_0_118180, S => \BIT_OS_SEL_0[1]\, Y => 
        HIEFFPLA_NET_0_118172);
    
    HIEFFPLA_INST_0_41981 : AND3C
      port map(A => HIEFFPLA_NET_0_119237, B => 
        HIEFFPLA_NET_0_119270, C => 
        \U50_PATTERNS/SM_BANK_SEL[14]\, Y => 
        HIEFFPLA_NET_0_119638);
    
    \U_ELK5_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]\ : DFN1C0
      port map(D => \U_ELK5_CH/U_SLAVE_1ELK/Q[1]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]_net_1\);
    
    \U_ELK2_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]\ : DFN1C0
      port map(D => \U_ELK2_CH/U_SLAVE_1ELK/Q[9]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]_net_1\);
    
    HIEFFPLA_INST_0_56871 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_1[5]\, B => 
        HIEFFPLA_NET_0_116762, S => HIEFFPLA_NET_0_117600, Y => 
        HIEFFPLA_NET_0_116783);
    
    HIEFFPLA_INST_0_48166 : MX2
      port map(A => HIEFFPLA_NET_0_118360, B => 
        HIEFFPLA_NET_0_118357, S => \BIT_OS_SEL_2[1]\, Y => 
        HIEFFPLA_NET_0_118359);
    
    HIEFFPLA_INST_0_41695 : MX2
      port map(A => HIEFFPLA_NET_0_119688, B => 
        \U50_PATTERNS/ELINK_RWA[12]\, S => 
        \U50_PATTERNS/SM_BANK_SEL_0[20]\, Y => 
        HIEFFPLA_NET_0_119708);
    
    HIEFFPLA_INST_0_46579 : NAND2B
      port map(A => \OP_MODE_c_4[1]\, B => \PATT_ELK_DAT_0[3]\, Y
         => HIEFFPLA_NET_0_118657);
    
    \U50_PATTERNS/ELINK_ADDRA_11[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120079, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_2, Q => 
        \U50_PATTERNS/ELINK_ADDRA_11[0]\);
    
    HIEFFPLA_INST_0_43955 : MX2
      port map(A => HIEFFPLA_NET_0_119566, B => 
        \U50_PATTERNS/TFC_DINA[6]\, S => HIEFFPLA_NET_0_119294, Y
         => HIEFFPLA_NET_0_119191);
    
    HIEFFPLA_INST_0_49905 : MX2
      port map(A => \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\, B
         => \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\, S => 
        \BIT_OS_SEL_6[2]\, Y => HIEFFPLA_NET_0_118045);
    
    HIEFFPLA_INST_0_37585 : AO1A
      port map(A => \ELKS_STRT_ADDR[0]\, B => 
        HIEFFPLA_NET_0_120219, C => HIEFFPLA_NET_0_120243, Y => 
        HIEFFPLA_NET_0_120254);
    
    HIEFFPLA_INST_0_56701 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_0[7]\, B => 
        HIEFFPLA_NET_0_116793, S => HIEFFPLA_NET_0_117602, Y => 
        HIEFFPLA_NET_0_116817);
    
    HIEFFPLA_INST_0_51872 : AX1
      port map(A => HIEFFPLA_NET_0_117682, B => 
        HIEFFPLA_NET_0_117686, C => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[5]\, Y => 
        HIEFFPLA_NET_0_117673);
    
    \P_MASTER_POR_B_pad/U0/U1\ : IOTRI_OB_EB
      port map(D => P_MASTER_POR_B_c, E => \VCC\, DOUT => 
        \P_MASTER_POR_B_pad/U0/NET1\, EOUT => 
        \P_MASTER_POR_B_pad/U0/NET2\);
    
    HIEFFPLA_INST_0_62316 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_3[4]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_4[4]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_4[0]\, Y => 
        HIEFFPLA_NET_0_116005);
    
    HIEFFPLA_INST_0_52872 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_19[3]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_20[3]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_1[0]\, Y => 
        HIEFFPLA_NET_0_117497);
    
    \U_ELK8_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]\ : DFN1C0
      port map(D => \U_ELK8_CH/U_SLAVE_1ELK/Q[14]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]_net_1\);
    
    HIEFFPLA_INST_0_55011 : AO1
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_3[6]_net_1\, B => 
        HIEFFPLA_NET_0_117203, C => HIEFFPLA_NET_0_117182, Y => 
        HIEFFPLA_NET_0_117141);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_27[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116069, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_13, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_27[1]\);
    
    \U50_PATTERNS/ELINK_BLKA[9]/U1\ : DFN1P0
      port map(D => HIEFFPLA_NET_0_119916, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_19, Q => 
        \U50_PATTERNS/ELINK_BLKA[9]\);
    
    HIEFFPLA_INST_0_48825 : AND2
      port map(A => \U_ELK19_CH/ELK_TX_DAT[0]\, B => 
        \U_ELK19_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118247);
    
    HIEFFPLA_INST_0_44078 : MX2
      port map(A => \U50_PATTERNS/TFC_STOP_ADDR_T[4]\, B => 
        \U50_PATTERNS/RD_USB_ADBUS[4]\, S => 
        HIEFFPLA_NET_0_119492, Y => HIEFFPLA_NET_0_119176);
    
    \U_ELK4_CH/U_SLAVE_1ELK/RECD_SER_WORD[7]\ : DFN1C0
      port map(D => \U_ELK4_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[7]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_4[7]\);
    
    \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[7]\ : DFN1C0
      port map(D => \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\);
    
    \U_ELK3_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL\ : DFN1C0
      port map(D => 
        \U_ELK3_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL_net_1\);
    
    \U50_PATTERNS/ELINKS_STOP_ADDR_T[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120113, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_7, Q => 
        \U50_PATTERNS/ELINKS_STOP_ADDR_T[6]\);
    
    HIEFFPLA_INST_0_45487 : AND3A
      port map(A => HIEFFPLA_NET_0_119437, B => 
        \U50_PATTERNS/WR_XFER_TYPE[1]_net_1\, C => 
        HIEFFPLA_NET_0_119367, Y => HIEFFPLA_NET_0_118904);
    
    \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[11]\ : DFN1C0
      port map(D => 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]_net_1\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[11]_net_1\);
    
    \U200A_TFC/LOC_STOP_ADDR[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120287, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_1, Q => \U200A_TFC/LOC_STOP_ADDR[3]\);
    
    HIEFFPLA_INST_0_38078 : NAND3C
      port map(A => \U200B_ELINKS/RX_SER_WORD_3DEL_i_0[3]\, B => 
        \U200B_ELINKS/RX_SER_WORD_3DEL_i_0[2]\, C => 
        HIEFFPLA_NET_0_120157, Y => HIEFFPLA_NET_0_120158);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_11[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116265, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_20, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_11[0]\);
    
    HIEFFPLA_INST_0_50319 : AND2
      port map(A => \U_ELK6_CH/ELK_TX_DAT[0]\, B => 
        \U_ELK6_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_117977);
    
    HIEFFPLA_INST_0_42109 : MX2
      port map(A => \U50_PATTERNS/OP_MODE[2]\, B => 
        \U50_PATTERNS/OP_MODE_T[2]\, S => HIEFFPLA_NET_0_119472, 
        Y => HIEFFPLA_NET_0_119615);
    
    \U50_PATTERNS/WR_XFER_TYPE[7]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118682, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c, Q => 
        \U50_PATTERNS/WR_XFER_TYPE[7]_net_1\);
    
    HIEFFPLA_INST_0_51441 : XA1A
      port map(A => HIEFFPLA_NET_0_117785, B => 
        \U_EXEC_MASTER/DEL_CNT[5]\, C => 
        \U_EXEC_MASTER/CCC_1_LOCK_STAT_1D_net_1\, Y => 
        HIEFFPLA_NET_0_117773);
    
    \U50_PATTERNS/ELINK_DINA_19[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119791, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_0, Q => 
        \U50_PATTERNS/ELINK_DINA_19[0]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_2[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116366, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_18, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_2[1]\);
    
    \U50_PATTERNS/U4E_REGCROSS/LOCAL_REG_VAL[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119068, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_6, Q => \OP_MODE_c[2]\);
    
    HIEFFPLA_INST_0_54847 : AND2B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_0[8]_net_1\, B => 
        HIEFFPLA_NET_0_117338, Y => HIEFFPLA_NET_0_117190);
    
    HIEFFPLA_INST_0_49642 : MX2
      port map(A => \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[3]_net_1\, B
         => \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\, S => 
        \BIT_OS_SEL_7[2]\, Y => HIEFFPLA_NET_0_118092);
    
    HIEFFPLA_INST_0_43670 : NAND2B
      port map(A => \U50_PATTERNS/SM_BANK_SEL_0[21]\, B => 
        \U50_PATTERNS/SM_BANK_SEL[16]\, Y => 
        HIEFFPLA_NET_0_119247);
    
    \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[14]\ : DFN1C0
      port map(D => 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[14]_net_1\);
    
    HIEFFPLA_INST_0_44748 : MX2
      port map(A => \OP_MODE_c_5[1]\, B => 
        \U50_PATTERNS/U4E_REGCROSS/SAMP_TWO[1]_net_1\, S => 
        HIEFFPLA_NET_0_119072, Y => HIEFFPLA_NET_0_119057);
    
    \U50_PATTERNS/ELINK_ADDRA_5[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119973, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_3, Q => 
        \U50_PATTERNS/ELINK_ADDRA_5[2]\);
    
    HIEFFPLA_INST_0_57740 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_6[4]\, B => 
        HIEFFPLA_NET_0_116611, S => HIEFFPLA_NET_0_117599, Y => 
        HIEFFPLA_NET_0_116628);
    
    HIEFFPLA_INST_0_42588 : AND3B
      port map(A => HIEFFPLA_NET_0_119452, B => 
        HIEFFPLA_NET_0_119499, C => HIEFFPLA_NET_0_119521, Y => 
        HIEFFPLA_NET_0_119505);
    
    \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[1]\ : DFN1C0
      port map(D => 
        \U_ELK15_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\);
    
    AFLSDF_INV_44 : INV
      port map(A => DCB_SALT_SEL_c, Y => \AFLSDF_INV_44\);
    
    \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[39]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117713, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_33, Q => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[39]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_16[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116512, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_16, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_16[0]\);
    
    HIEFFPLA_INST_0_38196 : MX2
      port map(A => \U50_PATTERNS/CHKSUM[5]\, B => 
        HIEFFPLA_NET_0_120130, S => HIEFFPLA_NET_0_119470, Y => 
        HIEFFPLA_NET_0_120138);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_30[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116356, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_18, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_30[0]\);
    
    \U_ELK10_CH/U_ELK1_CMD_TX/START_RISE\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118644, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_1, Q => 
        \U_ELK10_CH/U_ELK1_CMD_TX/START_RISE_net_1\);
    
    HIEFFPLA_INST_0_48573 : MX2
      port map(A => \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\, 
        B => \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[14]_net_1\, S => 
        \BIT_OS_SEL_2[2]\, Y => HIEFFPLA_NET_0_118293);
    
    HIEFFPLA_INST_0_40369 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_10[7]\, B => 
        HIEFFPLA_NET_0_119560, S => HIEFFPLA_NET_0_119239, Y => 
        HIEFFPLA_NET_0_119856);
    
    \U_MASTER_DES/U13C_MASTER_DESER/Q[1]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[1]_net_1\, CLK => 
        CCC_160M_FXD, CLR => P_MASTER_POR_B_c_34, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/Q[1]_net_1\);
    
    HIEFFPLA_INST_0_57439 : AND3
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_4[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_4[0]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_4[2]\, Y => 
        HIEFFPLA_NET_0_116683);
    
    HIEFFPLA_INST_0_44608 : MX2
      port map(A => \ELKS_STOP_ADDR[7]\, B => 
        \U50_PATTERNS/U4D_REGCROSS/SAMP_TWO[7]_net_1\, S => 
        HIEFFPLA_NET_0_119093, Y => HIEFFPLA_NET_0_119084);
    
    \U_ELK8_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL\ : DFN1C0
      port map(D => \U_ELK8_CH/ELK_IN_F_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/BEST_BIT_OS_VAL[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_117579, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_14, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_BIT_OS_VAL[1]\);
    
    HIEFFPLA_INST_0_59325 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_26[0]\, B => 
        HIEFFPLA_NET_0_116402, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_2[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116406);
    
    HIEFFPLA_INST_0_42853 : AND3B
      port map(A => HIEFFPLA_NET_0_119451, B => 
        \U50_PATTERNS/REG_STATE[0]_net_1\, C => 
        HIEFFPLA_NET_0_119429, Y => HIEFFPLA_NET_0_119447);
    
    \U_ELK13_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U0\ : IOPADP_BI
      port map(N2PIN => 
        \U_ELK13_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2_N2P\, D => 
        \U_ELK13_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, E => 
        \U_ELK13_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET2\, PAD => 
        ELK13_DAT_P, Y => 
        \U_ELK13_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\);
    
    HIEFFPLA_INST_0_52361 : AND2A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[8]_net_1\, B => 
        HIEFFPLA_NET_0_117571, Y => HIEFFPLA_NET_0_117575);
    
    HIEFFPLA_INST_0_60747 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_15[4]\, B => 
        HIEFFPLA_NET_0_117166, S => HIEFFPLA_NET_0_117356, Y => 
        HIEFFPLA_NET_0_116226);
    
    HIEFFPLA_INST_0_38921 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_14[7]\, B => 
        HIEFFPLA_NET_0_119516, S => HIEFFPLA_NET_0_119249, Y => 
        HIEFFPLA_NET_0_120048);
    
    \U_ELK13_CH/U_ELK1_CMD_TX/SER_OUT_FI\ : DFN1C0
      port map(D => 
        \U_ELK13_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_1, Q => 
        \U_ELK13_CH/U_ELK1_CMD_TX/SER_OUT_FI_net_1\);
    
    HIEFFPLA_INST_0_52073 : MX2
      port map(A => HIEFFPLA_NET_0_117633, B => 
        HIEFFPLA_NET_0_117632, S => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[4]\, Y => 
        HIEFFPLA_NET_0_117641);
    
    HIEFFPLA_INST_0_49662 : MX2
      port map(A => \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\, B
         => \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\, S => 
        \BIT_OS_SEL_7[2]\, Y => HIEFFPLA_NET_0_118089);
    
    HIEFFPLA_INST_0_111333 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_25[1]\, B => 
        HIEFFPLA_NET_0_116677, S => HIEFFPLA_NET_0_117394, Y => 
        HIEFFPLA_NET_0_116415);
    
    \U_ELK14_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]\ : DFN1C0
      port map(D => \U_ELK14_CH/U_SLAVE_1ELK/Q[14]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]_net_1\);
    
    HIEFFPLA_INST_0_52067 : MX2C
      port map(A => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[8]_net_1\, B => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[9]_net_1\, S => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[0]\, Y => 
        HIEFFPLA_NET_0_117642);
    
    HIEFFPLA_INST_0_43595 : NAND2B
      port map(A => \U50_PATTERNS/SM_BANK_SEL[21]\, B => 
        \U50_PATTERNS/SM_BANK_SEL[19]\, Y => 
        HIEFFPLA_NET_0_119272);
    
    HIEFFPLA_INST_0_37769 : AO1
      port map(A => HIEFFPLA_NET_0_120222, B => 
        HIEFFPLA_NET_0_120202, C => HIEFFPLA_NET_0_120194, Y => 
        HIEFFPLA_NET_0_120212);
    
    \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[8]\ : DFN1C0
      port map(D => 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\);
    
    HIEFFPLA_INST_0_44857 : NAND3C
      port map(A => HIEFFPLA_NET_0_119023, B => 
        HIEFFPLA_NET_0_119029, C => HIEFFPLA_NET_0_119028, Y => 
        HIEFFPLA_NET_0_119034);
    
    \U_ELK13_CH/U_SLAVE_1ELK/Q[5]\ : DFN1C0
      port map(D => \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/Q[5]_net_1\);
    
    HIEFFPLA_INST_0_52206 : MX2
      port map(A => HIEFFPLA_NET_0_161294, B => 
        HIEFFPLA_NET_0_161293, S => HIEFFPLA_NET_0_161292, Y => 
        HIEFFPLA_NET_0_117611);
    
    HIEFFPLA_INST_0_50953 : MX2
      port map(A => \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\, B
         => \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\, S => 
        \BIT_OS_SEL_3[2]\, Y => HIEFFPLA_NET_0_117858);
    
    \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[0]\ : DFN1C0
      port map(D => 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[0]_net_1\);
    
    HIEFFPLA_INST_0_41877 : AOI1C
      port map(A => \U50_PATTERNS/ELINK_RWA[3]\, B => 
        HIEFFPLA_NET_0_119645, C => HIEFFPLA_NET_0_119676, Y => 
        HIEFFPLA_NET_0_119677);
    
    HIEFFPLA_INST_0_40176 : AOI1D
      port map(A => HIEFFPLA_NET_0_119389, B => 
        HIEFFPLA_NET_0_119464, C => 
        \U50_PATTERNS/SM_BANK_SEL[10]\, Y => 
        HIEFFPLA_NET_0_119879);
    
    \U_ELK12_CH/U_SLAVE_1ELK/RECD_SER_WORD[6]\ : DFN1C0
      port map(D => \U_ELK12_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[6]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_12[6]\);
    
    HIEFFPLA_INST_0_46279 : AO1
      port map(A => HIEFFPLA_NET_0_119476, B => 
        \U50_PATTERNS/CHKSUM[7]\, C => HIEFFPLA_NET_0_118898, Y
         => HIEFFPLA_NET_0_118726);
    
    HIEFFPLA_INST_0_44236 : AND2A
      port map(A => \U50_PATTERNS/U4A_REGCROSS/DELCNT[0]_net_1\, 
        B => \U50_PATTERNS/U4A_REGCROSS/SYNC_SM[0]_net_1\, Y => 
        HIEFFPLA_NET_0_119155);
    
    HIEFFPLA_INST_0_60146 : AOI1C
      port map(A => HIEFFPLA_NET_0_116675, B => 
        HIEFFPLA_NET_0_116589, C => HIEFFPLA_NET_0_117211, Y => 
        HIEFFPLA_NET_0_116304);
    
    HIEFFPLA_INST_0_42877 : NAND2B
      port map(A => HIEFFPLA_NET_0_119452, B => 
        HIEFFPLA_NET_0_119443, Y => HIEFFPLA_NET_0_119439);
    
    HIEFFPLA_INST_0_46106 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_12[2]\, C => 
        \U50_PATTERNS/SM_BANK_SEL[7]\, Y => HIEFFPLA_NET_0_118764);
    
    \U_ELK4_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]\ : DFN1C0
      port map(D => \U_ELK4_CH/U_SLAVE_1ELK/Q[13]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_8[4]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_115966, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_19, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_8[4]\);
    
    \U_ELK7_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117928, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_10, Q => 
        \U_ELK7_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]_net_1\);
    
    \U_ELK3_CH/U_SLAVE_1ELK/RECD_SER_WORD[7]\ : DFN1C0
      port map(D => \U_ELK3_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[7]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_3[7]\);
    
    HIEFFPLA_INST_0_49616 : AND2A
      port map(A => \OP_MODE_c_5[1]\, B => \PATT_ELK_DAT_3[5]\, Y
         => HIEFFPLA_NET_0_118098);
    
    HIEFFPLA_INST_0_57570 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_5[4]\, B => 
        HIEFFPLA_NET_0_116640, S => HIEFFPLA_NET_0_117121, Y => 
        HIEFFPLA_NET_0_116657);
    
    \U50_PATTERNS/ELINK_ADDRA_7[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119958, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_5, Q => 
        \U50_PATTERNS/ELINK_ADDRA_7[1]\);
    
    HIEFFPLA_INST_0_61364 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_21[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_22[1]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_3[0]\, Y => 
        HIEFFPLA_NET_0_116137);
    
    HIEFFPLA_INST_0_55069 : AND3A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[3]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[6]_net_1\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[7]_net_1\, Y => 
        HIEFFPLA_NET_0_117128);
    
    HIEFFPLA_INST_0_47049 : MX2
      port map(A => HIEFFPLA_NET_0_118580, B => 
        HIEFFPLA_NET_0_118565, S => \BIT_OS_SEL[0]\, Y => 
        \U_ELK11_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[7]\);
    
    HIEFFPLA_INST_0_61148 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_1[3]\, 
        B => HIEFFPLA_NET_0_117186, S => HIEFFPLA_NET_0_117149, Y
         => HIEFFPLA_NET_0_116167);
    
    HIEFFPLA_INST_0_43709 : NAND3C
      port map(A => HIEFFPLA_NET_0_119242, B => 
        HIEFFPLA_NET_0_119259, C => HIEFFPLA_NET_0_119261, Y => 
        HIEFFPLA_NET_0_119235);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_9[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_115965, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_20, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_9[0]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/BEST_SEQCNT[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117441, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_8, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_SEQCNT[1]\);
    
    HIEFFPLA_INST_0_46207 : AO1A
      port map(A => HIEFFPLA_NET_0_118921, B => 
        \U50_PATTERNS/SM_BANK_SEL[0]\, C => HIEFFPLA_NET_0_118742, 
        Y => HIEFFPLA_NET_0_118743);
    
    \U_ELK7_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]\ : DFN1C0
      port map(D => \U_ELK7_CH/U_SLAVE_1ELK/Q[9]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]_net_1\);
    
    HIEFFPLA_INST_0_59047 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_23[0]\, B => 
        HIEFFPLA_NET_0_116680, S => HIEFFPLA_NET_0_116438, Y => 
        HIEFFPLA_NET_0_116442);
    
    HIEFFPLA_INST_0_57111 : AO1A
      port map(A => HIEFFPLA_NET_0_116745, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_2[3]\, C => 
        HIEFFPLA_NET_0_116739, Y => HIEFFPLA_NET_0_116740);
    
    HIEFFPLA_INST_0_43006 : NAND3B
      port map(A => \U50_PATTERNS/REG_STATE[1]_net_1\, B => 
        \U50_PATTERNS/USB_RXF_B\, C => HIEFFPLA_NET_0_119429, Y
         => HIEFFPLA_NET_0_119405);
    
    HIEFFPLA_INST_0_43601 : NAND3C
      port map(A => HIEFFPLA_NET_0_119274, B => 
        HIEFFPLA_NET_0_119281, C => HIEFFPLA_NET_0_119273, Y => 
        HIEFFPLA_NET_0_119271);
    
    HIEFFPLA_INST_0_40333 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_10[3]\, B => 
        HIEFFPLA_NET_0_119574, S => HIEFFPLA_NET_0_119239, Y => 
        HIEFFPLA_NET_0_119860);
    
    HIEFFPLA_INST_0_38966 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_15[4]\, B => 
        HIEFFPLA_NET_0_119519, S => HIEFFPLA_NET_0_119297, Y => 
        HIEFFPLA_NET_0_120043);
    
    \U50_PATTERNS/U108_PATT_ELINK_BLK/DPRT_512X9_SRAM_R0C0\ : 
        RAM4K9
      generic map(MEMORYFILE => "DPRT_512X9_SRAM_R0C0.mem")

      port map(ADDRA11 => AFLSDF_GND, ADDRA10 => AFLSDF_GND, 
        ADDRA9 => AFLSDF_GND, ADDRA8 => \GND\, ADDRA7 => 
        \U50_PATTERNS/ELINK_ADDRA_8[7]\, ADDRA6 => 
        \U50_PATTERNS/ELINK_ADDRA_8[6]\, ADDRA5 => 
        \U50_PATTERNS/ELINK_ADDRA_8[5]\, ADDRA4 => 
        \U50_PATTERNS/ELINK_ADDRA_8[4]\, ADDRA3 => 
        \U50_PATTERNS/ELINK_ADDRA_8[3]\, ADDRA2 => 
        \U50_PATTERNS/ELINK_ADDRA_8[2]\, ADDRA1 => 
        \U50_PATTERNS/ELINK_ADDRA_8[1]\, ADDRA0 => 
        \U50_PATTERNS/ELINK_ADDRA_8[0]\, ADDRB11 => AFLSDF_GND, 
        ADDRB10 => AFLSDF_GND, ADDRB9 => AFLSDF_GND, ADDRB8 => 
        \GND\, ADDRB7 => \ELKS_ADDRB[7]\, ADDRB6 => 
        \ELKS_ADDRB_0[6]\, ADDRB5 => \ELKS_ADDRB[5]\, ADDRB4 => 
        \ELKS_ADDRB_0[4]\, ADDRB3 => \ELKS_ADDRB[3]\, ADDRB2 => 
        \ELKS_ADDRB_0[2]\, ADDRB1 => \ELKS_ADDRB[1]\, ADDRB0 => 
        \ELKS_ADDRB[0]\, DINA8 => \GND\, DINA7 => 
        \U50_PATTERNS/ELINK_DINA_8[7]\, DINA6 => 
        \U50_PATTERNS/ELINK_DINA_8[6]\, DINA5 => 
        \U50_PATTERNS/ELINK_DINA_8[5]\, DINA4 => 
        \U50_PATTERNS/ELINK_DINA_8[4]\, DINA3 => 
        \U50_PATTERNS/ELINK_DINA_8[3]\, DINA2 => 
        \U50_PATTERNS/ELINK_DINA_8[2]\, DINA1 => 
        \U50_PATTERNS/ELINK_DINA_8[1]\, DINA0 => 
        \U50_PATTERNS/ELINK_DINA_8[0]\, DINB8 => \GND\, DINB7 => 
        \ELK_RX_SER_WORD_8[7]\, DINB6 => \ELK_RX_SER_WORD_8[6]\, 
        DINB5 => \ELK_RX_SER_WORD_8[5]\, DINB4 => 
        \ELK_RX_SER_WORD_8[4]\, DINB3 => \ELK_RX_SER_WORD_8[3]\, 
        DINB2 => \ELK_RX_SER_WORD_8[2]\, DINB1 => 
        \ELK_RX_SER_WORD_8[1]\, DINB0 => \ELK_RX_SER_WORD_8[0]\, 
        WIDTHA0 => \VCC\, WIDTHA1 => \VCC\, WIDTHB0 => \VCC\, 
        WIDTHB1 => \VCC\, PIPEA => \VCC\, PIPEB => \VCC\, WMODEA
         => \GND\, WMODEB => \GND\, BLKA => 
        \U50_PATTERNS/ELINK_BLKA[8]\, BLKB => ELKS_RAM_BLKB_EN, 
        WENA => \U50_PATTERNS/ELINK_RWA[8]\, WENB => ELKS_RWB, 
        CLKA => CLK60MHZ, CLKB => CLK_40M_GL, RESET => 
        P_USB_MASTER_EN_c_0, DOUTA8 => OPEN, DOUTA7 => 
        \U50_PATTERNS/ELINK_DOUTA_8[7]\, DOUTA6 => 
        \U50_PATTERNS/ELINK_DOUTA_8[6]\, DOUTA5 => 
        \U50_PATTERNS/ELINK_DOUTA_8[5]\, DOUTA4 => 
        \U50_PATTERNS/ELINK_DOUTA_8[4]\, DOUTA3 => 
        \U50_PATTERNS/ELINK_DOUTA_8[3]\, DOUTA2 => 
        \U50_PATTERNS/ELINK_DOUTA_8[2]\, DOUTA1 => 
        \U50_PATTERNS/ELINK_DOUTA_8[1]\, DOUTA0 => 
        \U50_PATTERNS/ELINK_DOUTA_8[0]\, DOUTB8 => OPEN, DOUTB7
         => \PATT_ELK_DAT_8[7]\, DOUTB6 => \PATT_ELK_DAT_8[6]\, 
        DOUTB5 => \PATT_ELK_DAT_8[5]\, DOUTB4 => 
        \PATT_ELK_DAT_8[4]\, DOUTB3 => \PATT_ELK_DAT_8[3]\, 
        DOUTB2 => \PATT_ELK_DAT_8[2]\, DOUTB1 => 
        \PATT_ELK_DAT_8[1]\, DOUTB0 => \PATT_ELK_DAT_8[0]\);
    
    HIEFFPLA_INST_0_55144 : AO1
      port map(A => HIEFFPLA_NET_0_117128, B => 
        HIEFFPLA_NET_0_117584, C => HIEFFPLA_NET_0_117085, Y => 
        HIEFFPLA_NET_0_117113);
    
    HIEFFPLA_INST_0_41924 : NAND2B
      port map(A => \U50_PATTERNS/ELINK_RWA[12]\, B => 
        HIEFFPLA_NET_0_119659, Y => HIEFFPLA_NET_0_119660);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_25[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116095, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_10, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_25[0]\);
    
    HIEFFPLA_INST_0_43937 : MX2
      port map(A => HIEFFPLA_NET_0_119570, B => 
        \U50_PATTERNS/TFC_DINA[4]\, S => HIEFFPLA_NET_0_119294, Y
         => HIEFFPLA_NET_0_119193);
    
    HIEFFPLA_INST_0_57976 : AO1
      port map(A => HIEFFPLA_NET_0_116620, B => 
        HIEFFPLA_NET_0_116649, C => HIEFFPLA_NET_0_116589, Y => 
        HIEFFPLA_NET_0_116586);
    
    HIEFFPLA_INST_0_43167 : AND3A
      port map(A => HIEFFPLA_NET_0_119477, B => 
        HIEFFPLA_NET_0_119393, C => 
        \U50_PATTERNS/REG_STATE_0[5]_net_1\, Y => 
        HIEFFPLA_NET_0_119356);
    
    \U50_PATTERNS/U4B_REGCROSS/LOCAL_REG_VAL[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119127, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_19, Q => \TFC_STOP_ADDR[6]\);
    
    HIEFFPLA_INST_0_56243 : AND2A
      port map(A => DCB_SALT_SEL_c, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/RECD_SER_WORD[4]_net_1\, 
        Y => \TFC_RX_SER_WORD[4]\);
    
    HIEFFPLA_INST_0_63047 : AND3
      port map(A => HIEFFPLA_NET_0_115903, B => 
        HIEFFPLA_NET_0_115899, C => HIEFFPLA_NET_0_115901, Y => 
        HIEFFPLA_NET_0_115904);
    
    \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[5]\ : DFN1C0
      port map(D => 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\);
    
    HIEFFPLA_INST_0_54528 : NAND2
      port map(A => HIEFFPLA_NET_0_117208, B => 
        HIEFFPLA_NET_0_116678, Y => HIEFFPLA_NET_0_117254);
    
    HIEFFPLA_INST_0_47328 : MX2
      port map(A => \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\, 
        B => \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[14]_net_1\, S => 
        \BIT_OS_SEL_6[2]\, Y => HIEFFPLA_NET_0_118518);
    
    \U_ELK17_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]\ : DFN1C0
      port map(D => \U_ELK17_CH/U_SLAVE_1ELK/Q[5]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]_net_1\);
    
    \U_ELK17_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]\ : DFN1C0
      port map(D => \U_ELK17_CH/U_SLAVE_1ELK/Q[13]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]_net_1\);
    
    HIEFFPLA_INST_0_59558 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_29[0]\, B => 
        HIEFFPLA_NET_0_116680, S => HIEFFPLA_NET_0_117129, Y => 
        HIEFFPLA_NET_0_116378);
    
    HIEFFPLA_INST_0_62520 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_7[1]\, 
        B => HIEFFPLA_NET_0_117114, S => HIEFFPLA_NET_0_117174, Y
         => HIEFFPLA_NET_0_115979);
    
    \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[3]\ : DFN1C0
      port map(D => 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[3]_net_1\);
    
    \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[13]\ : DFN1C0
      port map(D => \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\, 
        CLK => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[13]_net_1\);
    
    HIEFFPLA_INST_0_63040 : NOR3A
      port map(A => HIEFFPLA_NET_0_115913, B => 
        HIEFFPLA_NET_0_115907, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[7]\, Y => 
        HIEFFPLA_NET_0_115906);
    
    HIEFFPLA_INST_0_55596 : MX2
      port map(A => HIEFFPLA_NET_0_116161, B => 
        HIEFFPLA_NET_0_116266, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_1[3]\, Y => 
        HIEFFPLA_NET_0_117016);
    
    \U_ELK12_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118560, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_15, Q => 
        \U_ELK12_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]_net_1\);
    
    HIEFFPLA_INST_0_42189 : MX2
      port map(A => \U50_PATTERNS/OP_MODE_T[4]\, B => 
        \U50_PATTERNS/RD_USB_ADBUS[4]\, S => 
        HIEFFPLA_NET_0_119440, Y => HIEFFPLA_NET_0_119605);
    
    AFLSDF_INV_18 : INV
      port map(A => DCB_SALT_SEL_c, Y => \AFLSDF_INV_18\);
    
    \U_ELK7_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117929, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_14, Q => 
        \U_ELK7_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]_net_1\);
    
    HIEFFPLA_INST_0_53336 : AND2B
      port map(A => \BIT_OS_SEL[2]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_SEL[3]_net_1\, Y
         => HIEFFPLA_NET_0_117423);
    
    \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[8]\ : DFN1C0
      port map(D => 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\);
    
    \U_ELK3_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]\ : DFN1C0
      port map(D => \U_ELK3_CH/U_SLAVE_1ELK/Q[2]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]_net_1\);
    
    \U_ELK19_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118243, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_4, Q => 
        \U_ELK19_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]_net_1\);
    
    HIEFFPLA_INST_0_38156 : MX2
      port map(A => \U50_PATTERNS/CHKSUM[1]\, B => 
        HIEFFPLA_NET_0_120134, S => HIEFFPLA_NET_0_119470, Y => 
        HIEFFPLA_NET_0_120142);
    
    \U_ELK14_CH/U_ELK1_SERDAT_SOURCE/SERDAT[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118462, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_6, Q => 
        \U_ELK14_CH/ELK_TX_DAT[1]\);
    
    HIEFFPLA_INST_0_41359 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_5[5]\, B => 
        HIEFFPLA_NET_0_119567, S => HIEFFPLA_NET_0_119251, Y => 
        HIEFFPLA_NET_0_119746);
    
    \U_ELK7_CH/U_SLAVE_1ELK/Q[3]\ : DFN1C0
      port map(D => \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/Q[3]_net_1\);
    
    \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[4]\ : DFN1C0
      port map(D => 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\);
    
    HIEFFPLA_INST_0_62810 : AOI1D
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[8]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[0]_net_1\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/TUNE_CLKPHASE[2]\, Y => 
        HIEFFPLA_NET_0_115944);
    
    \U_ELK1_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]\ : DFN1C0
      port map(D => \U_ELK1_CH/U_SLAVE_1ELK/Q[8]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]_net_1\);
    
    HIEFFPLA_INST_0_62364 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_4[2]\, 
        B => HIEFFPLA_NET_0_117131, S => HIEFFPLA_NET_0_117148, Y
         => HIEFFPLA_NET_0_115998);
    
    \U_EXEC_MASTER/MPOR_B_32_0\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117787, CLK => CLK_40M_GL, CLR
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_0\, Q => 
        P_MASTER_POR_B_c_32_0);
    
    \U_ELK2_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118151, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_8, Q => 
        \U_ELK2_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]_net_1\);
    
    HIEFFPLA_INST_0_47961 : MX2
      port map(A => \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\, 
        B => \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[12]_net_1\, S => 
        \BIT_OS_SEL_2[2]\, Y => HIEFFPLA_NET_0_118398);
    
    \U_ELK1_CH/U_ELK1_SERDAT_SOURCE/SERDAT[6]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118187, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_11, Q => 
        \U_ELK1_CH/ELK_TX_DAT[6]\);
    
    \P_OP_MODE6_EE_pad/U0/U1\ : IOTRI_OB_EB
      port map(D => \OP_MODE_c[6]\, E => \VCC\, DOUT => 
        \P_OP_MODE6_EE_pad/U0/NET1\, EOUT => 
        \P_OP_MODE6_EE_pad/U0/NET2\);
    
    HIEFFPLA_INST_0_50985 : MX2
      port map(A => HIEFFPLA_NET_0_117870, B => 
        HIEFFPLA_NET_0_117868, S => \BIT_OS_SEL_5[0]\, Y => 
        \U_ELK8_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[1]\);
    
    \U_ELK18_CH/U_SLAVE_1ELK/Q[2]\ : DFN1C0
      port map(D => \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/Q[2]_net_1\);
    
    HIEFFPLA_INST_0_61028 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_2[3]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_18[3]\, S
         => \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_4[4]_net_1\, 
        Y => HIEFFPLA_NET_0_116183);
    
    \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[8]\ : DFN1C0
      port map(D => \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_11[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116554, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_8, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_11[0]\);
    
    HIEFFPLA_INST_0_62015 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_12[4]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_28[4]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_3[4]_net_1\, Y
         => HIEFFPLA_NET_0_116046);
    
    HIEFFPLA_INST_0_58405 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_14[2]\, B => 
        HIEFFPLA_NET_0_116522, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_1[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116526);
    
    HIEFFPLA_INST_0_54464 : MX2
      port map(A => HIEFFPLA_NET_0_116471, B => 
        HIEFFPLA_NET_0_116281, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[3]_net_1\, Y => 
        HIEFFPLA_NET_0_117262);
    
    HIEFFPLA_INST_0_42309 : AND2A
      port map(A => HIEFFPLA_NET_0_119275, B => 
        \U50_PATTERNS/RD_USB_ADBUS[1]\, Y => 
        HIEFFPLA_NET_0_119576);
    
    \U_ELK19_CH/U_ELK1_SERDAT_SOURCE/SERDAT[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118237, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_15, Q => 
        \U_ELK19_CH/ELK_TX_DAT[1]\);
    
    HIEFFPLA_INST_0_57898 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_7[3]\, B => 
        HIEFFPLA_NET_0_116581, S => HIEFFPLA_NET_0_117113, Y => 
        HIEFFPLA_NET_0_116600);
    
    HIEFFPLA_INST_0_49113 : AND2A
      port map(A => \OP_MODE_c_5[1]\, B => \PATT_ELK_DAT_1[0]\, Y
         => HIEFFPLA_NET_0_118193);
    
    HIEFFPLA_INST_0_40156 : AOI1D
      port map(A => HIEFFPLA_NET_0_119389, B => 
        HIEFFPLA_NET_0_119464, C => 
        \U50_PATTERNS/SM_BANK_SEL[14]\, Y => 
        HIEFFPLA_NET_0_119887);
    
    \U50_PATTERNS/SM_BANK_SEL_0[20]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119300, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_1_0, Q => 
        \U50_PATTERNS/SM_BANK_SEL_0[20]\);
    
    \U50_PATTERNS/ELINK_DINA_0[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119865, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_5, Q => 
        \U50_PATTERNS/ELINK_DINA_0[6]\);
    
    \U50_PATTERNS/ELINK_ADDRA_12[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120066, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_2_0, Q => 
        \U50_PATTERNS/ELINK_ADDRA_12[5]\);
    
    HIEFFPLA_INST_0_49859 : AND2
      port map(A => CLK_40M_GL, B => 
        \U_ELK4_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0_net_1\, Y => 
        HIEFFPLA_NET_0_118059);
    
    HIEFFPLA_INST_0_43721 : AND2B
      port map(A => HIEFFPLA_NET_0_119262, B => 
        HIEFFPLA_NET_0_119270, Y => HIEFFPLA_NET_0_119232);
    
    HIEFFPLA_INST_0_50587 : AND2
      port map(A => \U_ELK7_CH/ELK_TX_DAT[1]\, B => 
        \U_ELK7_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_117928);
    
    HIEFFPLA_INST_0_51107 : NAND2B
      port map(A => \OP_MODE_c_3[1]\, B => \PATT_ELK_DAT_9[2]\, Y
         => HIEFFPLA_NET_0_117831);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_14[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116232, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_2, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_14[3]\);
    
    HIEFFPLA_INST_0_59912 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_3[0]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_19[0]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_4[4]_net_1\, Y
         => HIEFFPLA_NET_0_116335);
    
    HIEFFPLA_INST_0_51879 : AX1C
      port map(A => \U_MASTER_DES/U13A_ADJ_160M/BITCNT[6]\, B => 
        HIEFFPLA_NET_0_117690, C => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[7]\, Y => 
        HIEFFPLA_NET_0_117672);
    
    HIEFFPLA_INST_0_40585 : MX2
      port map(A => HIEFFPLA_NET_0_119560, B => 
        \U50_PATTERNS/ELINK_DINA_13[7]\, S => 
        HIEFFPLA_NET_0_119285, Y => HIEFFPLA_NET_0_119832);
    
    \U_ELK5_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118018, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_2, Q => 
        \U_ELK5_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]_net_1\);
    
    HIEFFPLA_INST_0_52201 : AND3A
      port map(A => \U_MASTER_DES/U13A_ADJ_160M/BITCNT[3]\, B => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[1]\, C => 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM[0]_net_1\, Y => 
        HIEFFPLA_NET_0_117612);
    
    \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117061, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_26, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[0]_net_1\);
    
    HIEFFPLA_INST_0_58622 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_1[3]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_17[3]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[4]_net_1\, Y
         => HIEFFPLA_NET_0_116497);
    
    HIEFFPLA_INST_0_56591 : AND3
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[7]_net_1\, B => 
        HIEFFPLA_NET_0_117424, C => HIEFFPLA_NET_0_117427, Y => 
        HIEFFPLA_NET_0_116832);
    
    HIEFFPLA_INST_0_56355 : AO1
      port map(A => HIEFFPLA_NET_0_117431, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[3]_net_1\, C => 
        HIEFFPLA_NET_0_116863, Y => HIEFFPLA_NET_0_116887);
    
    HIEFFPLA_INST_0_58169 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_10[3]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_26[3]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_2[4]_net_1\, Y
         => HIEFFPLA_NET_0_116555);
    
    \U_ELK12_CH/U_SLAVE_1ELK/Q[13]\ : DFN1C0
      port map(D => \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[13]_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/Q[13]_net_1\);
    
    HIEFFPLA_INST_0_52854 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_19[0]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_20[0]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_1[0]\, Y => 
        HIEFFPLA_NET_0_117500);
    
    HIEFFPLA_INST_0_45453 : AO1
      port map(A => HIEFFPLA_NET_0_119244, B => 
        \U50_PATTERNS/ELINK_DOUTA_2[2]\, C => 
        HIEFFPLA_NET_0_118810, Y => HIEFFPLA_NET_0_118911);
    
    HIEFFPLA_INST_0_37471 : MX2
      port map(A => \U200A_TFC/LOC_STRT_ADDR[3]\, B => 
        \TFC_STRT_ADDR[3]\, S => \U200A_TFC/GP_PG_SM_0[10]_net_1\, 
        Y => HIEFFPLA_NET_0_120279);
    
    \U_ELK4_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118067, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_1, Q => 
        \U_ELK4_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]_net_1\);
    
    \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[2]\ : DFN1C0
      port map(D => 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[2]_net_1\);
    
    HIEFFPLA_INST_0_62547 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_7[4]\, 
        B => HIEFFPLA_NET_0_117100, S => HIEFFPLA_NET_0_117174, Y
         => HIEFFPLA_NET_0_115976);
    
    HIEFFPLA_INST_0_56927 : NAND2B
      port map(A => HIEFFPLA_NET_0_116768, B => 
        HIEFFPLA_NET_0_117370, Y => HIEFFPLA_NET_0_116773);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_5[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116321, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_1, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_5[1]\);
    
    \U200A_TFC/ADDR_POINTER[6]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120356, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_30, Q => \TFC_ADDRB[6]\);
    
    HIEFFPLA_INST_0_61580 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_23[3]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_24[3]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[0]\, Y => 
        HIEFFPLA_NET_0_116106);
    
    HIEFFPLA_INST_0_58036 : NAND2A
      port map(A => HIEFFPLA_NET_0_116585, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_7[7]\, Y => 
        HIEFFPLA_NET_0_116573);
    
    \U_ELK4_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]\ : DFN1C0
      port map(D => \U_ELK4_CH/U_SLAVE_1ELK/Q[3]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]_net_1\);
    
    \U_ELK7_CH/ELK_IN_F\ : DFN1C0
      port map(D => \U_ELK7_CH/ELK_IN_DDR_F\, CLK => CCC_160M_ADJ, 
        CLR => DEV_RST_B_c, Q => \U_ELK7_CH/ELK_IN_F_net_1\);
    
    \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[14]\ : DFN1C0
      port map(D => 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[14]_net_1\);
    
    HIEFFPLA_INST_0_53094 : MX2
      port map(A => HIEFFPLA_NET_0_117554, B => 
        HIEFFPLA_NET_0_117550, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[2]\, Y => 
        HIEFFPLA_NET_0_117466);
    
    HIEFFPLA_INST_0_45043 : AO1A
      port map(A => \U50_PATTERNS/USB_TXE_B\, B => 
        HIEFFPLA_NET_0_119479, C => HIEFFPLA_NET_0_119375, Y => 
        HIEFFPLA_NET_0_118992);
    
    \U50_PATTERNS/U4D_REGCROSS/LOCAL_REG_VAL[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119084, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_3, Q => \ELKS_STOP_ADDR[7]\);
    
    HIEFFPLA_INST_0_56794 : XA1C
      port map(A => HIEFFPLA_NET_0_116805, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_0[5]\, C => 
        HIEFFPLA_NET_0_117179, Y => HIEFFPLA_NET_0_116795);
    
    HIEFFPLA_INST_0_53768 : AOI1D
      port map(A => HIEFFPLA_NET_0_117184, B => 
        HIEFFPLA_NET_0_117388, C => HIEFFPLA_NET_0_117336, Y => 
        HIEFFPLA_NET_0_117355);
    
    \U_ELK8_CH/U_SLAVE_1ELK/Q[4]\ : DFN1C0
      port map(D => \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/Q[4]_net_1\);
    
    HIEFFPLA_INST_0_48134 : MX2
      port map(A => \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[2]_net_1\, 
        B => \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\, S => 
        \BIT_OS_SEL_1[2]\, Y => HIEFFPLA_NET_0_118364);
    
    \U_ELK6_CH/U_ELK1_SERDAT_SOURCE/SERDAT[7]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117961, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_2, Q => 
        \U_ELK6_CH/ELK_TX_DAT[7]\);
    
    HIEFFPLA_INST_0_53795 : MX2
      port map(A => HIEFFPLA_NET_0_117290, B => 
        HIEFFPLA_NET_0_117408, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[2]_net_1\, Y
         => HIEFFPLA_NET_0_117351);
    
    \U200A_TFC/RX_SER_WORD_3DEL[7]\ : DFN1P0
      port map(D => \AFLSDF_INV_59\, CLK => CLK_40M_GL, PRE => 
        P_MASTER_POR_B_c_24, Q => 
        \U200A_TFC/RX_SER_WORD_3DEL_i_0[7]\);
    
    HIEFFPLA_INST_0_45695 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_19[3]\, C => 
        \U50_PATTERNS/SM_BANK_SEL[0]\, Y => HIEFFPLA_NET_0_118863);
    
    \U_ELK11_CH/U_ELK1_SERDAT_SOURCE/SERDAT[6]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118592, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_0, Q => 
        \U_ELK11_CH/ELK_TX_DAT[6]\);
    
    \U_ELK6_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117975, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_9, Q => 
        \U_ELK6_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]_net_1\);
    
    \U_ELK14_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL\ : DFN1C0
      port map(D => \U_ELK14_CH/ELK_IN_R_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL_net_1\);
    
    \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[6]\ : DFN1C0
      port map(D => 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\);
    
    HIEFFPLA_INST_0_56209 : NAND2A
      port map(A => HIEFFPLA_NET_0_116945, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/MAX_CNT[7]\, Y => 
        HIEFFPLA_NET_0_116929);
    
    \U_ELK3_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118107, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_12, Q => 
        \U_ELK3_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]_net_1\);
    
    \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[1]\ : DFN1C0
      port map(D => 
        \U_ELK1_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\);
    
    ELK0_SYNC_DET : DFN1C0
      port map(D => HIEFFPLA_NET_0_116926, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_25, Q => P_ELK0_SYNC_DET_c);
    
    \U_ELK0_CMD_TX/SER_OUT_FDEL\ : DFN1P0
      port map(D => \U_ELK0_CMD_TX/SER_OUT_FI_i\, CLK => 
        CCC_160M_FXD, PRE => MASTER_SALT_POR_B_i_0_i_10, Q => 
        ELK0_OUT_F_i_0);
    
    \U50_PATTERNS/REG_STATE[4]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119480, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_22_0, Q => 
        \U50_PATTERNS/REG_STATE[4]_net_1\);
    
    HIEFFPLA_INST_0_56073 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/MAX_CNT[1]\, 
        B => HIEFFPLA_NET_0_116938, S => HIEFFPLA_NET_0_117084, Y
         => HIEFFPLA_NET_0_116953);
    
    \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[9]\ : DFN1C0
      port map(D => 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\);
    
    \U50_PATTERNS/ELINK_ADDRA_0[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120091, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_18, Q => 
        \U50_PATTERNS/ELINK_ADDRA_0[4]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_30[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116355, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_18, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_30[1]\);
    
    \U_ELK16_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118377, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_10, Q => 
        \U_ELK16_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]_net_1\);
    
    HIEFFPLA_INST_0_53483 : MX2
      port map(A => HIEFFPLA_NET_0_117368, B => 
        HIEFFPLA_NET_0_117409, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[1]_net_1\, Y
         => HIEFFPLA_NET_0_117401);
    
    HIEFFPLA_INST_0_59525 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_28[3]\, B => 
        HIEFFPLA_NET_0_116815, S => HIEFFPLA_NET_0_117094, Y => 
        HIEFFPLA_NET_0_116383);
    
    HIEFFPLA_INST_0_51930 : AND3A
      port map(A => \U_MASTER_DES/U13A_ADJ_160M/BITCNT[5]\, B => 
        HIEFFPLA_NET_0_117684, C => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[31]_net_1\, Y => 
        HIEFFPLA_NET_0_117664);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_11[4]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116261, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_20, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_11[4]\);
    
    \U_ELK3_CH/U_SLAVE_1ELK/RECD_SER_WORD[2]\ : DFN1C0
      port map(D => \U_ELK3_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[2]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_3[2]\);
    
    \U_ELK15_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]\ : DFN1C0
      port map(D => \U_ELK15_CH/U_SLAVE_1ELK/Q[4]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]_net_1\);
    
    \U50_PATTERNS/ELINK_ADDRA_3[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119988, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_1, Q => 
        \U50_PATTERNS/ELINK_ADDRA_3[3]\);
    
    HIEFFPLA_INST_0_39920 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_9[6]\, B => 
        HIEFFPLA_NET_0_119517, S => HIEFFPLA_NET_0_119292, Y => 
        HIEFFPLA_NET_0_119937);
    
    \U_EXEC_MASTER/MPOR_B_4\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117787, CLK => CLK_40M_GL, CLR
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_1\, Q => 
        P_MASTER_POR_B_c_4);
    
    HIEFFPLA_INST_0_46877 : AND2A
      port map(A => \OP_MODE_c[1]\, B => \PATT_ELK_DAT_11[5]\, Y
         => HIEFFPLA_NET_0_118593);
    
    HIEFFPLA_INST_0_55066 : AND2A
      port map(A => HIEFFPLA_NET_0_117395, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[6]_net_1\, Y => 
        HIEFFPLA_NET_0_117129);
    
    \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[6]\ : DFN1C0
      port map(D => 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\);
    
    \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[9]\ : DFN1C0
      port map(D => \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\);
    
    \U50_PATTERNS/U4B_REGCROSS/DELCNT[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119134, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_30, Q => 
        \U50_PATTERNS/U4B_REGCROSS/DELCNT[0]_net_1\);
    
    HIEFFPLA_INST_0_57851 : XA1C
      port map(A => HIEFFPLA_NET_0_116604, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_6[8]\, C => 
        HIEFFPLA_NET_0_117179, Y => HIEFFPLA_NET_0_116607);
    
    \U50_PATTERNS/ELINK_DINA_5[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119745, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_14, Q => 
        \U50_PATTERNS/ELINK_DINA_5[6]\);
    
    HIEFFPLA_INST_0_44529 : XO1
      port map(A => \U50_PATTERNS/U4C_REGCROSS/SAMP_TWO[0]_net_1\, 
        B => \ELKS_STRT_ADDR[0]\, C => HIEFFPLA_NET_0_119097, Y
         => HIEFFPLA_NET_0_119101);
    
    HIEFFPLA_INST_0_41894 : AND2
      port map(A => HIEFFPLA_NET_0_119389, B => 
        \U50_PATTERNS/SM_BANK_SEL[13]\, Y => 
        HIEFFPLA_NET_0_119671);
    
    AFLSDF_INV_3 : INV
      port map(A => EXT_INT_REF_SEL_c, Y => \AFLSDF_INV_3\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_17[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116203, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_7, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_17[2]\);
    
    \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[0]\ : DFN1C0
      port map(D => 
        \U_ELK5_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\);
    
    HIEFFPLA_INST_0_49515 : MX2
      port map(A => HIEFFPLA_NET_0_118130, B => 
        HIEFFPLA_NET_0_118127, S => \BIT_OS_SEL_1[0]\, Y => 
        \U_ELK2_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[4]\);
    
    HIEFFPLA_INST_0_48905 : MX2
      port map(A => \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\, 
        B => \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\, S => 
        \BIT_OS_SEL[2]\, Y => HIEFFPLA_NET_0_118226);
    
    HIEFFPLA_INST_0_48768 : MX2
      port map(A => HIEFFPLA_NET_0_118269, B => 
        HIEFFPLA_NET_0_118267, S => \BIT_OS_SEL_2[0]\, Y => 
        \U_ELK18_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[4]\);
    
    \U50_PATTERNS/ELINK_DINA_14[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119829, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_16, Q => 
        \U50_PATTERNS/ELINK_DINA_14[2]\);
    
    HIEFFPLA_INST_0_45164 : NAND3C
      port map(A => HIEFFPLA_NET_0_118801, B => 
        HIEFFPLA_NET_0_118879, C => HIEFFPLA_NET_0_118964, Y => 
        HIEFFPLA_NET_0_118974);
    
    HIEFFPLA_INST_0_43479 : MX2
      port map(A => \U50_PATTERNS/SM_BANK_SEL[4]\, B => 
        HIEFFPLA_NET_0_119214, S => HIEFFPLA_NET_0_118691, Y => 
        HIEFFPLA_NET_0_119306);
    
    HIEFFPLA_INST_0_56109 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/MAX_CNT[5]\, 
        B => HIEFFPLA_NET_0_116934, S => HIEFFPLA_NET_0_117084, Y
         => HIEFFPLA_NET_0_116949);
    
    HIEFFPLA_INST_0_51192 : MX2
      port map(A => HIEFFPLA_NET_0_117816, B => 
        HIEFFPLA_NET_0_117812, S => \BIT_OS_SEL_3[1]\, Y => 
        HIEFFPLA_NET_0_117814);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_29[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116378, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_4, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_29[0]\);
    
    \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[14]\ : DFN1C0
      port map(D => \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[14]_net_1\);
    
    HIEFFPLA_INST_0_42197 : MX2
      port map(A => \U50_PATTERNS/OP_MODE_T[5]\, B => 
        \U50_PATTERNS/RD_USB_ADBUS[5]\, S => 
        HIEFFPLA_NET_0_119440, Y => HIEFFPLA_NET_0_119604);
    
    HIEFFPLA_INST_0_43946 : MX2
      port map(A => HIEFFPLA_NET_0_119567, B => 
        \U50_PATTERNS/TFC_DINA[5]\, S => HIEFFPLA_NET_0_119294, Y
         => HIEFFPLA_NET_0_119192);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_31[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116020, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_9, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_31[0]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_28[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116384, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_2, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_28[2]\);
    
    HIEFFPLA_INST_0_48465 : MX2
      port map(A => \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\, 
        B => \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[13]_net_1\, S => 
        \BIT_OS_SEL_0[2]\, Y => HIEFFPLA_NET_0_118307);
    
    \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[2]\ : DFN1C0
      port map(D => \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\);
    
    HIEFFPLA_INST_0_39398 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_2[4]\, B => 
        HIEFFPLA_NET_0_119519, S => HIEFFPLA_NET_0_119278, Y => 
        HIEFFPLA_NET_0_119995);
    
    HIEFFPLA_INST_0_56492 : AO1
      port map(A => HIEFFPLA_NET_0_117428, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[8]_net_1\, C => 
        HIEFFPLA_NET_0_116836, Y => HIEFFPLA_NET_0_116852);
    
    \U_ELK19_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL\ : DFN1C0
      port map(D => \U_ELK19_CH/ELK_IN_R_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL_net_1\);
    
    \U50_PATTERNS/ELINK_ADDRA_16[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120037, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_8, Q => 
        \U50_PATTERNS/ELINK_ADDRA_16[2]\);
    
    HIEFFPLA_INST_0_61481 : MX2
      port map(A => HIEFFPLA_NET_0_117190, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_23[0]\, S => 
        HIEFFPLA_NET_0_117151, Y => HIEFFPLA_NET_0_116120);
    
    HIEFFPLA_INST_0_42898 : AND2A
      port map(A => \U50_PATTERNS/REG_STATE[5]_net_1\, B => 
        \U50_PATTERNS/REG_STATE[2]_net_1\, Y => 
        HIEFFPLA_NET_0_119430);
    
    HIEFFPLA_INST_0_49427 : MX2
      port map(A => HIEFFPLA_NET_0_118129, B => 
        HIEFFPLA_NET_0_118139, S => \BIT_OS_SEL[1]\, Y => 
        HIEFFPLA_NET_0_118132);
    
    HIEFFPLA_INST_0_50776 : MX2
      port map(A => HIEFFPLA_NET_0_117915, B => 
        HIEFFPLA_NET_0_117913, S => \BIT_OS_SEL[0]\, Y => 
        \U_ELK7_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[6]\);
    
    HIEFFPLA_INST_0_37465 : MX2
      port map(A => \U200A_TFC/LOC_STRT_ADDR[2]\, B => 
        \TFC_STRT_ADDR[2]\, S => \U200A_TFC/GP_PG_SM_0[10]_net_1\, 
        Y => HIEFFPLA_NET_0_120280);
    
    HIEFFPLA_INST_0_44600 : MX2
      port map(A => \ELKS_STOP_ADDR[6]\, B => 
        \U50_PATTERNS/U4D_REGCROSS/SAMP_TWO[6]_net_1\, S => 
        HIEFFPLA_NET_0_119093, Y => HIEFFPLA_NET_0_119085);
    
    HIEFFPLA_INST_0_41961 : AND3C
      port map(A => HIEFFPLA_NET_0_119255, B => 
        HIEFFPLA_NET_0_119262, C => 
        \U50_PATTERNS/SM_BANK_SEL[15]\, Y => 
        HIEFFPLA_NET_0_119645);
    
    HIEFFPLA_INST_0_51312 : MX2
      port map(A => \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\, 
        B => \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[14]_net_1\, S => 
        \BIT_OS_SEL_5[2]\, Y => HIEFFPLA_NET_0_117798);
    
    HIEFFPLA_INST_0_54719 : NAND3B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[1]_net_1\, B => 
        HIEFFPLA_NET_0_117246, C => HIEFFPLA_NET_0_117251, Y => 
        HIEFFPLA_NET_0_117218);
    
    HIEFFPLA_INST_0_51017 : MX2
      port map(A => HIEFFPLA_NET_0_117859, B => 
        HIEFFPLA_NET_0_117869, S => \BIT_OS_SEL_5[0]\, Y => 
        \U_ELK8_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[5]\);
    
    \U_EXEC_MASTER/MPOR_SALT_B_6\ : DFI1P0
      port map(D => HIEFFPLA_NET_0_117781, CLK => CLK_40M_GL, PRE
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_2\, QN => 
        MASTER_SALT_POR_B_i_0_i_6);
    
    HIEFFPLA_INST_0_46248 : AO1
      port map(A => HIEFFPLA_NET_0_119476, B => 
        \U50_PATTERNS/CHKSUM[1]\, C => HIEFFPLA_NET_0_118904, Y
         => HIEFFPLA_NET_0_118732);
    
    HIEFFPLA_INST_0_45760 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_9[3]\, C => 
        \U50_PATTERNS/SM_BANK_SEL[10]\, Y => 
        HIEFFPLA_NET_0_118850);
    
    HIEFFPLA_INST_0_39749 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_7[3]\, B => 
        HIEFFPLA_NET_0_119520, S => HIEFFPLA_NET_0_119289, Y => 
        HIEFFPLA_NET_0_119956);
    
    HIEFFPLA_INST_0_57519 : XA1B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_4[7]\, B => 
        HIEFFPLA_NET_0_116682, C => HIEFFPLA_NET_0_117179, Y => 
        HIEFFPLA_NET_0_116664);
    
    \U_ELK6_CH/U_ELK1_CMD_TX/SER_OUT_RDEL\ : DFN1C0
      port map(D => \U_ELK6_CH/U_ELK1_CMD_TX/SER_OUT_RI_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_16, Q
         => \U_ELK6_CH/ELK_OUT_R\);
    
    \U200B_ELINKS/RX_SER_WORD_2DEL[6]\ : DFN1C0
      port map(D => \U200B_ELINKS/RX_SER_WORD_1DEL[6]_net_1\, CLK
         => CLK_40M_GL, CLR => P_MASTER_POR_B_c_26, Q => 
        \U200B_ELINKS/RX_SER_WORD_2DEL[6]_net_1\);
    
    HIEFFPLA_INST_0_55715 : MX2
      port map(A => HIEFFPLA_NET_0_115971, B => 
        HIEFFPLA_NET_0_116224, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_2[3]\, Y => 
        HIEFFPLA_NET_0_117000);
    
    HIEFFPLA_INST_0_56448 : AND3
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[10]_net_1\, B
         => HIEFFPLA_NET_0_117427, C => HIEFFPLA_NET_0_117423, Y
         => HIEFFPLA_NET_0_116865);
    
    HIEFFPLA_INST_0_52558 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_1[0]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_2[0]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[0]\, Y => 
        HIEFFPLA_NET_0_117548);
    
    HIEFFPLA_INST_0_49306 : MX2
      port map(A => HIEFFPLA_NET_0_118173, B => 
        HIEFFPLA_NET_0_118158, S => \BIT_OS_SEL_1[1]\, Y => 
        HIEFFPLA_NET_0_118160);
    
    HIEFFPLA_INST_0_46160 : AO1
      port map(A => HIEFFPLA_NET_0_119241, B => 
        \U50_PATTERNS/ELINK_DOUTA_1[1]\, C => 
        HIEFFPLA_NET_0_118928, Y => HIEFFPLA_NET_0_118753);
    
    \U_ELK8_CH/U_SLAVE_1ELK/Q[10]\ : DFN1C0
      port map(D => \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/Q[10]_net_1\);
    
    \U_ELK6_CH/U_SLAVE_1ELK/RECD_SER_WORD[7]\ : DFN1C0
      port map(D => \U_ELK6_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[7]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_6[7]\);
    
    HIEFFPLA_INST_0_54520 : MX2
      port map(A => HIEFFPLA_NET_0_117317, B => 
        HIEFFPLA_NET_0_117299, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[2]_net_1\, Y => 
        HIEFFPLA_NET_0_117255);
    
    HIEFFPLA_INST_0_40190 : AOI1D
      port map(A => HIEFFPLA_NET_0_119389, B => 
        HIEFFPLA_NET_0_119464, C => \U50_PATTERNS/SM_BANK_SEL[5]\, 
        Y => HIEFFPLA_NET_0_119877);
    
    HIEFFPLA_INST_0_51444 : AND2A
      port map(A => HIEFFPLA_NET_0_117771, B => 
        \U_EXEC_MASTER/CCC_1_LOCK_STAT_1D_net_1\, Y => 
        HIEFFPLA_NET_0_117772);
    
    \U_ELK12_CH/U_SLAVE_1ELK/Q[9]\ : DFN1C0
      port map(D => \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/Q[9]_net_1\);
    
    HIEFFPLA_INST_0_37400 : AO1C
      port map(A => \U200A_TFC/N_232_li\, B => ALIGN_ACTIVE, C
         => P_USB_MASTER_EN_c_22_0, Y => HIEFFPLA_NET_0_120291);
    
    \U50_PATTERNS/ELINK_BLKA[17]/U1\ : DFN1P0
      port map(D => HIEFFPLA_NET_0_119927, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_20, Q => 
        \U50_PATTERNS/ELINK_BLKA[17]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_13[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116249, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_1, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_13[1]\);
    
    \U_ELK6_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117977, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_9, Q => 
        \U_ELK6_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]_net_1\);
    
    HIEFFPLA_INST_0_38633 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_10[7]\, B => 
        HIEFFPLA_NET_0_119516, S => HIEFFPLA_NET_0_119239, Y => 
        HIEFFPLA_NET_0_120080);
    
    HIEFFPLA_INST_0_58002 : AND3B
      port map(A => HIEFFPLA_NET_0_117179, B => 
        HIEFFPLA_NET_0_116575, C => HIEFFPLA_NET_0_116590, Y => 
        HIEFFPLA_NET_0_116580);
    
    HIEFFPLA_INST_0_56653 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_0[2]\, B => 
        HIEFFPLA_NET_0_116798, S => HIEFFPLA_NET_0_117602, Y => 
        HIEFFPLA_NET_0_116822);
    
    HIEFFPLA_INST_0_55173 : AND3B
      port map(A => HIEFFPLA_NET_0_117071, B => 
        HIEFFPLA_NET_0_117105, C => HIEFFPLA_NET_0_117086, Y => 
        HIEFFPLA_NET_0_117106);
    
    \U_ELK19_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]\ : DFN1C0
      port map(D => \U_ELK19_CH/U_SLAVE_1ELK/Q[9]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]_net_1\);
    
    \U_ELK8_CH/U_SLAVE_1ELK/Q[1]\ : DFN1C0
      port map(D => \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/Q[1]_net_1\);
    
    \U_ELK12_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118556, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_12, Q => 
        \U_ELK12_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]_net_1\);
    
    HIEFFPLA_INST_0_56960 : AOI1A
      port map(A => HIEFFPLA_NET_0_116779, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_1[0]\, C => 
        HIEFFPLA_NET_0_116764, Y => HIEFFPLA_NET_0_116765);
    
    \U50_PATTERNS/ELINK_DINA_15[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119820, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_16, Q => 
        \U50_PATTERNS/ELINK_DINA_15[3]\);
    
    HIEFFPLA_INST_0_42961 : AND3C
      port map(A => \U50_PATTERNS/REG_STATE[5]_net_1\, B => 
        \U50_PATTERNS/WR_XFER_TYPE[1]_net_1\, C => 
        HIEFFPLA_NET_0_118692, Y => HIEFFPLA_NET_0_119415);
    
    \U50_PATTERNS/USB_OE_BI/U1\ : DFN1P0
      port map(D => HIEFFPLA_NET_0_119045, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_19, Q => USB_OE_BI);
    
    HIEFFPLA_INST_0_45630 : NAND3C
      port map(A => HIEFFPLA_NET_0_118710, B => 
        HIEFFPLA_NET_0_118720, C => HIEFFPLA_NET_0_118729, Y => 
        HIEFFPLA_NET_0_118877);
    
    HIEFFPLA_INST_0_42735 : AND3C
      port map(A => HIEFFPLA_NET_0_119379, B => 
        \U50_PATTERNS/REG_STATE_0[4]_net_1\, C => 
        HIEFFPLA_NET_0_119442, Y => HIEFFPLA_NET_0_119472);
    
    HIEFFPLA_INST_0_61991 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_12[0]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_28[0]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_3[4]_net_1\, Y
         => HIEFFPLA_NET_0_116050);
    
    HIEFFPLA_INST_0_54738 : NAND3B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[3]_net_1\, B => 
        HIEFFPLA_NET_0_117238, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[0]_net_1\, Y => 
        HIEFFPLA_NET_0_117212);
    
    HIEFFPLA_INST_0_62373 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_4[3]\, 
        B => HIEFFPLA_NET_0_117075, S => HIEFFPLA_NET_0_117148, Y
         => HIEFFPLA_NET_0_115997);
    
    HIEFFPLA_INST_0_57431 : AO1A
      port map(A => HIEFFPLA_NET_0_116681, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_4[3]\, C => 
        HIEFFPLA_NET_0_116685, Y => HIEFFPLA_NET_0_116686);
    
    HIEFFPLA_INST_0_52227 : AND3
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[7]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[2]_net_1\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[7]_net_1\, Y => 
        HIEFFPLA_NET_0_117606);
    
    HIEFFPLA_INST_0_46816 : MX2
      port map(A => HIEFFPLA_NET_0_118626, B => 
        HIEFFPLA_NET_0_118608, S => \BIT_OS_SEL[1]\, Y => 
        HIEFFPLA_NET_0_118610);
    
    HIEFFPLA_INST_0_55691 : MX2
      port map(A => HIEFFPLA_NET_0_115974, B => 
        HIEFFPLA_NET_0_116217, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_2[3]\, Y => 
        HIEFFPLA_NET_0_117003);
    
    HIEFFPLA_INST_0_50116 : NAND2B
      port map(A => \OP_MODE_c_5[1]\, B => \PATT_ELK_DAT_5[7]\, Y
         => HIEFFPLA_NET_0_118006);
    
    \U_ELK16_CH/U_SLAVE_1ELK/Q[7]\ : DFN1C0
      port map(D => \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/Q[7]_net_1\);
    
    \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_2S_1\ : DFN1C0
      port map(D => 
        \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_1S_net_1\, CLK
         => CLK60MHZ, CLR => P_MASTER_POR_B_c_0_0, Q => 
        P_USB_MASTER_EN_c_1);
    
    HIEFFPLA_INST_0_47885 : MX2
      port map(A => \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[2]_net_1\, 
        B => \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\, S => 
        \BIT_OS_SEL_1[2]\, Y => HIEFFPLA_NET_0_118409);
    
    HIEFFPLA_INST_0_46376 : AO1
      port map(A => HIEFFPLA_NET_0_119241, B => 
        \U50_PATTERNS/ELINK_DOUTA_1[0]\, C => 
        HIEFFPLA_NET_0_118845, Y => HIEFFPLA_NET_0_118703);
    
    HIEFFPLA_INST_0_60324 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_9[0]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_25[0]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[4]_net_1\, Y
         => HIEFFPLA_NET_0_116281);
    
    \U_ELK4_CH/U_SLAVE_1ELK/RECD_SER_WORD[2]\ : DFN1C0
      port map(D => \U_ELK4_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[2]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_4[2]\);
    
    HIEFFPLA_INST_0_44971 : AO1A
      port map(A => HIEFFPLA_NET_0_118991, B => 
        HIEFFPLA_NET_0_119632, C => HIEFFPLA_NET_0_119298, Y => 
        HIEFFPLA_NET_0_119009);
    
    \U_ELK19_CH/U_SLAVE_1ELK/Q[7]\ : DFN1C0
      port map(D => \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/Q[7]_net_1\);
    
    \U_ELK13_CH/U_SLAVE_1ELK/RECD_SER_WORD[2]\ : DFN1C0
      port map(D => \U_ELK13_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[2]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_13[2]\);
    
    HIEFFPLA_INST_0_43560 : AND2B
      port map(A => \U50_PATTERNS/SM_BANK_SEL[20]\, B => 
        \U50_PATTERNS/SM_BANK_SEL_0[21]\, Y => 
        HIEFFPLA_NET_0_119294);
    
    HIEFFPLA_INST_0_61091 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_3[1]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_19[1]\, S
         => \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_1[4]_net_1\, 
        Y => HIEFFPLA_NET_0_116175);
    
    HIEFFPLA_INST_0_62996 : NAND3A
      port map(A => HIEFFPLA_NET_0_115905, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[4]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[3]\, Y => 
        HIEFFPLA_NET_0_115920);
    
    \U50_PATTERNS/ELINK_ADDRA_13[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120056, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_3, Q => 
        \U50_PATTERNS/ELINK_ADDRA_13[7]\);
    
    \U_ELK5_CH/U_SLAVE_1ELK/RECD_SER_WORD[4]\ : DFN1C0
      port map(D => \U_ELK5_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[4]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_5[4]\);
    
    HIEFFPLA_INST_0_43533 : MX2
      port map(A => \U50_PATTERNS/SM_BANK_SEL_0[20]\, B => 
        HIEFFPLA_NET_0_119467, S => HIEFFPLA_NET_0_118691, Y => 
        HIEFFPLA_NET_0_119300);
    
    HIEFFPLA_INST_0_46581 : AND2A
      port map(A => \OP_MODE_c_4[1]\, B => \PATT_ELK_DAT_0[5]\, Y
         => HIEFFPLA_NET_0_118655);
    
    HIEFFPLA_INST_0_45977 : NAND3C
      port map(A => HIEFFPLA_NET_0_118942, B => 
        HIEFFPLA_NET_0_118953, C => HIEFFPLA_NET_0_118698, Y => 
        HIEFFPLA_NET_0_118798);
    
    \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[1]\ : DFN1C0
      port map(D => 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[1]_net_1\);
    
    HIEFFPLA_INST_0_61649 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_8[3]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_24[3]\, S
         => \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_4[4]_net_1\, 
        Y => HIEFFPLA_NET_0_116097);
    
    HIEFFPLA_INST_0_59474 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_11[0]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_27[0]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_5[4]_net_1\, Y
         => HIEFFPLA_NET_0_116390);
    
    \U_TFC_CMD_TX/SER_CMD_WORD_F[0]\ : DFN1C0
      port map(D => \U_TFC_CMD_TX/N_SER_CMD_WORD_F[0]\, CLK => 
        CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_TFC_CMD_TX/SER_CMD_WORD_F[0]_net_1\);
    
    HIEFFPLA_INST_0_54747 : AND3A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[1]_net_1\, B => 
        HIEFFPLA_NET_0_117251, C => HIEFFPLA_NET_0_117244, Y => 
        HIEFFPLA_NET_0_117209);
    
    HIEFFPLA_INST_0_161261 : DFN1C0
      port map(D => \TFC_IN_F\, CLK => CCC_160M_ADJ, CLR => 
        P_MASTER_POR_B_c_31_0, Q => HIEFFPLA_NET_0_161294);
    
    HIEFFPLA_INST_0_50833 : MX2
      port map(A => 
        \U_ELK8_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]_net_1\, B => 
        \U_ELK8_CH/ELK_TX_DAT[6]\, S => 
        \U_ELK8_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_117884);
    
    HIEFFPLA_INST_0_48527 : MX2
      port map(A => HIEFFPLA_NET_0_118313, B => 
        HIEFFPLA_NET_0_118308, S => \BIT_OS_SEL_3[0]\, Y => 
        \U_ELK17_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[5]\);
    
    HIEFFPLA_INST_0_59014 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_22[3]\, B => 
        HIEFFPLA_NET_0_116815, S => HIEFFPLA_NET_0_117095, Y => 
        HIEFFPLA_NET_0_116447);
    
    HIEFFPLA_INST_0_55826 : MX2
      port map(A => HIEFFPLA_NET_0_117018, B => 
        HIEFFPLA_NET_0_117006, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[2]\, Y => 
        HIEFFPLA_NET_0_116985);
    
    HIEFFPLA_INST_0_58412 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_14[3]\, B => 
        HIEFFPLA_NET_0_116521, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_1[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116525);
    
    HIEFFPLA_INST_0_47376 : AND2A
      port map(A => \OP_MODE_c[1]\, B => \PATT_ELK_DAT_13[6]\, Y
         => HIEFFPLA_NET_0_118502);
    
    \U_ELK1_CH/U_SLAVE_1ELK/Q[3]\ : DFN1C0
      port map(D => \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/Q[3]_net_1\);
    
    \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[5]\ : DFN1C0
      port map(D => 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\);
    
    HIEFFPLA_INST_0_43747 : AND3A
      port map(A => \U50_PATTERNS/RD_USB_ADBUS[3]\, B => 
        HIEFFPLA_NET_0_119592, C => 
        \U50_PATTERNS/RD_USB_ADBUS[2]\, Y => 
        HIEFFPLA_NET_0_119224);
    
    HIEFFPLA_INST_0_43635 : AND2B
      port map(A => \U50_PATTERNS/SM_BANK_SEL[21]\, B => 
        \U50_PATTERNS/SM_BANK_SEL[2]\, Y => HIEFFPLA_NET_0_119260);
    
    HIEFFPLA_INST_0_62400 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_5[1]\, 
        B => HIEFFPLA_NET_0_117114, S => HIEFFPLA_NET_0_117172, Y
         => HIEFFPLA_NET_0_115994);
    
    HIEFFPLA_INST_0_48294 : MX2
      port map(A => HIEFFPLA_NET_0_118351, B => 
        HIEFFPLA_NET_0_118340, S => \BIT_OS_SEL_3[0]\, Y => 
        \U_ELK16_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[7]\);
    
    \U50_PATTERNS/U4E_REGCROSS/SAMP_TWO[4]\ : DFN1C0
      port map(D => \U50_PATTERNS/U4E_REGCROSS/SAMP_ONE[4]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_23, Q => 
        \U50_PATTERNS/U4E_REGCROSS/SAMP_TWO[4]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_26[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116079, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_12, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_26[1]\);
    
    \U_ELK19_CH/U_SLAVE_1ELK/RECD_SER_WORD[1]\ : DFN1C0
      port map(D => \U_ELK19_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[1]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_19[1]\);
    
    HIEFFPLA_INST_0_61022 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_2[2]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_18[2]\, S
         => \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_4[4]_net_1\, 
        Y => HIEFFPLA_NET_0_116184);
    
    \U50_PATTERNS/TFC_STRT_ADDR_T[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119162, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_4, Q => 
        \U50_PATTERNS/TFC_STRT_ADDR_T[2]\);
    
    HIEFFPLA_INST_0_50278 : MX2
      port map(A => HIEFFPLA_NET_0_117990, B => 
        HIEFFPLA_NET_0_118004, S => \BIT_OS_SEL_0[0]\, Y => 
        \U_ELK5_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[6]\);
    
    \U_ELK17_CH/U_SLAVE_1ELK/Q[14]\ : DFN1C0
      port map(D => \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[14]_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/Q[14]_net_1\);
    
    HIEFFPLA_INST_0_56226 : AND3C
      port map(A => \ELK_RX_SER_WORD_0[5]\, B => 
        \ELK_RX_SER_WORD_0[4]\, C => HIEFFPLA_NET_0_116925, Y => 
        HIEFFPLA_NET_0_116926);
    
    \U_ELK2_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118150, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_8, Q => 
        \U_ELK2_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]_net_1\);
    
    \U50_PATTERNS/ELINKS_STOP_ADDR_T[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120116, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_7, Q => 
        \U50_PATTERNS/ELINKS_STOP_ADDR_T[3]\);
    
    \P_OP_MODE1_SPE_pad/U0/U0\ : IOPAD_TRI_U
      port map(D => \P_OP_MODE1_SPE_pad/U0/NET1\, E => 
        \P_OP_MODE1_SPE_pad/U0/NET2\, PAD => P_OP_MODE1_SPE);
    
    HIEFFPLA_INST_0_40050 : MX2
      port map(A => HIEFFPLA_NET_0_119886, B => 
        \U50_PATTERNS/ELINK_BLKA[6]\, S => 
        \U50_PATTERNS/SM_BANK_SEL[20]\, Y => 
        HIEFFPLA_NET_0_119919);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_15[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116227, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_4, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_15[3]\);
    
    HIEFFPLA_INST_0_62502 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_6[4]\, 
        B => HIEFFPLA_NET_0_117100, S => HIEFFPLA_NET_0_117132, Y
         => HIEFFPLA_NET_0_115981);
    
    HIEFFPLA_INST_0_43567 : AND2A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/SM_BANK_SEL[3]\, Y => HIEFFPLA_NET_0_119288);
    
    \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[1]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_SER_IN_F_1DEL_net_1\, 
        CLK => CCC_160M_ADJ, CLR => P_MASTER_POR_B_c_34_0, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[1]_net_1\);
    
    \U_ELK13_CH/U_SLAVE_1ELK/Q[9]\ : DFN1C0
      port map(D => \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/Q[9]_net_1\);
    
    HIEFFPLA_INST_0_52594 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_9[2]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_10[2]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[0]\, Y => 
        HIEFFPLA_NET_0_117542);
    
    HIEFFPLA_INST_0_38242 : MX2
      port map(A => \U50_PATTERNS/ELINKS_STOP_ADDR[0]\, B => 
        \U50_PATTERNS/ELINKS_STOP_ADDR_T[0]\, S => 
        HIEFFPLA_NET_0_119472, Y => HIEFFPLA_NET_0_120127);
    
    \U_ELK14_CH/U_ELK1_SERDAT_SOURCE/SERDAT[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118463, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_6, Q => 
        \U_ELK14_CH/ELK_TX_DAT[0]\);
    
    \U50_PATTERNS/U106_PATT_ELINK_BLK/DPRT_512X9_SRAM_R0C0\ : 
        RAM4K9
      generic map(MEMORYFILE => "DPRT_512X9_SRAM_R0C0.mem")

      port map(ADDRA11 => AFLSDF_GND, ADDRA10 => AFLSDF_GND, 
        ADDRA9 => AFLSDF_GND, ADDRA8 => \GND\, ADDRA7 => 
        \U50_PATTERNS/ELINK_ADDRA_6[7]\, ADDRA6 => 
        \U50_PATTERNS/ELINK_ADDRA_6[6]\, ADDRA5 => 
        \U50_PATTERNS/ELINK_ADDRA_6[5]\, ADDRA4 => 
        \U50_PATTERNS/ELINK_ADDRA_6[4]\, ADDRA3 => 
        \U50_PATTERNS/ELINK_ADDRA_6[3]\, ADDRA2 => 
        \U50_PATTERNS/ELINK_ADDRA_6[2]\, ADDRA1 => 
        \U50_PATTERNS/ELINK_ADDRA_6[1]\, ADDRA0 => 
        \U50_PATTERNS/ELINK_ADDRA_6[0]\, ADDRB11 => AFLSDF_GND, 
        ADDRB10 => AFLSDF_GND, ADDRB9 => AFLSDF_GND, ADDRB8 => 
        \GND\, ADDRB7 => \ELKS_ADDRB[7]\, ADDRB6 => 
        \ELKS_ADDRB_0[6]\, ADDRB5 => \ELKS_ADDRB[5]\, ADDRB4 => 
        \ELKS_ADDRB_0[4]\, ADDRB3 => \ELKS_ADDRB[3]\, ADDRB2 => 
        \ELKS_ADDRB_0[2]\, ADDRB1 => \ELKS_ADDRB[1]\, ADDRB0 => 
        \ELKS_ADDRB[0]\, DINA8 => \GND\, DINA7 => 
        \U50_PATTERNS/ELINK_DINA_6[7]\, DINA6 => 
        \U50_PATTERNS/ELINK_DINA_6[6]\, DINA5 => 
        \U50_PATTERNS/ELINK_DINA_6[5]\, DINA4 => 
        \U50_PATTERNS/ELINK_DINA_6[4]\, DINA3 => 
        \U50_PATTERNS/ELINK_DINA_6[3]\, DINA2 => 
        \U50_PATTERNS/ELINK_DINA_6[2]\, DINA1 => 
        \U50_PATTERNS/ELINK_DINA_6[1]\, DINA0 => 
        \U50_PATTERNS/ELINK_DINA_6[0]\, DINB8 => \GND\, DINB7 => 
        \ELK_RX_SER_WORD_6[7]\, DINB6 => \ELK_RX_SER_WORD_6[6]\, 
        DINB5 => \ELK_RX_SER_WORD_6[5]\, DINB4 => 
        \ELK_RX_SER_WORD_6[4]\, DINB3 => \ELK_RX_SER_WORD_6[3]\, 
        DINB2 => \ELK_RX_SER_WORD_6[2]\, DINB1 => 
        \ELK_RX_SER_WORD_6[1]\, DINB0 => \ELK_RX_SER_WORD_6[0]\, 
        WIDTHA0 => \VCC\, WIDTHA1 => \VCC\, WIDTHB0 => \VCC\, 
        WIDTHB1 => \VCC\, PIPEA => \VCC\, PIPEB => \VCC\, WMODEA
         => \GND\, WMODEB => \GND\, BLKA => 
        \U50_PATTERNS/ELINK_BLKA[6]\, BLKB => ELKS_RAM_BLKB_EN, 
        WENA => \U50_PATTERNS/ELINK_RWA[6]\, WENB => ELKS_RWB, 
        CLKA => CLK60MHZ, CLKB => CLK_40M_GL, RESET => 
        P_USB_MASTER_EN_c_0, DOUTA8 => OPEN, DOUTA7 => 
        \U50_PATTERNS/ELINK_DOUTA_6[7]\, DOUTA6 => 
        \U50_PATTERNS/ELINK_DOUTA_6[6]\, DOUTA5 => 
        \U50_PATTERNS/ELINK_DOUTA_6[5]\, DOUTA4 => 
        \U50_PATTERNS/ELINK_DOUTA_6[4]\, DOUTA3 => 
        \U50_PATTERNS/ELINK_DOUTA_6[3]\, DOUTA2 => 
        \U50_PATTERNS/ELINK_DOUTA_6[2]\, DOUTA1 => 
        \U50_PATTERNS/ELINK_DOUTA_6[1]\, DOUTA0 => 
        \U50_PATTERNS/ELINK_DOUTA_6[0]\, DOUTB8 => OPEN, DOUTB7
         => \PATT_ELK_DAT_6[7]\, DOUTB6 => \PATT_ELK_DAT_6[6]\, 
        DOUTB5 => \PATT_ELK_DAT_6[5]\, DOUTB4 => 
        \PATT_ELK_DAT_6[4]\, DOUTB3 => \PATT_ELK_DAT_6[3]\, 
        DOUTB2 => \PATT_ELK_DAT_6[2]\, DOUTB1 => 
        \PATT_ELK_DAT_6[1]\, DOUTB0 => \PATT_ELK_DAT_6[0]\);
    
    HIEFFPLA_INST_0_50857 : NAND2B
      port map(A => \OP_MODE_c_0[1]\, B => \PATT_ELK_DAT_8[1]\, Y
         => HIEFFPLA_NET_0_117877);
    
    HIEFFPLA_INST_0_47111 : MX2
      port map(A => 
        \U_ELK12_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]_net_1\, B => 
        \U_ELK12_CH/ELK_TX_DAT[5]\, S => 
        \U_ELK12_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118556);
    
    HIEFFPLA_INST_0_42240 : AND3C
      port map(A => \U50_PATTERNS/RD_USB_ADBUS[1]\, B => 
        \U50_PATTERNS/RD_USB_ADBUS[0]\, C => 
        HIEFFPLA_NET_0_119208, Y => HIEFFPLA_NET_0_119594);
    
    HIEFFPLA_INST_0_38615 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_10[5]\, B => 
        HIEFFPLA_NET_0_119518, S => HIEFFPLA_NET_0_119239, Y => 
        HIEFFPLA_NET_0_120082);
    
    HIEFFPLA_INST_0_54822 : MX2
      port map(A => HIEFFPLA_NET_0_116183, B => 
        HIEFFPLA_NET_0_116072, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[3]_net_1\, Y => 
        HIEFFPLA_NET_0_117195);
    
    HIEFFPLA_INST_0_54840 : NAND2B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[1]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[5]_net_1\, Y => 
        HIEFFPLA_NET_0_117192);
    
    HIEFFPLA_INST_0_43743 : AND3A
      port map(A => \U50_PATTERNS/RD_USB_ADBUS[3]\, B => 
        HIEFFPLA_NET_0_119591, C => 
        \U50_PATTERNS/RD_USB_ADBUS[2]\, Y => 
        HIEFFPLA_NET_0_119225);
    
    HIEFFPLA_INST_0_40999 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_19[5]\, B => 
        HIEFFPLA_NET_0_119567, S => HIEFFPLA_NET_0_119293, Y => 
        HIEFFPLA_NET_0_119786);
    
    \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[4]\ : DFN1C0
      port map(D => \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\);
    
    HIEFFPLA_INST_0_44664 : MX2
      port map(A => \OP_MODE_c[1]\, B => 
        \U50_PATTERNS/U4E_REGCROSS/SAMP_TWO[1]_net_1\, S => 
        HIEFFPLA_NET_0_119072, Y => HIEFFPLA_NET_0_119069);
    
    HIEFFPLA_INST_0_45747 : AO1
      port map(A => HIEFFPLA_NET_0_119254, B => 
        \U50_PATTERNS/ELINK_DOUTA_6[0]\, C => 
        HIEFFPLA_NET_0_118769, Y => HIEFFPLA_NET_0_118853);
    
    \U_ELK14_CH/ELK_IN_R\ : DFN1C0
      port map(D => \U_ELK14_CH/ELK_IN_DDR_R\, CLK => 
        CCC_160M_ADJ, CLR => DEV_RST_B_c, Q => 
        \U_ELK14_CH/ELK_IN_R_net_1\);
    
    \U50_PATTERNS/TFC_STOP_ADDR[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119185, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_8, Q => 
        \U50_PATTERNS/TFC_STOP_ADDR[3]\);
    
    HIEFFPLA_INST_0_53927 : MX2
      port map(A => HIEFFPLA_NET_0_117309, B => 
        HIEFFPLA_NET_0_117302, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[2]_net_1\, Y
         => HIEFFPLA_NET_0_117332);
    
    HIEFFPLA_INST_0_46088 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_7[0]\, C => 
        \U50_PATTERNS/SM_BANK_SEL[12]\, Y => 
        HIEFFPLA_NET_0_118769);
    
    \U50_PATTERNS/ELINK_ADDRA_12[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120068, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_2_0, Q => 
        \U50_PATTERNS/ELINK_ADDRA_12[3]\);
    
    HIEFFPLA_INST_0_42286 : AND2B
      port map(A => \U50_PATTERNS/RD_USB_ADBUS[0]\, B => 
        \U50_PATTERNS/RD_USB_ADBUS[7]\, Y => 
        HIEFFPLA_NET_0_119582);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_25[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116093, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_10, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_25[2]\);
    
    HIEFFPLA_INST_0_42559 : AND3B
      port map(A => \U50_PATTERNS/REG_ADDR[8]\, B => 
        HIEFFPLA_NET_0_119509, C => \U50_PATTERNS/REG_ADDR[7]\, Y
         => HIEFFPLA_NET_0_119511);
    
    \U_ELK4_CH/U_SLAVE_1ELK/Q[4]\ : DFN1C0
      port map(D => \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/Q[4]_net_1\);
    
    \U_ELK19_CH/U_ELK1_SERDAT_SOURCE/SERDAT[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118238, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_15, Q => 
        \U_ELK19_CH/ELK_TX_DAT[0]\);
    
    HIEFFPLA_INST_0_48069 : MX2
      port map(A => \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[0]_net_1\, 
        B => \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\, S => 
        \BIT_OS_SEL_1[2]\, Y => HIEFFPLA_NET_0_118384);
    
    HIEFFPLA_INST_0_42805 : AND3C
      port map(A => HIEFFPLA_NET_0_119573, B => 
        \U50_PATTERNS/REG_STATE_0[4]_net_1\, C => 
        HIEFFPLA_NET_0_119412, Y => HIEFFPLA_NET_0_119459);
    
    \U_EXEC_MASTER/MPOR_SALT_B_8\ : DFI1P0
      port map(D => HIEFFPLA_NET_0_117781, CLK => CLK_40M_GL, PRE
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_2\, QN => 
        MASTER_SALT_POR_B_i_0_i_8);
    
    \U50_PATTERNS/U3_USB_DAT_BUS/_BIBUF_F_24U[0]_/U0/U1\ : 
        IOBI_IRC_OB_EB
      port map(D => \U50_PATTERNS/WR_USB_ADBUS[0]\, CLR => 
        \AFLSDF_INV_4\, E => \U50_PATTERNS/TrienAux\, ICLK => 
        CLK60MHZ, YIN => 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[0]\\\\/U0/NET3\, 
        DOUT => 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[0]\\\\/U0/NET1\, 
        EOUT => 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[0]\\\\/U0/NET2\, 
        Y => \U50_PATTERNS/RD_USB_ADBUS[0]\);
    
    \U50_PATTERNS/U4E_REGCROSS/SAMP_ONE[0]\ : DFN1C0
      port map(D => \U50_PATTERNS/OP_MODE[0]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c, Q => 
        \U50_PATTERNS/U4E_REGCROSS/SAMP_ONE[0]_net_1\);
    
    HIEFFPLA_INST_0_45482 : AND3A
      port map(A => HIEFFPLA_NET_0_119437, B => 
        \U50_PATTERNS/WR_XFER_TYPE[0]_net_1\, C => 
        HIEFFPLA_NET_0_119367, Y => HIEFFPLA_NET_0_118905);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_22[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116450, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_15, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_22[0]\);
    
    \U_ELK5_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]\ : DFN1C0
      port map(D => \U_ELK5_CH/U_SLAVE_1ELK/Q[9]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_17[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116204, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_7, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_17[1]\);
    
    HIEFFPLA_INST_0_43165 : NAND3B
      port map(A => \U50_PATTERNS/USB_TXE_B\, B => 
        \U50_PATTERNS/REG_STATE_0[5]_net_1\, C => 
        \U50_PATTERNS/REG_STATE[4]_net_1\, Y => 
        HIEFFPLA_NET_0_119357);
    
    HIEFFPLA_INST_0_47621 : NAND2B
      port map(A => \OP_MODE_c_2[1]\, B => \PATT_ELK_DAT_14[2]\, 
        Y => HIEFFPLA_NET_0_118461);
    
    HIEFFPLA_INST_0_43108 : AND2
      port map(A => \U50_PATTERNS/REG_STATE[5]_net_1\, B => 
        HIEFFPLA_NET_0_119005, Y => HIEFFPLA_NET_0_119374);
    
    \U_ELK16_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]\ : DFN1C0
      port map(D => \U_ELK16_CH/U_SLAVE_1ELK/Q[12]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]_net_1\);
    
    HIEFFPLA_INST_0_46594 : MX2
      port map(A => 
        \U_ELK10_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]_net_1\, B => 
        \U_ELK10_CH/ELK_TX_DAT[4]\, S => 
        \U_ELK10_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118650);
    
    HIEFFPLA_INST_0_63113 : XA1C
      port map(A => HIEFFPLA_NET_0_115916, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[9]\, C => 
        HIEFFPLA_NET_0_117081, Y => HIEFFPLA_NET_0_115885);
    
    HIEFFPLA_INST_0_45362 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_19[7]\, C => 
        \U50_PATTERNS/SM_BANK_SEL[0]\, Y => HIEFFPLA_NET_0_118930);
    
    HIEFFPLA_INST_0_42794 : AOI1C
      port map(A => HIEFFPLA_NET_0_119385, B => 
        HIEFFPLA_NET_0_119463, C => HIEFFPLA_NET_0_119478, Y => 
        HIEFFPLA_NET_0_119461);
    
    HIEFFPLA_INST_0_39146 : MX2
      port map(A => HIEFFPLA_NET_0_119524, B => 
        \U50_PATTERNS/ELINK_ADDRA_18[0]\, S => 
        HIEFFPLA_NET_0_119264, Y => HIEFFPLA_NET_0_120023);
    
    \U_ELK9_CH/U_ELK1_SERDAT_SOURCE/SERDAT[5]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117828, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_7, Q => 
        \U_ELK9_CH/ELK_TX_DAT[5]\);
    
    \U50_PATTERNS/TFC_STOP_ADDR_T[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119175, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_15, Q => 
        \U50_PATTERNS/TFC_STOP_ADDR_T[5]\);
    
    HIEFFPLA_INST_0_58257 : MX2
      port map(A => HIEFFPLA_NET_0_116687, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_12[2]\, S => 
        HIEFFPLA_NET_0_117210, Y => HIEFFPLA_NET_0_116544);
    
    HIEFFPLA_INST_0_57504 : XA1B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_4[4]\, B => 
        HIEFFPLA_NET_0_116673, C => HIEFFPLA_NET_0_117179, Y => 
        HIEFFPLA_NET_0_116667);
    
    HIEFFPLA_INST_0_55762 : MX2
      port map(A => HIEFFPLA_NET_0_116995, B => 
        HIEFFPLA_NET_0_117035, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[4]\, Y => 
        HIEFFPLA_NET_0_116993);
    
    HIEFFPLA_INST_0_42345 : AND2B
      port map(A => \U50_PATTERNS/RD_USB_ADBUS[1]\, B => 
        \U50_PATTERNS/RD_USB_ADBUS[0]\, Y => 
        HIEFFPLA_NET_0_119562);
    
    HIEFFPLA_INST_0_52240 : AO1
      port map(A => HIEFFPLA_NET_0_117591, B => 
        HIEFFPLA_NET_0_117592, C => HIEFFPLA_NET_0_117179, Y => 
        HIEFFPLA_NET_0_117602);
    
    \U_ELK14_CH/U_SLAVE_1ELK/RECD_SER_WORD[7]\ : DFN1C0
      port map(D => \U_ELK14_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[7]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_14[7]\);
    
    \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[3]\ : DFN1C0
      port map(D => 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[3]_net_1\);
    
    \U50_PATTERNS/U4E_REGCROSS/LOCAL_REG_VAL[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119066, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_6, Q => \OP_MODE[4]\);
    
    HIEFFPLA_INST_0_45894 : AO1
      port map(A => HIEFFPLA_NET_0_119283, B => 
        \U50_PATTERNS/ELINK_DOUTA_13[2]\, C => 
        HIEFFPLA_NET_0_118764, Y => HIEFFPLA_NET_0_118818);
    
    HIEFFPLA_INST_0_37112 : AND3B
      port map(A => \U200A_TFC/LOC_STRT_ADDR[3]\, B => 
        HIEFFPLA_NET_0_120293, C => HIEFFPLA_NET_0_120328, Y => 
        HIEFFPLA_NET_0_120345);
    
    HIEFFPLA_INST_0_54512 : MX2
      port map(A => HIEFFPLA_NET_0_117305, B => 
        HIEFFPLA_NET_0_117286, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[2]_net_1\, Y => 
        HIEFFPLA_NET_0_117256);
    
    \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[2]\ : DFN1C0
      port map(D => \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\);
    
    HIEFFPLA_INST_0_45940 : AND3B
      port map(A => HIEFFPLA_NET_0_119426, B => 
        HIEFFPLA_NET_0_119379, C => \U50_PATTERNS/OP_MODE[6]\, Y
         => HIEFFPLA_NET_0_118806);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_28[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116053, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_15, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_28[2]\);
    
    HIEFFPLA_INST_0_55588 : MX2
      port map(A => HIEFFPLA_NET_0_116197, B => 
        HIEFFPLA_NET_0_116089, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_1[3]\, Y => 
        HIEFFPLA_NET_0_117017);
    
    HIEFFPLA_INST_0_46684 : MX2
      port map(A => \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\, 
        B => \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[11]_net_1\, S => 
        \BIT_OS_SEL_5[2]\, Y => HIEFFPLA_NET_0_118628);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_31[4]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116016, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_10, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_31[4]\);
    
    HIEFFPLA_INST_0_58595 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_17[1]\, B => 
        HIEFFPLA_NET_0_116677, S => HIEFFPLA_NET_0_117161, Y => 
        HIEFFPLA_NET_0_116500);
    
    \U_ELK7_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]\ : DFN1C0
      port map(D => \U_ELK7_CH/U_SLAVE_1ELK/Q[3]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_9[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116285, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_6, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_9[0]\);
    
    HIEFFPLA_INST_0_55192 : AND2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[6]_net_1\, B => 
        HIEFFPLA_NET_0_117336, Y => HIEFFPLA_NET_0_117098);
    
    HIEFFPLA_INST_0_50174 : MX2
      port map(A => HIEFFPLA_NET_0_117999, B => 
        HIEFFPLA_NET_0_117995, S => \BIT_OS_SEL_6[1]\, Y => 
        HIEFFPLA_NET_0_117997);
    
    HIEFFPLA_INST_0_41999 : AO1A
      port map(A => HIEFFPLA_NET_0_119629, B => 
        HIEFFPLA_NET_0_118693, C => HIEFFPLA_NET_0_119634, Y => 
        HIEFFPLA_NET_0_119635);
    
    HIEFFPLA_INST_0_113940 : AO18
      port map(A => HIEFFPLA_NET_0_115809, B => \ELKS_ADDRB[2]\, 
        C => \U200B_ELINKS/LOC_STOP_ADDR[2]\, Y => 
        HIEFFPLA_NET_0_115813);
    
    HIEFFPLA_INST_0_56303 : NAND3C
      port map(A => HIEFFPLA_NET_0_116873, B => 
        HIEFFPLA_NET_0_116881, C => HIEFFPLA_NET_0_116889, Y => 
        HIEFFPLA_NET_0_116897);
    
    HIEFFPLA_INST_0_50768 : MX2
      port map(A => HIEFFPLA_NET_0_117905, B => 
        HIEFFPLA_NET_0_117915, S => \BIT_OS_SEL_5[0]\, Y => 
        \U_ELK7_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[5]\);
    
    HIEFFPLA_INST_0_48254 : MX2
      port map(A => HIEFFPLA_NET_0_118352, B => 
        HIEFFPLA_NET_0_118350, S => \BIT_OS_SEL_3[0]\, Y => 
        \U_ELK16_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[2]\);
    
    \U_ELK14_CH/ELK_IN_F\ : DFN1C0
      port map(D => \U_ELK14_CH/ELK_IN_DDR_F\, CLK => 
        CCC_160M_ADJ, CLR => DEV_RST_B_c, Q => 
        \U_ELK14_CH/ELK_IN_F_net_1\);
    
    \U200B_ELINKS/GP_PG_SM[9]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120205, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_29, Q => 
        \U200B_ELINKS/GP_PG_SM[9]_net_1\);
    
    HIEFFPLA_INST_0_50662 : MX2
      port map(A => \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[3]_net_1\, B
         => \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\, S => 
        \BIT_OS_SEL_4[2]\, Y => HIEFFPLA_NET_0_117909);
    
    HIEFFPLA_INST_0_46431 : NAND3B
      port map(A => HIEFFPLA_NET_0_119452, B => 
        HIEFFPLA_NET_0_118690, C => HIEFFPLA_NET_0_119020, Y => 
        HIEFFPLA_NET_0_118691);
    
    HIEFFPLA_INST_0_45188 : NAND3C
      port map(A => HIEFFPLA_NET_0_118797, B => 
        HIEFFPLA_NET_0_118874, C => HIEFFPLA_NET_0_118960, Y => 
        HIEFFPLA_NET_0_118969);
    
    \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[11]\ : DFN1C0
      port map(D => 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]_net_1\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[11]_net_1\);
    
    \U50_PATTERNS/REG_ADDR[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119531, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_10, Q => \U50_PATTERNS/REG_ADDR[2]\);
    
    HIEFFPLA_INST_0_52550 : MX2
      port map(A => HIEFFPLA_NET_0_117489, B => 
        HIEFFPLA_NET_0_117485, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_2[3]\, Y => 
        HIEFFPLA_NET_0_117549);
    
    HIEFFPLA_INST_0_41858 : OA1A
      port map(A => HIEFFPLA_NET_0_119231, B => 
        \U50_PATTERNS/ELINK_RWA[18]\, C => HIEFFPLA_NET_0_119651, 
        Y => HIEFFPLA_NET_0_119681);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_2[6]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116749, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_5, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_2[6]\);
    
    \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[14]\ : DFN1C0
      port map(D => \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\, 
        CLK => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[14]_net_1\);
    
    \U50_PATTERNS/ELINK_RWA[16]/U1\ : DFN1P0
      port map(D => HIEFFPLA_NET_0_119704, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_12, Q => 
        \U50_PATTERNS/ELINK_RWA[16]\);
    
    HIEFFPLA_INST_0_37578 : AND3
      port map(A => HIEFFPLA_NET_0_120258, B => \TFC_ADDRB[5]\, C
         => \TFC_ADDRB[4]\, Y => HIEFFPLA_NET_0_120256);
    
    HIEFFPLA_INST_0_56221 : AND3A
      port map(A => \ELK_RX_SER_WORD_0[0]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/RECD_SER_WORD[2]_net_1\, 
        C => 
        \U_MASTER_DES/U13C_MASTER_DESER/RECD_SER_WORD[1]_net_1\, 
        Y => HIEFFPLA_NET_0_116927);
    
    \U50_PATTERNS/SM_BANK_SEL[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119305, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_7, Q => 
        \U50_PATTERNS/SM_BANK_SEL[5]\);
    
    HIEFFPLA_INST_0_47704 : MX2
      port map(A => \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\, 
        B => \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[12]_net_1\, S => 
        \BIT_OS_SEL_2[2]\, Y => HIEFFPLA_NET_0_118444);
    
    \U_ELK10_CH/U_SLAVE_1ELK/Q[3]\ : DFN1C0
      port map(D => \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/Q[3]_net_1\);
    
    AFLSDF_INV_54 : INV
      port map(A => \U200A_TFC/RX_SER_WORD_2DEL[3]_net_1\, Y => 
        \AFLSDF_INV_54\);
    
    \U_ELK7_CH/U_ELK1_SERDAT_SOURCE/SERDAT[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117921, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_3, Q => 
        \U_ELK7_CH/ELK_TX_DAT[2]\);
    
    \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[9]\ : DFN1C0
      port map(D => \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\);
    
    HIEFFPLA_INST_0_60774 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_31[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_15[1]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[4]_net_1\, Y
         => HIEFFPLA_NET_0_116222);
    
    HIEFFPLA_INST_0_57788 : NAND3
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_6[0]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_6[2]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_6[1]\, Y => 
        HIEFFPLA_NET_0_116623);
    
    HIEFFPLA_INST_0_43685 : AND2A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/SM_BANK_SEL[18]\, Y => 
        HIEFFPLA_NET_0_119241);
    
    \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[13]\ : DFN1C0
      port map(D => 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[13]_net_1\);
    
    \U_ELK5_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]\ : DFN1C0
      port map(D => \U_ELK5_CH/U_SLAVE_1ELK/Q[0]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]_net_1\);
    
    HIEFFPLA_INST_0_59139 : MX2
      port map(A => HIEFFPLA_NET_0_116426, B => 
        HIEFFPLA_NET_0_116423, S => HIEFFPLA_NET_0_117249, Y => 
        HIEFFPLA_NET_0_116430);
    
    HIEFFPLA_INST_0_51585 : AX1C
      port map(A => HIEFFPLA_NET_0_117747, B => 
        HIEFFPLA_NET_0_117753, C => HIEFFPLA_NET_0_117733, Y => 
        HIEFFPLA_NET_0_117739);
    
    HIEFFPLA_INST_0_51076 : MX2
      port map(A => 
        \U_ELK9_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]_net_1\, B => 
        \U_ELK9_CH/ELK_TX_DAT[4]\, S => 
        \U_ELK9_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_117840);
    
    HIEFFPLA_INST_0_51722 : NAND2B
      port map(A => 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM_0[4]_net_1\, B => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[77]_net_1\, Y => 
        HIEFFPLA_NET_0_117704);
    
    \U200B_ELINKS/ADDR_POINTER[4]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120164, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_32, Q => \ELKS_ADDRB[4]\);
    
    \U50_PATTERNS/ELINK_ADDRA_11[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120078, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_2, Q => 
        \U50_PATTERNS/ELINK_ADDRA_11[1]\);
    
    HIEFFPLA_INST_0_48331 : MX2
      port map(A => 
        \U_ELK17_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]_net_1\, B => 
        \U_ELK17_CH/ELK_TX_DAT[2]\, S => 
        \U_ELK17_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118336);
    
    HIEFFPLA_INST_0_40079 : AOI1D
      port map(A => HIEFFPLA_NET_0_119389, B => 
        HIEFFPLA_NET_0_119464, C => 
        \U50_PATTERNS/SM_BANK_SEL[19]\, Y => 
        HIEFFPLA_NET_0_119914);
    
    \U_ELK1_CH/U_ELK1_SERDAT_SOURCE/SERDAT[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118193, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_11, Q => 
        \U_ELK1_CH/ELK_TX_DAT[0]\);
    
    HIEFFPLA_INST_0_46009 : AND3B
      port map(A => HIEFFPLA_NET_0_119426, B => 
        HIEFFPLA_NET_0_119379, C => \U50_PATTERNS/OP_MODE[7]\, Y
         => HIEFFPLA_NET_0_118788);
    
    \U_ELK10_CH/U_SLAVE_1ELK/RECD_SER_WORD[5]\ : DFN1C0
      port map(D => \U_ELK10_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[5]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_10[5]\);
    
    \U50_PATTERNS/SM_BANK_SEL[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119322, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_7, Q => 
        \U50_PATTERNS/SM_BANK_SEL[0]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/Q[10]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[10]_net_1\, CLK => 
        CCC_160M_FXD, CLR => P_MASTER_POR_B_c_23, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/Q[10]_net_1\);
    
    HIEFFPLA_INST_0_57145 : XA1B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_2[4]\, B => 
        HIEFFPLA_NET_0_116743, C => HIEFFPLA_NET_0_117179, Y => 
        HIEFFPLA_NET_0_116731);
    
    HIEFFPLA_INST_0_44649 : XOR2
      port map(A => \ELKS_STOP_ADDR[7]\, B => 
        \U50_PATTERNS/U4D_REGCROSS/SAMP_TWO[7]_net_1\, Y => 
        HIEFFPLA_NET_0_119074);
    
    HIEFFPLA_INST_0_46534 : AND3A
      port map(A => \U50_PATTERNS/REG_STATE_0[2]_net_1\, B => 
        \U50_PATTERNS/REG_STATE[4]_net_1\, C => 
        HIEFFPLA_NET_0_119367, Y => HIEFFPLA_NET_0_118670);
    
    \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[1]\ : DFN1C0
      port map(D => 
        \U_ELK18_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_6[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116632, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_12, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_6[0]\);
    
    \U_ELK6_CH/U_SLAVE_1ELK/Q[1]\ : DFN1C0
      port map(D => \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/Q[1]_net_1\);
    
    \U50_PATTERNS/ELINK_RWA[11]/U1\ : DFN1P0
      port map(D => HIEFFPLA_NET_0_119709, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_11, Q => 
        \U50_PATTERNS/ELINK_RWA[11]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_15[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116230, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_4, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_15[0]\);
    
    HIEFFPLA_INST_0_42885 : NAND3C
      port map(A => \U50_PATTERNS/REG_STATE[1]_net_1\, B => 
        \U50_PATTERNS/REG_STATE[3]_net_1\, C => 
        \U50_PATTERNS/REG_STATE[4]_net_1\, Y => 
        HIEFFPLA_NET_0_119436);
    
    \U50_PATTERNS/ELINK_DINA_5[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119744, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_14, Q => 
        \U50_PATTERNS/ELINK_DINA_5[7]\);
    
    \U50_PATTERNS/RD_XFER_TYPE[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119547, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c, Q => 
        \U50_PATTERNS/RD_XFER_TYPE[2]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_6[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116630, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_12, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_6[2]\);
    
    HIEFFPLA_INST_0_57692 : AOI1A
      port map(A => HIEFFPLA_NET_0_116647, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_5[4]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_5[5]\, Y => 
        HIEFFPLA_NET_0_116634);
    
    HIEFFPLA_INST_0_44537 : XOR2
      port map(A => \ELKS_STRT_ADDR[3]\, B => 
        \U50_PATTERNS/U4C_REGCROSS/SAMP_TWO[3]_net_1\, Y => 
        HIEFFPLA_NET_0_119098);
    
    HIEFFPLA_INST_0_48979 : MX2
      port map(A => \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\, 
        B => \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\, S => 
        \BIT_OS_SEL[2]\, Y => HIEFFPLA_NET_0_118215);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_28[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116054, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_15, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_28[1]\);
    
    \U50_PATTERNS/OP_MODE[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119610, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_15, Q => \U50_PATTERNS/OP_MODE[7]\);
    
    HIEFFPLA_INST_0_57267 : NAND3A
      port map(A => HIEFFPLA_NET_0_116711, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_3[4]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_3[5]\, Y => 
        HIEFFPLA_NET_0_116712);
    
    HIEFFPLA_INST_0_50005 : MX2
      port map(A => HIEFFPLA_NET_0_118049, B => 
        HIEFFPLA_NET_0_118043, S => \BIT_OS_SEL_0[0]\, Y => 
        \U_ELK4_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[3]\);
    
    HIEFFPLA_INST_0_41911 : AND2A
      port map(A => \U50_PATTERNS/ELINK_RWA[0]\, B => 
        HIEFFPLA_NET_0_119664, Y => HIEFFPLA_NET_0_119665);
    
    \U_ELK4_CH/U_ELK1_CMD_TX/SER_OUT_FI\ : DFI1C0
      port map(D => 
        \U_ELK4_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_4, QN
         => \U_ELK4_CH/U_ELK1_CMD_TX/SER_OUT_FI_i\);
    
    \U_GEN_REF_CLK/GEN_40M_REF\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117728, CLK => Y, CLR => 
        DEV_RST_B_c, Q => CLK40M_10NS_REF);
    
    \U_ELK2_CH/U_SLAVE_1ELK/RECD_SER_WORD[0]\ : DFN1C0
      port map(D => \U_ELK2_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[0]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_2[0]\);
    
    \U50_PATTERNS/TFC_DINA[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119194, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_4, Q => \U50_PATTERNS/TFC_DINA[3]\);
    
    HIEFFPLA_INST_0_60357 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_9[3]\, B => 
        HIEFFPLA_NET_0_116815, S => HIEFFPLA_NET_0_117393, Y => 
        HIEFFPLA_NET_0_116276);
    
    HIEFFPLA_INST_0_53801 : AND3
      port map(A => HIEFFPLA_NET_0_117135, B => 
        HIEFFPLA_NET_0_117334, C => HIEFFPLA_NET_0_117325, Y => 
        HIEFFPLA_NET_0_117350);
    
    HIEFFPLA_INST_0_51501 : NAND2B
      port map(A => \U_EXEC_MASTER/PRESCALE[2]\, B => 
        \U_EXEC_MASTER/PRESCALE[3]\, Y => HIEFFPLA_NET_0_117763);
    
    \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[9]\ : DFN1C0
      port map(D => 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\);
    
    \U_ELK16_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]\ : DFN1C0
      port map(D => \U_ELK16_CH/U_SLAVE_1ELK/Q[14]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]_net_1\);
    
    HIEFFPLA_INST_0_55572 : MX2
      port map(A => HIEFFPLA_NET_0_116163, B => 
        HIEFFPLA_NET_0_116268, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_1[3]\, Y => 
        HIEFFPLA_NET_0_117019);
    
    \U50_PATTERNS/U3_USB_DAT_BUS/_BIBUF_F_24U[6]_/U0/U1\ : 
        IOBI_IRC_OB_EB
      port map(D => \U50_PATTERNS/WR_USB_ADBUS[6]\, CLR => 
        \AFLSDF_INV_10\, E => \U50_PATTERNS/TrienAux\, ICLK => 
        CLK60MHZ, YIN => 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[6]\\\\/U0/NET3\, 
        DOUT => 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[6]\\\\/U0/NET1\, 
        EOUT => 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[6]\\\\/U0/NET2\, 
        Y => \U50_PATTERNS/RD_USB_ADBUS[6]\);
    
    HIEFFPLA_INST_0_46003 : AND3B
      port map(A => HIEFFPLA_NET_0_119426, B => 
        HIEFFPLA_NET_0_119379, C => \U50_PATTERNS/OP_MODE[4]\, Y
         => HIEFFPLA_NET_0_118790);
    
    HIEFFPLA_INST_0_49327 : MX2
      port map(A => 
        \U_ELK2_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]_net_1\, B => 
        \U_ELK2_CH/ELK_TX_DAT[2]\, S => 
        \U_ELK2_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118156);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_22[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116130, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_5, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_22[0]\);
    
    HIEFFPLA_INST_0_45100 : MX2
      port map(A => HIEFFPLA_NET_0_118974, B => 
        \U50_PATTERNS/WR_USB_ADBUS[2]\, S => 
        HIEFFPLA_NET_0_119486, Y => HIEFFPLA_NET_0_118983);
    
    \U_ELK8_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117887, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_3[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116722, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_7, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_3[3]\);
    
    AFLSDF_INV_48 : INV
      port map(A => DCB_SALT_SEL_c, Y => \AFLSDF_INV_48\);
    
    HIEFFPLA_INST_0_40630 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_14[4]\, B => 
        HIEFFPLA_NET_0_119570, S => HIEFFPLA_NET_0_119249, Y => 
        HIEFFPLA_NET_0_119827);
    
    \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[72]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117707, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_33, Q => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[72]_net_1\);
    
    \U_EXEC_MASTER/USB_MASTER_EN/TEST_SM[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117752, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_24, Q => 
        \U_EXEC_MASTER/USB_MASTER_EN/TEST_SM[1]_net_1\);
    
    HIEFFPLA_INST_0_48146 : MX2
      port map(A => \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\, 
        B => \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\, S => 
        \BIT_OS_SEL_1[2]\, Y => HIEFFPLA_NET_0_118362);
    
    \U50_PATTERNS/U4E_REGCROSS/SAMP_ONE[5]\ : DFN1C0
      port map(D => \U50_PATTERNS/OP_MODE[5]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c, Q => 
        \U50_PATTERNS/U4E_REGCROSS/SAMP_ONE[5]_net_1\);
    
    HIEFFPLA_INST_0_43574 : AND2A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/SM_BANK_SEL[6]\, Y => HIEFFPLA_NET_0_119283);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_23[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116120, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_6, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_23[0]\);
    
    HIEFFPLA_INST_0_58476 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_15[3]\, B => 
        HIEFFPLA_NET_0_116815, S => HIEFFPLA_NET_0_117098, Y => 
        HIEFFPLA_NET_0_116517);
    
    HIEFFPLA_INST_0_49078 : MX2
      port map(A => 
        \U_ELK1_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]_net_1\, B => 
        \U_ELK1_CH/ELK_TX_DAT[2]\, S => 
        \U_ELK1_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118201);
    
    \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[14]\ : DFN1C0
      port map(D => 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]_net_1\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[14]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117045, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_16_0, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[0]\);
    
    HIEFFPLA_INST_0_58948 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_21[1]\, B => 
        HIEFFPLA_NET_0_116677, S => HIEFFPLA_NET_0_117093, Y => 
        HIEFFPLA_NET_0_116455);
    
    HIEFFPLA_INST_0_42531 : OA1A
      port map(A => HIEFFPLA_NET_0_119433, B => 
        HIEFFPLA_NET_0_119010, C => \U50_PATTERNS/REG_ADDR[4]\, Y
         => HIEFFPLA_NET_0_119519);
    
    \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[4]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_115935, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_24_0, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[4]_net_1\);
    
    \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[0]\ : DFN1C0
      port map(D => 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[0]_net_1\);
    
    HIEFFPLA_INST_0_49435 : MX2
      port map(A => \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\, B
         => \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\, S => 
        \BIT_OS_SEL_7[2]\, Y => HIEFFPLA_NET_0_118131);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_20[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116160, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_2, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_20[0]\);
    
    \U_ELK5_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118015, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_2, Q => 
        \U_ELK5_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]_net_1\);
    
    \U_EXEC_MASTER/MPOR_B_18\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117787, CLK => CLK_40M_GL, CLR
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_1\, Q => 
        P_MASTER_POR_B_c_18);
    
    HIEFFPLA_INST_0_45589 : AO1A
      port map(A => HIEFFPLA_NET_0_119622, B => 
        \U50_PATTERNS/TFC_STOP_ADDR[4]\, C => 
        HIEFFPLA_NET_0_118777, Y => HIEFFPLA_NET_0_118885);
    
    \U_MASTER_DES/U13C_MASTER_DESER/MAX_CNT[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_116953, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_16, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/MAX_CNT[1]\);
    
    \U_ELK9_CH/U_SLAVE_1ELK/RECD_SER_WORD[1]\ : DFN1C0
      port map(D => \U_ELK9_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[1]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_9[1]\);
    
    \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[4]\ : DFN1C0
      port map(D => 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\);
    
    HIEFFPLA_INST_0_48457 : MX2
      port map(A => HIEFFPLA_NET_0_118312, B => 
        HIEFFPLA_NET_0_118309, S => \BIT_OS_SEL_1[1]\, Y => 
        HIEFFPLA_NET_0_118308);
    
    HIEFFPLA_INST_0_47507 : MX2
      port map(A => HIEFFPLA_NET_0_118490, B => 
        HIEFFPLA_NET_0_118486, S => \BIT_OS_SEL_4[0]\, Y => 
        \U_ELK13_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[2]\);
    
    HIEFFPLA_INST_0_56731 : NAND3B
      port map(A => HIEFFPLA_NET_0_116800, B => 
        HIEFFPLA_NET_0_116808, C => HIEFFPLA_NET_0_116802, Y => 
        HIEFFPLA_NET_0_116813);
    
    HIEFFPLA_INST_0_57533 : AXOI4
      port map(A => HIEFFPLA_NET_0_117085, B => 
        HIEFFPLA_NET_0_117121, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_5[0]\, Y => 
        HIEFFPLA_NET_0_116661);
    
    HIEFFPLA_INST_0_51678 : MX2
      port map(A => \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[46]\, B
         => \U_MASTER_DES/PHASE_ADJ_160_L[0]\, S => 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM_0[4]_net_1\, Y => 
        HIEFFPLA_NET_0_117726);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_27[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116070, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_13, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_27[0]\);
    
    \U200B_ELINKS/GP_PG_SM[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120213, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_29, Q => 
        \U200B_ELINKS/GP_PG_SM[3]_net_1\);
    
    HIEFFPLA_INST_0_52678 : MX2
      port map(A => HIEFFPLA_NET_0_117480, B => 
        HIEFFPLA_NET_0_117476, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[4]\, Y => 
        HIEFFPLA_NET_0_117528);
    
    \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[5]\ : DFN1C0
      port map(D => \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\);
    
    HIEFFPLA_INST_0_57434 : NAND3C
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_4[7]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_4[6]\, C => 
        HIEFFPLA_NET_0_116674, Y => HIEFFPLA_NET_0_116685);
    
    HIEFFPLA_INST_0_51365 : MX2
      port map(A => HIEFFPLA_NET_0_117774, B => 
        \U_EXEC_MASTER/DEL_CNT[4]\, S => HIEFFPLA_NET_0_117796, Y
         => HIEFFPLA_NET_0_117791);
    
    HIEFFPLA_INST_0_58275 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_13[0]\, B => 
        HIEFFPLA_NET_0_116538, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_0[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116542);
    
    \U200B_ELINKS/R_BLKB/U1\ : DFN1P0
      port map(D => HIEFFPLA_NET_0_120154, CLK => CLK_40M_GL, PRE
         => P_MASTER_POR_B_c_13, Q => ELKS_RAM_BLKB_EN);
    
    HIEFFPLA_INST_0_59111 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_24[0]\, B => 
        HIEFFPLA_NET_0_116430, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_2[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116434);
    
    HIEFFPLA_INST_0_51554 : AND3
      port map(A => HIEFFPLA_NET_0_117744, B => 
        \U_EXEC_MASTER/USB_MASTER_EN/T_CNT60M[7]_net_1\, C => 
        \U_EXEC_MASTER/USB_MASTER_EN/T_CNT60M[4]_net_1\, Y => 
        HIEFFPLA_NET_0_117745);
    
    \U_ELK16_CH/ELK_IN_F\ : DFN1C0
      port map(D => \U_ELK16_CH/ELK_IN_DDR_F\, CLK => 
        CCC_160M_ADJ, CLR => DEV_RST_B_c, Q => 
        \U_ELK16_CH/ELK_IN_F_net_1\);
    
    \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[7]\ : DFN1C0
      port map(D => \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_1[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117022, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_17_0, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_1[3]\);
    
    \U_ELK1_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118199, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_7, Q => 
        \U_ELK1_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]_net_1\);
    
    \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[4]\ : DFN1C0
      port map(D => \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\);
    
    HIEFFPLA_INST_0_55310 : AND3B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[0]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[2]_net_1\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[3]_net_1\, Y => 
        HIEFFPLA_NET_0_117064);
    
    HIEFFPLA_INST_0_42026 : NAND2B
      port map(A => \U50_PATTERNS/ELK_N_ACTIVE_net_1\, B => 
        \U50_PATTERNS/REG_STATE_0[5]_net_1\, Y => 
        HIEFFPLA_NET_0_119629);
    
    HIEFFPLA_INST_0_37591 : AO1A
      port map(A => \ELKS_STRT_ADDR[1]\, B => 
        HIEFFPLA_NET_0_120219, C => HIEFFPLA_NET_0_120242, Y => 
        HIEFFPLA_NET_0_120252);
    
    HIEFFPLA_INST_0_40963 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_19[1]\, B => 
        HIEFFPLA_NET_0_119576, S => HIEFFPLA_NET_0_119293, Y => 
        HIEFFPLA_NET_0_119790);
    
    \U_ELK5_CH/U_ELK1_SERDAT_SOURCE/SERDAT[6]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118007, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i, Q => 
        \U_ELK5_CH/ELK_TX_DAT[6]\);
    
    \U_ELK12_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL\ : DFN1C0
      port map(D => 
        \U_ELK12_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL_net_1\);
    
    \U_ELK10_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]\ : DFN1C0
      port map(D => \U_ELK10_CH/U_SLAVE_1ELK/Q[0]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]_net_1\);
    
    \U_ELK4_CH/U_ELK1_SERDAT_SOURCE/SERDAT[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118056, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_16, Q => 
        \U_ELK4_CH/ELK_TX_DAT[2]\);
    
    \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[11]\ : DFN1C0
      port map(D => \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\);
    
    HIEFFPLA_INST_0_49674 : MX2
      port map(A => \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\, B
         => \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[11]_net_1\, S => 
        \BIT_OS_SEL_7[2]\, Y => HIEFFPLA_NET_0_118087);
    
    HIEFFPLA_INST_0_45942 : AND3A
      port map(A => HIEFFPLA_NET_0_119376, B => 
        \U50_PATTERNS/TFC_STRT_ADDR[7]\, C => 
        HIEFFPLA_NET_0_119431, Y => HIEFFPLA_NET_0_118805);
    
    \U50_PATTERNS/U4B_REGCROSS/LOCAL_REG_VAL[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119130, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_19, Q => \TFC_STOP_ADDR[3]\);
    
    \U_ELK17_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U3\ : IOBI_ID_OD_EB
      port map(DR => \U_ELK17_CH/ELK_OUT_R\, DF => 
        \U_ELK17_CH/ELK_OUT_F\, CLR => \GND\, E => 
        \AFLSDF_INV_29\, ICLK => CCC_160M_ADJ, OCLK => 
        CCC_160M_FXD, YIN => 
        \U_ELK17_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\, DOUT => 
        OPEN, EOUT => 
        \U_ELK17_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET3\, YR => OPEN, 
        YF => OPEN);
    
    \U50_PATTERNS/ELINK_DINA_15[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119818, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_16, Q => 
        \U50_PATTERNS/ELINK_DINA_15[5]\);
    
    HIEFFPLA_INST_0_38498 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_0[0]\, B => 
        HIEFFPLA_NET_0_119524, S => HIEFFPLA_NET_0_119272, Y => 
        HIEFFPLA_NET_0_120095);
    
    \U_ELK19_CH/U_SLAVE_1ELK/RECD_SER_WORD[5]\ : DFN1C0
      port map(D => \U_ELK19_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[5]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_19[5]\);
    
    HIEFFPLA_INST_0_55734 : AND3B
      port map(A => HIEFFPLA_NET_0_117185, B => 
        HIEFFPLA_NET_0_117087, C => HIEFFPLA_NET_0_117027, Y => 
        HIEFFPLA_NET_0_116997);
    
    HIEFFPLA_INST_0_47105 : MX2
      port map(A => 
        \U_ELK12_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]_net_1\, B => 
        \U_ELK12_CH/ELK_TX_DAT[3]\, S => 
        \U_ELK12_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118557);
    
    \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[8]\ : DFN1C0
      port map(D => 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\);
    
    \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[1]\ : DFN1C0
      port map(D => 
        \U_ELK7_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\);
    
    \U_ELK18_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118287, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_0, Q => 
        \U_ELK18_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]_net_1\);
    
    HIEFFPLA_INST_0_44086 : MX2
      port map(A => \U50_PATTERNS/TFC_STOP_ADDR_T[5]\, B => 
        \U50_PATTERNS/RD_USB_ADBUS[5]\, S => 
        HIEFFPLA_NET_0_119492, Y => HIEFFPLA_NET_0_119175);
    
    HIEFFPLA_INST_0_111335 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_25[0]\, B => 
        HIEFFPLA_NET_0_116735, S => HIEFFPLA_NET_0_117394, Y => 
        HIEFFPLA_NET_0_116409);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_20[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116159, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_2, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_20[1]\);
    
    \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[12]\ : DFN1C0
      port map(D => \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\, 
        CLK => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\);
    
    HIEFFPLA_INST_0_52666 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_17[2]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_18[2]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_3[0]\, Y => 
        HIEFFPLA_NET_0_117530);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_4[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_115997, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_13, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_4[3]\);
    
    \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[3]\ : DFN1C0
      port map(D => \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\);
    
    HIEFFPLA_INST_0_41368 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_5[6]\, B => 
        HIEFFPLA_NET_0_119566, S => HIEFFPLA_NET_0_119251, Y => 
        HIEFFPLA_NET_0_119745);
    
    HIEFFPLA_INST_0_48238 : MX2
      port map(A => HIEFFPLA_NET_0_118341, B => 
        HIEFFPLA_NET_0_118356, S => \BIT_OS_SEL_3[0]\, Y => 
        \U_ELK16_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[0]\);
    
    \U50_PATTERNS/ELINKS_STOP_ADDR[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120127, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_14, Q => 
        \U50_PATTERNS/ELINKS_STOP_ADDR[0]\);
    
    HIEFFPLA_INST_0_47580 : AND2
      port map(A => \U_ELK14_CH/ELK_TX_DAT[0]\, B => 
        \U_ELK14_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118472);
    
    \U200B_ELINKS/RX_SER_WORD_1DEL[4]\ : DFN1C0
      port map(D => \ELK_RX_SER_WORD_0[4]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_23, Q => 
        \U200B_ELINKS/RX_SER_WORD_1DEL[4]_net_1\);
    
    HIEFFPLA_INST_0_52140 : AND3C
      port map(A => 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM_0[4]_net_1\, B => 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM[3]_net_1\, C => 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM[5]_net_1\, Y => 
        HIEFFPLA_NET_0_117628);
    
    HIEFFPLA_INST_0_48370 : AND2A
      port map(A => \OP_MODE_c_6[1]\, B => \PATT_ELK_DAT_17[4]\, 
        Y => HIEFFPLA_NET_0_118324);
    
    HIEFFPLA_INST_0_55580 : MX2
      port map(A => HIEFFPLA_NET_0_116162, B => 
        HIEFFPLA_NET_0_116267, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_1[3]\, Y => 
        HIEFFPLA_NET_0_117018);
    
    HIEFFPLA_INST_0_51402 : NAND2A
      port map(A => HIEFFPLA_NET_0_117782, B => 
        \U_EXEC_MASTER/DEL_CNT[4]\, Y => HIEFFPLA_NET_0_117785);
    
    HIEFFPLA_INST_0_47017 : MX2
      port map(A => HIEFFPLA_NET_0_118579, B => 
        HIEFFPLA_NET_0_118576, S => \BIT_OS_SEL[0]\, Y => 
        \U_ELK11_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[3]\);
    
    \U_ELK4_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]\ : DFN1C0
      port map(D => \U_ELK4_CH/U_SLAVE_1ELK/Q[5]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]_net_1\);
    
    \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[10]\ : DFN1C0
      port map(D => \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\);
    
    \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[6]\ : DFN1C0
      port map(D => 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\);
    
    HIEFFPLA_INST_0_63227 : MX2
      port map(A => \U_TFC_CMD_TX/SER_CMD_WORD_R[1]_net_1\, B => 
        \TFC_TX_DAT[5]\, S => \U_TFC_CMD_TX/START_RISE_net_1\, Y
         => \U_TFC_CMD_TX/N_SER_CMD_WORD_R[2]\);
    
    HIEFFPLA_INST_0_40148 : AOI1C
      port map(A => \U50_PATTERNS/ELINK_BLKA[4]\, B => 
        HIEFFPLA_NET_0_119643, C => HIEFFPLA_NET_0_119889, Y => 
        HIEFFPLA_NET_0_119890);
    
    HIEFFPLA_INST_0_56045 : MX2
      port map(A => HIEFFPLA_NET_0_116970, B => 
        HIEFFPLA_NET_0_116962, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[1]\, Y => 
        HIEFFPLA_NET_0_116957);
    
    HIEFFPLA_INST_0_53973 : MX2
      port map(A => HIEFFPLA_NET_0_117382, B => 
        HIEFFPLA_NET_0_117312, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[0]_net_1\, Y
         => HIEFFPLA_NET_0_117325);
    
    HIEFFPLA_INST_0_47393 : MX2
      port map(A => HIEFFPLA_NET_0_118497, B => 
        HIEFFPLA_NET_0_118493, S => \BIT_OS_SEL_3[1]\, Y => 
        HIEFFPLA_NET_0_118498);
    
    HIEFFPLA_INST_0_54676 : MX2
      port map(A => HIEFFPLA_NET_0_117233, B => 
        HIEFFPLA_NET_0_117412, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[1]_net_1\, Y => 
        HIEFFPLA_NET_0_117224);
    
    HIEFFPLA_INST_0_56254 : AND3
      port map(A => HIEFFPLA_NET_0_116924, B => 
        HIEFFPLA_NET_0_116905, C => \TFC_RX_SER_WORD[7]\, Y => 
        HIEFFPLA_NET_0_116906);
    
    \U_ELK12_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]\ : DFN1C0
      port map(D => \U_ELK12_CH/U_SLAVE_1ELK/Q[3]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]_net_1\);
    
    HIEFFPLA_INST_0_52365 : AND2A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[8]_net_1\, B => 
        HIEFFPLA_NET_0_117569, Y => HIEFFPLA_NET_0_117573);
    
    \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[9]\ : DFN1C0
      port map(D => 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\);
    
    \U_ELK10_CH/U_SLAVE_1ELK/Q[12]\ : DFN1C0
      port map(D => \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/Q[12]_net_1\);
    
    \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[5]\\\\/U0/U0\ : 
        IOPAD_BI_U
      port map(D => 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[5]\\\\/U0/NET1\, 
        E => 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[5]\\\\/U0/NET2\, 
        Y => 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[5]\\\\/U0/NET3\, 
        PAD => BIDIR_USB_ADBUS(5));
    
    HIEFFPLA_INST_0_54596 : AND3A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[2]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[4]_net_1\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[1]_net_1\, Y => 
        HIEFFPLA_NET_0_117236);
    
    HIEFFPLA_INST_0_54592 : NAND3A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[4]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[2]_net_1\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[1]_net_1\, Y => 
        HIEFFPLA_NET_0_117238);
    
    HIEFFPLA_INST_0_49981 : MX2
      port map(A => HIEFFPLA_NET_0_118026, B => 
        HIEFFPLA_NET_0_118038, S => \BIT_OS_SEL_0[0]\, Y => 
        \U_ELK4_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[0]\);
    
    HIEFFPLA_INST_0_45289 : AO1
      port map(A => HIEFFPLA_NET_0_119244, B => 
        \U50_PATTERNS/ELINK_DOUTA_2[0]\, C => 
        HIEFFPLA_NET_0_118949, Y => HIEFFPLA_NET_0_118950);
    
    HIEFFPLA_INST_0_42704 : AO1C
      port map(A => \U50_PATTERNS/REG_STATE[0]_net_1\, B => 
        \U50_PATTERNS/REG_STATE[1]_net_1\, C => 
        \U50_PATTERNS/REG_STATE_0[2]_net_1\, Y => 
        HIEFFPLA_NET_0_119479);
    
    HIEFFPLA_INST_0_111191 : NAND3
      port map(A => HIEFFPLA_NET_0_115918, B => 
        HIEFFPLA_NET_0_115915, C => HIEFFPLA_NET_0_115913, Y => 
        HIEFFPLA_NET_0_115848);
    
    HIEFFPLA_INST_0_59387 : AO1
      port map(A => HIEFFPLA_NET_0_116620, B => 
        HIEFFPLA_NET_0_117411, C => HIEFFPLA_NET_0_116589, Y => 
        HIEFFPLA_NET_0_116398);
    
    HIEFFPLA_INST_0_46357 : NAND3C
      port map(A => HIEFFPLA_NET_0_118856, B => 
        HIEFFPLA_NET_0_118862, C => HIEFFPLA_NET_0_118866, Y => 
        HIEFFPLA_NET_0_118708);
    
    HIEFFPLA_INST_0_45999 : AND3B
      port map(A => HIEFFPLA_NET_0_119426, B => 
        HIEFFPLA_NET_0_119379, C => \U50_PATTERNS/OP_MODE[2]\, Y
         => HIEFFPLA_NET_0_118792);
    
    \U_TFC_SERDAT_SOURCE/SERDAT[7]\ : DFN1C0
      port map(D => \U_TFC_SERDAT_SOURCE/N_SERDAT[7]\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \TFC_TX_DAT[7]\);
    
    HIEFFPLA_INST_0_52788 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_11[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_12[1]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_1[0]\, Y => 
        HIEFFPLA_NET_0_117511);
    
    HIEFFPLA_INST_0_42041 : AND3
      port map(A => \U50_PATTERNS/TFC_DOUTA[3]\, B => 
        HIEFFPLA_NET_0_118997, C => HIEFFPLA_NET_0_119365, Y => 
        HIEFFPLA_NET_0_119625);
    
    HIEFFPLA_INST_0_41681 : MX2
      port map(A => HIEFFPLA_NET_0_119690, B => 
        \U50_PATTERNS/ELINK_RWA[10]\, S => 
        \U50_PATTERNS/SM_BANK_SEL_0[20]\, Y => 
        HIEFFPLA_NET_0_119710);
    
    HIEFFPLA_INST_0_40567 : MX2
      port map(A => HIEFFPLA_NET_0_119567, B => 
        \U50_PATTERNS/ELINK_DINA_13[5]\, S => 
        HIEFFPLA_NET_0_119285, Y => HIEFFPLA_NET_0_119834);
    
    HIEFFPLA_INST_0_48005 : MX2
      port map(A => HIEFFPLA_NET_0_118399, B => 
        HIEFFPLA_NET_0_118395, S => \BIT_OS_SEL_3[0]\, Y => 
        \U_ELK15_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[2]\);
    
    \U_ELK16_CH/U_SLAVE_1ELK/Q[2]\ : DFN1C0
      port map(D => \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/Q[2]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/Q[3]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[3]_net_1\, CLK => 
        CCC_160M_FXD, CLR => P_MASTER_POR_B_c_34, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/Q[3]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/PHASE_ADJ[4]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[4]_net_1\, CLK
         => CLK_40M_GL, CLR => P_MASTER_POR_B_c, Q => 
        \U_MASTER_DES/PHASE_ADJ_160_L[4]\);
    
    \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[6]\ : DFN1C0
      port map(D => \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\);
    
    HIEFFPLA_INST_0_39353 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_1[7]\, B => 
        HIEFFPLA_NET_0_119516, S => HIEFFPLA_NET_0_119243, Y => 
        HIEFFPLA_NET_0_120000);
    
    \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[11]\ : DFN1C0
      port map(D => 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[11]_net_1\);
    
    HIEFFPLA_INST_0_62986 : MX2
      port map(A => HIEFFPLA_NET_0_115885, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[9]\, S => 
        HIEFFPLA_NET_0_117073, Y => HIEFFPLA_NET_0_115921);
    
    HIEFFPLA_INST_0_47590 : MX2
      port map(A => 
        \U_ELK14_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]_net_1\, B => 
        \U_ELK14_CH/ELK_TX_DAT[4]\, S => 
        \U_ELK14_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118470);
    
    HIEFFPLA_INST_0_50597 : MX2
      port map(A => 
        \U_ELK7_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]_net_1\, B => 
        \U_ELK7_CH/ELK_TX_DAT[5]\, S => 
        \U_ELK7_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_117926);
    
    HIEFFPLA_INST_0_45559 : AO1A
      port map(A => HIEFFPLA_NET_0_119475, B => 
        \U50_PATTERNS/ELINKS_STOP_ADDR[7]\, C => 
        HIEFFPLA_NET_0_118805, Y => HIEFFPLA_NET_0_118890);
    
    HIEFFPLA_INST_0_58282 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_13[1]\, B => 
        HIEFFPLA_NET_0_116537, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_0[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116541);
    
    \U_ELK3_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]\ : DFN1C0
      port map(D => \U_ELK3_CH/U_SLAVE_1ELK/Q[12]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]_net_1\);
    
    \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[4]\ : DFN1C0
      port map(D => \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\);
    
    \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[2]\ : DFN1C0
      port map(D => 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[2]_net_1\);
    
    HIEFFPLA_INST_0_42634 : AOI1C
      port map(A => HIEFFPLA_NET_0_119408, B => 
        HIEFFPLA_NET_0_119553, C => 
        \U50_PATTERNS/REG_STATE_0[4]_net_1\, Y => 
        HIEFFPLA_NET_0_119495);
    
    \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[3]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[1]_net_1\, CLK => 
        CCC_160M_ADJ, CLR => P_MASTER_POR_B_c_34_0, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[3]_net_1\);
    
    \DEV_RST_B_pad/U0/U1\ : IOIN_IB
      port map(YIN => \DEV_RST_B_pad/U0/NET1\, Y => DEV_RST_B_c);
    
    HIEFFPLA_INST_0_45292 : AO1A
      port map(A => HIEFFPLA_NET_0_118828, B => 
        \U50_PATTERNS/SM_BANK_SEL[4]\, C => HIEFFPLA_NET_0_118820, 
        Y => HIEFFPLA_NET_0_118949);
    
    HIEFFPLA_INST_0_111900 : AO1A
      port map(A => \U50_PATTERNS/RD_USB_ADBUS[6]\, B => 
        HIEFFPLA_NET_0_119557, C => \U50_PATTERNS/USB_RXF_B\, Y
         => HIEFFPLA_NET_0_115824);
    
    \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[5]\ : DFN1C0
      port map(D => \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\);
    
    AFLSDF_INV_10 : INV
      port map(A => P_USB_MASTER_EN_c_22_0, Y => \AFLSDF_INV_10\);
    
    HIEFFPLA_INST_0_59730 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_30[0]\, B => 
        HIEFFPLA_NET_0_116350, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_1[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116356);
    
    HIEFFPLA_INST_0_53763 : AO1E
      port map(A => HIEFFPLA_NET_0_116678, B => 
        HIEFFPLA_NET_0_116593, C => HIEFFPLA_NET_0_117328, Y => 
        HIEFFPLA_NET_0_117357);
    
    HIEFFPLA_INST_0_43018 : AO1D
      port map(A => HIEFFPLA_NET_0_119380, B => 
        HIEFFPLA_NET_0_119432, C => HIEFFPLA_NET_0_119375, Y => 
        HIEFFPLA_NET_0_119401);
    
    \U_EXEC_MASTER/USB_MASTER_EN/CNT_EN_60M1S\ : DFN1C0
      port map(D => 
        \U_EXEC_MASTER/USB_MASTER_EN/CNT_EN_60M0S_net_1\, CLK => 
        CLK60MHZ, CLR => P_MASTER_POR_B_c_23, Q => 
        \U_EXEC_MASTER/USB_MASTER_EN/CNT_EN_60M1S_net_1\);
    
    HIEFFPLA_INST_0_57419 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_4[8]\, B => 
        HIEFFPLA_NET_0_116663, S => HIEFFPLA_NET_0_117122, Y => 
        HIEFFPLA_NET_0_116688);
    
    HIEFFPLA_INST_0_44352 : MX2
      port map(A => \TFC_STOP_ADDR[1]\, B => 
        \U50_PATTERNS/U4B_REGCROSS/SAMP_TWO[1]_net_1\, S => 
        HIEFFPLA_NET_0_119135, Y => HIEFFPLA_NET_0_119132);
    
    HIEFFPLA_INST_0_47174 : MX2
      port map(A => \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\, 
        B => \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\, S => 
        \BIT_OS_SEL_4[2]\, Y => HIEFFPLA_NET_0_118539);
    
    HIEFFPLA_INST_0_45162 : NAND3C
      port map(A => HIEFFPLA_NET_0_118880, B => 
        HIEFFPLA_NET_0_118732, C => HIEFFPLA_NET_0_118803, Y => 
        HIEFFPLA_NET_0_118975);
    
    HIEFFPLA_INST_0_38063 : NAND2A
      port map(A => \U200B_ELINKS/RX_SER_WORD_2DEL[0]_net_1\, B
         => \U200B_ELINKS/RX_SER_WORD_2DEL[1]_net_1\, Y => 
        HIEFFPLA_NET_0_120162);
    
    \U50_PATTERNS/U4D_REGCROSS/SAMP_ONE[5]\ : DFN1C0
      port map(D => \U50_PATTERNS/ELINKS_STOP_ADDR[5]\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_25, Q => 
        \U50_PATTERNS/U4D_REGCROSS/SAMP_ONE[5]_net_1\);
    
    HIEFFPLA_INST_0_55468 : MX2
      port map(A => HIEFFPLA_NET_0_116110, B => 
        HIEFFPLA_NET_0_116014, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[3]\, Y => 
        HIEFFPLA_NET_0_117033);
    
    HIEFFPLA_INST_0_48116 : AND2
      port map(A => CLK_40M_GL, B => 
        \U_ELK16_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0_net_1\, Y => 
        HIEFFPLA_NET_0_118374);
    
    HIEFFPLA_INST_0_41953 : AND3C
      port map(A => HIEFFPLA_NET_0_119265, B => 
        HIEFFPLA_NET_0_119261, C => 
        \U50_PATTERNS/SM_BANK_SEL[17]\, Y => 
        HIEFFPLA_NET_0_119648);
    
    \U_ELK17_CH/U_ELK1_CMD_TX/SER_OUT_FI\ : DFN1C0
      port map(D => 
        \U_ELK17_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_0, Q => 
        \U_ELK17_CH/U_ELK1_CMD_TX/SER_OUT_FI_net_1\);
    
    HIEFFPLA_INST_0_44240 : MX2
      port map(A => \TFC_STRT_ADDR[0]\, B => 
        \U50_PATTERNS/U4A_REGCROSS/SAMP_TWO[0]_net_1\, S => 
        HIEFFPLA_NET_0_119156, Y => HIEFFPLA_NET_0_119154);
    
    \U_ELK5_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]\ : DFN1C0
      port map(D => \U_ELK5_CH/U_SLAVE_1ELK/Q[4]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]_net_1\);
    
    \U200A_TFC/GP_PG_SM[5]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120316, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_28, Q => 
        \U200A_TFC/GP_PG_SM[5]_net_1\);
    
    HIEFFPLA_INST_0_58009 : XA1C
      port map(A => HIEFFPLA_NET_0_116590, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_7[5]\, C => 
        HIEFFPLA_NET_0_117179, Y => HIEFFPLA_NET_0_116579);
    
    HIEFFPLA_INST_0_55082 : NAND3C
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[8]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[0]_net_1\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[5]_net_1\, Y => 
        HIEFFPLA_NET_0_117125);
    
    HIEFFPLA_INST_0_37850 : AO1E
      port map(A => \OP_MODE_c[6]\, B => HIEFFPLA_NET_0_120190, C
         => \U200B_ELINKS/GP_PG_SM[2]_net_1\, Y => 
        HIEFFPLA_NET_0_120191);
    
    HIEFFPLA_INST_0_61166 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_1[0]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_2[0]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_1[0]\, Y => 
        HIEFFPLA_NET_0_116165);
    
    HIEFFPLA_INST_0_42698 : AND3C
      port map(A => HIEFFPLA_NET_0_119510, B => 
        HIEFFPLA_NET_0_119410, C => HIEFFPLA_NET_0_119459, Y => 
        HIEFFPLA_NET_0_119480);
    
    \U_ELK13_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]\ : DFN1C0
      port map(D => \U_ELK13_CH/U_SLAVE_1ELK/Q[13]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]_net_1\);
    
    \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[8]\ : DFN1C0
      port map(D => \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\);
    
    HIEFFPLA_INST_0_38458 : MX2
      port map(A => \U50_PATTERNS/ELINKS_STRT_ADDR_T[3]\, B => 
        \U50_PATTERNS/RD_USB_ADBUS[3]\, S => 
        HIEFFPLA_NET_0_119493, Y => HIEFFPLA_NET_0_120100);
    
    \U_ELK2_CH/U_SLAVE_1ELK/RECD_SER_WORD[6]\ : DFN1C0
      port map(D => \U_ELK2_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[6]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_2[6]\);
    
    HIEFFPLA_INST_0_46871 : AND2
      port map(A => CLK_40M_GL, B => 
        \U_ELK11_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0_net_1\, Y => 
        HIEFFPLA_NET_0_118599);
    
    \U_ELK15_CH/U_SLAVE_1ELK/Q[7]\ : DFN1C0
      port map(D => \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/Q[7]_net_1\);
    
    HIEFFPLA_INST_0_46511 : AND3B
      port map(A => \U50_PATTERNS/RD_USB_ADBUS[5]\, B => 
        \U50_PATTERNS/WR_XFER_TYPE[0]_net_1\, C => 
        \U50_PATTERNS/RD_USB_ADBUS[1]\, Y => 
        HIEFFPLA_NET_0_118676);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_2[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116032, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_10, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_2[3]\);
    
    \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[14]\ : DFN1C0
      port map(D => \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[14]_net_1\);
    
    HIEFFPLA_INST_0_63150 : AND3
      port map(A => HIEFFPLA_NET_0_117125, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[0]_net_1\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[1]_net_1\, Y => 
        HIEFFPLA_NET_0_115876);
    
    HIEFFPLA_INST_0_55406 : AO1
      port map(A => HIEFFPLA_NET_0_117087, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[3]\, C => 
        HIEFFPLA_NET_0_117008, Y => HIEFFPLA_NET_0_117042);
    
    HIEFFPLA_INST_0_53126 : MX2
      port map(A => HIEFFPLA_NET_0_117546, B => 
        HIEFFPLA_NET_0_117542, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[3]\, Y => 
        HIEFFPLA_NET_0_117462);
    
    HIEFFPLA_INST_0_111664 : MX2
      port map(A => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[7]_net_1\, B => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[71]_net_1\, S => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[6]\, Y => 
        HIEFFPLA_NET_0_115834);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_31[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116343, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_20, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_31[0]\);
    
    HIEFFPLA_INST_0_50674 : MX2
      port map(A => \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\, B
         => \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\, S => 
        \BIT_OS_SEL_4[2]\, Y => HIEFFPLA_NET_0_117907);
    
    \U_ELK10_CH/U_ELK1_SERDAT_SOURCE/SERDAT[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118641, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_17, Q => 
        \U_ELK10_CH/ELK_TX_DAT[2]\);
    
    \U50_PATTERNS/WR_XFER_TYPE[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118687, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c, Q => 
        \U50_PATTERNS/WR_XFER_TYPE[2]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_23[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116441, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_17_0, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_23[1]\);
    
    HIEFFPLA_INST_0_43191 : NAND3C
      port map(A => HIEFFPLA_NET_0_119340, B => 
        HIEFFPLA_NET_0_119342, C => HIEFFPLA_NET_0_119344, Y => 
        HIEFFPLA_NET_0_119350);
    
    \U50_PATTERNS/ELINK_RWA[19]/U1\ : DFN1P0
      port map(D => HIEFFPLA_NET_0_119701, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_12, Q => 
        \U50_PATTERNS/ELINK_RWA[19]\);
    
    HIEFFPLA_INST_0_43130 : NAND3C
      port map(A => HIEFFPLA_NET_0_119350, B => 
        HIEFFPLA_NET_0_119420, C => HIEFFPLA_NET_0_119361, Y => 
        HIEFFPLA_NET_0_119364);
    
    \U_ELK1_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]\ : DFN1C0
      port map(D => \U_ELK1_CH/U_SLAVE_1ELK/Q[5]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]_net_1\);
    
    HIEFFPLA_INST_0_60330 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_9[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_25[1]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[4]_net_1\, Y
         => HIEFFPLA_NET_0_116280);
    
    \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[3]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_WRD_40M_FIXED[3]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_27, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[3]_net_1\);
    
    HIEFFPLA_INST_0_61613 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_24[3]\, B => 
        HIEFFPLA_NET_0_117186, S => HIEFFPLA_NET_0_117074, Y => 
        HIEFFPLA_NET_0_116102);
    
    HIEFFPLA_INST_0_54277 : MX2
      port map(A => HIEFFPLA_NET_0_116443, B => 
        HIEFFPLA_NET_0_116524, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_2[3]_net_1\, Y
         => HIEFFPLA_NET_0_117286);
    
    \U_ELK0_CMD_TX/SER_CMD_WORD_R[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118665, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_14, Q => 
        \U_ELK0_CMD_TX/SER_CMD_WORD_R[0]_net_1\);
    
    HIEFFPLA_INST_0_57528 : AND3
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_4[6]\, B => 
        HIEFFPLA_NET_0_116672, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_4[7]\, Y => 
        HIEFFPLA_NET_0_116662);
    
    HIEFFPLA_INST_0_47871 : NAND2B
      port map(A => \OP_MODE_c_6[1]\, B => \PATT_ELK_DAT_15[3]\, 
        Y => HIEFFPLA_NET_0_118415);
    
    HIEFFPLA_INST_0_42264 : AND2B
      port map(A => \U50_PATTERNS/USB_RXF_B\, B => 
        \U50_PATTERNS/RD_USB_ADBUS[6]\, Y => 
        HIEFFPLA_NET_0_119586);
    
    \U50_PATTERNS/TFC_STOP_ADDR[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119183, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_8, Q => 
        \U50_PATTERNS/TFC_STOP_ADDR[5]\);
    
    HIEFFPLA_INST_0_49368 : AND2A
      port map(A => \OP_MODE_c_1[1]\, B => \PATT_ELK_DAT_2[6]\, Y
         => HIEFFPLA_NET_0_118142);
    
    HIEFFPLA_INST_0_53182 : MX2
      port map(A => HIEFFPLA_NET_0_117531, B => 
        HIEFFPLA_NET_0_117523, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_2[3]\, Y => 
        HIEFFPLA_NET_0_117455);
    
    HIEFFPLA_INST_0_41883 : AOI1B
      port map(A => HIEFFPLA_NET_0_119389, B => 
        \U50_PATTERNS/SM_BANK_SEL[15]\, C => 
        HIEFFPLA_NET_0_119644, Y => HIEFFPLA_NET_0_119675);
    
    \U_MASTER_DES/U13C_MASTER_DESER/ARB_WRD_40M_FIXED[8]\ : 
        DFN1C0
      port map(D => \U_MASTER_DES/U13C_MASTER_DESER/Q[8]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_26, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_WRD_40M_FIXED[8]_net_1\);
    
    HIEFFPLA_INST_0_48620 : AND2A
      port map(A => \OP_MODE_c_2[1]\, B => \PATT_ELK_DAT_18[5]\, 
        Y => HIEFFPLA_NET_0_118278);
    
    \U50_PATTERNS/ELINK_ADDRA_4[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119980, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_2_0, Q => 
        \U50_PATTERNS/ELINK_ADDRA_4[3]\);
    
    HIEFFPLA_INST_0_55882 : MX2
      port map(A => HIEFFPLA_NET_0_116967, B => 
        HIEFFPLA_NET_0_116993, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[1]\, Y => 
        HIEFFPLA_NET_0_116978);
    
    HIEFFPLA_INST_0_47463 : MX2
      port map(A => \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\, 
        B => \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[13]_net_1\, S => 
        \BIT_OS_SEL_3[2]\, Y => HIEFFPLA_NET_0_118488);
    
    HIEFFPLA_INST_0_52224 : AND3B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[7]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[0]_net_1\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[7]_net_1\, Y => 
        HIEFFPLA_NET_0_117607);
    
    HIEFFPLA_INST_0_56246 : AND2
      port map(A => DCB_SALT_SEL_c, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/RECD_SER_WORD[6]_net_1\, 
        Y => \ELK_RX_SER_WORD_0[6]\);
    
    HIEFFPLA_INST_0_47128 : NAND2B
      port map(A => \OP_MODE_c_3[1]\, B => \PATT_ELK_DAT_12[7]\, 
        Y => HIEFFPLA_NET_0_118546);
    
    HIEFFPLA_INST_0_41557 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_8[3]\, B => 
        HIEFFPLA_NET_0_119574, S => HIEFFPLA_NET_0_119291, Y => 
        HIEFFPLA_NET_0_119724);
    
    \U50_PATTERNS/ELINK_DINA_18[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119797, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_21, Q => 
        \U50_PATTERNS/ELINK_DINA_18[2]\);
    
    HIEFFPLA_INST_0_50612 : AND2A
      port map(A => \OP_MODE_c_4[1]\, B => \PATT_ELK_DAT_7[5]\, Y
         => HIEFFPLA_NET_0_117918);
    
    HIEFFPLA_INST_0_45259 : AO1
      port map(A => HIEFFPLA_NET_0_119241, B => 
        \U50_PATTERNS/ELINK_DOUTA_1[2]\, C => 
        HIEFFPLA_NET_0_118835, Y => HIEFFPLA_NET_0_118956);
    
    \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[9]\ : DFN1C0
      port map(D => \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\);
    
    \U_ELK6_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL\ : DFN1C0
      port map(D => \U_ELK6_CH/ELK_IN_F_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL_net_1\);
    
    \U_ELK3_CH/U_SLAVE_1ELK/Q[14]\ : DFN1C0
      port map(D => \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[14]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/Q[14]_net_1\);
    
    HIEFFPLA_INST_0_40549 : MX2
      port map(A => HIEFFPLA_NET_0_119574, B => 
        \U50_PATTERNS/ELINK_DINA_13[3]\, S => 
        HIEFFPLA_NET_0_119285, Y => HIEFFPLA_NET_0_119836);
    
    HIEFFPLA_INST_0_50808 : MX2
      port map(A => \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[0]_net_1\, B
         => \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\, S => 
        \BIT_OS_SEL_4[2]\, Y => HIEFFPLA_NET_0_117889);
    
    HIEFFPLA_INST_0_47531 : MX2
      port map(A => HIEFFPLA_NET_0_118495, B => 
        HIEFFPLA_NET_0_118492, S => \BIT_OS_SEL_4[0]\, Y => 
        \U_ELK13_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[5]\);
    
    HIEFFPLA_INST_0_42356 : NOR3A
      port map(A => HIEFFPLA_NET_0_119565, B => 
        HIEFFPLA_NET_0_119582, C => HIEFFPLA_NET_0_119581, Y => 
        HIEFFPLA_NET_0_119558);
    
    \U50_PATTERNS/TFC_STRT_ADDR_T[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119164, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_4, Q => 
        \U50_PATTERNS/TFC_STRT_ADDR_T[0]\);
    
    \U_ELK14_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL\ : DFN1C0
      port map(D => \U_ELK14_CH/ELK_IN_F_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL_net_1\);
    
    \U50_PATTERNS/ELINK_DINA_18[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119799, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_20, Q => 
        \U50_PATTERNS/ELINK_DINA_18[0]\);
    
    \U_ELK12_CH/U_SLAVE_1ELK/Q[3]\ : DFN1C0
      port map(D => \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/Q[3]_net_1\);
    
    HIEFFPLA_INST_0_54253 : MX2
      port map(A => HIEFFPLA_NET_0_116568, B => 
        HIEFFPLA_NET_0_116286, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_1[3]_net_1\, Y
         => HIEFFPLA_NET_0_117289);
    
    \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[3]\ : DFN1C0
      port map(D => 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[3]_net_1\);
    
    HIEFFPLA_INST_0_45606 : NAND3C
      port map(A => HIEFFPLA_NET_0_118716, B => 
        HIEFFPLA_NET_0_118725, C => HIEFFPLA_NET_0_118733, Y => 
        HIEFFPLA_NET_0_118881);
    
    HIEFFPLA_INST_0_45390 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_19[0]\, C => 
        \U50_PATTERNS/SM_BANK_SEL[0]\, Y => HIEFFPLA_NET_0_118922);
    
    HIEFFPLA_INST_0_47829 : AND2
      port map(A => \U_ELK15_CH/ELK_TX_DAT[0]\, B => 
        \U_ELK15_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118427);
    
    HIEFFPLA_INST_0_45300 : NAND3C
      port map(A => HIEFFPLA_NET_0_118818, B => 
        HIEFFPLA_NET_0_118826, C => HIEFFPLA_NET_0_118829, Y => 
        HIEFFPLA_NET_0_118947);
    
    \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[1]\ : DFN1C0
      port map(D => 
        \U_ELK9_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\);
    
    \U_ELK7_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]\ : DFN1C0
      port map(D => \U_ELK7_CH/U_SLAVE_1ELK/Q[0]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]_net_1\);
    
    \U_ELK19_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]\ : DFN1C0
      port map(D => \U_ELK19_CH/U_SLAVE_1ELK/Q[11]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]_net_1\);
    
    HIEFFPLA_INST_0_52273 : NAND3B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[7]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[5]_net_1\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[0]_net_1\, Y => 
        HIEFFPLA_NET_0_117595);
    
    \U_ELK2_CH/U_ELK1_SERDAT_SOURCE/SERDAT[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118146, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_13, Q => 
        \U_ELK2_CH/ELK_TX_DAT[2]\);
    
    HIEFFPLA_INST_0_43660 : NAND2B
      port map(A => \U50_PATTERNS/SM_BANK_SEL_0[21]\, B => 
        \U50_PATTERNS/SM_BANK_SEL[14]\, Y => 
        HIEFFPLA_NET_0_119251);
    
    \U_ELK11_CH/U_ELK1_CMD_TX/SER_OUT_FI\ : DFN1C0
      port map(D => 
        \U_ELK11_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_2, Q => 
        \U_ELK11_CH/U_ELK1_CMD_TX/SER_OUT_FI_net_1\);
    
    \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[5]\ : DFN1C0
      port map(D => \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\);
    
    \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[1]\ : DFN1C0
      port map(D => 
        \U_ELK10_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\);
    
    HIEFFPLA_INST_0_62334 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_3[2]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_4[2]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_4[0]\, Y => 
        HIEFFPLA_NET_0_116002);
    
    HIEFFPLA_INST_0_58975 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_5[2]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_21[2]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_5[4]_net_1\, Y
         => HIEFFPLA_NET_0_116452);
    
    HIEFFPLA_INST_0_49033 : MX2
      port map(A => HIEFFPLA_NET_0_118224, B => 
        HIEFFPLA_NET_0_118222, S => \BIT_OS_SEL_2[0]\, Y => 
        \U_ELK19_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[6]\);
    
    \U50_PATTERNS/ELINK_DINA_13[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119839, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_14, Q => 
        \U50_PATTERNS/ELINK_DINA_13[0]\);
    
    HIEFFPLA_INST_0_48397 : MX2
      port map(A => \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[3]_net_1\, 
        B => \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\, S => 
        \BIT_OS_SEL_0[2]\, Y => HIEFFPLA_NET_0_118317);
    
    \U_EXEC_MASTER/MPOR_B_13\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117787, CLK => CLK_40M_GL, CLR
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_1\, Q => 
        P_MASTER_POR_B_c_13);
    
    \U_ELK16_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2\ : IOPADN_BI
      port map(DB => \U_ELK16_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, 
        E => \U_ELK16_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET3\, PAD
         => ELK16_DAT_N, N2POUT => 
        \U_ELK16_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2_N2P\);
    
    HIEFFPLA_INST_0_56064 : AXOI4
      port map(A => HIEFFPLA_NET_0_117112, B => 
        HIEFFPLA_NET_0_117084, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/MAX_CNT[0]\, Y => 
        HIEFFPLA_NET_0_116954);
    
    \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[11]\ : DFN1C0
      port map(D => \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\);
    
    \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[7]\ : DFN1C0
      port map(D => 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\);
    
    HIEFFPLA_INST_0_56239 : AND2A
      port map(A => DCB_SALT_SEL_c, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/RECD_SER_WORD[2]_net_1\, 
        Y => \TFC_RX_SER_WORD[2]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_16[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116214, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_5, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_16[1]\);
    
    HIEFFPLA_INST_0_57655 : AOI1A
      port map(A => HIEFFPLA_NET_0_116648, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_5[0]\, C => 
        HIEFFPLA_NET_0_116641, Y => HIEFFPLA_NET_0_116642);
    
    \U50_PATTERNS/U4A_REGCROSS/SAMP_ONE[2]\ : DFN1C0
      port map(D => \U50_PATTERNS/TFC_STRT_ADDR[2]\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_32, Q => 
        \U50_PATTERNS/U4A_REGCROSS/SAMP_ONE[2]_net_1\);
    
    \U_ELK12_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]\ : DFN1C0
      port map(D => \U_ELK12_CH/U_SLAVE_1ELK/Q[13]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]_net_1\);
    
    HIEFFPLA_INST_0_52824 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_7[3]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_8[3]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_2[0]\, Y => 
        HIEFFPLA_NET_0_117505);
    
    \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[3]\ : DFN1C0
      port map(D => \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\);
    
    \U50_PATTERNS/U4A_REGCROSS/SAMP_ONE[7]\ : DFN1C0
      port map(D => \U50_PATTERNS/TFC_STRT_ADDR[7]\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_32_0, Q => 
        \U50_PATTERNS/U4A_REGCROSS/SAMP_ONE[7]_net_1\);
    
    \U50_PATTERNS/ELINK_ADDRA_3[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119989, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_1, Q => 
        \U50_PATTERNS/ELINK_ADDRA_3[2]\);
    
    \U50_PATTERNS/ELINK_ADDRA_18[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120020, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_12, Q => 
        \U50_PATTERNS/ELINK_ADDRA_18[3]\);
    
    HIEFFPLA_INST_0_38606 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_10[4]\, B => 
        HIEFFPLA_NET_0_119519, S => HIEFFPLA_NET_0_119239, Y => 
        HIEFFPLA_NET_0_120083);
    
    \U50_PATTERNS/TFC_STRT_ADDR_T[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119163, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_4, Q => 
        \U50_PATTERNS/TFC_STRT_ADDR_T[1]\);
    
    HIEFFPLA_INST_0_38229 : AND2A
      port map(A => HIEFFPLA_NET_0_119452, B => 
        \U50_PATTERNS/RD_USB_ADBUS[3]\, Y => 
        HIEFFPLA_NET_0_120132);
    
    HIEFFPLA_INST_0_37673 : NAND2B
      port map(A => \U200B_ELINKS/GP_PG_SM[2]_net_1\, B => 
        \U200B_ELINKS/GP_PG_SM[3]_net_1\, Y => 
        HIEFFPLA_NET_0_120234);
    
    HIEFFPLA_INST_0_44504 : MX2
      port map(A => \ELKS_STRT_ADDR[7]\, B => 
        \U50_PATTERNS/U4C_REGCROSS/SAMP_TWO[7]_net_1\, S => 
        HIEFFPLA_NET_0_119114, Y => HIEFFPLA_NET_0_119105);
    
    HIEFFPLA_INST_0_40945 : MX2
      port map(A => HIEFFPLA_NET_0_119560, B => 
        \U50_PATTERNS/ELINK_DINA_18[7]\, S => 
        HIEFFPLA_NET_0_119264, Y => HIEFFPLA_NET_0_119792);
    
    \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[12]\ : DFN1C0
      port map(D => 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[12]_net_1\);
    
    \U50_PATTERNS/SI_CNT[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119332, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_5, Q => \U50_PATTERNS/SI_CNT[2]\);
    
    HIEFFPLA_INST_0_45887 : AO1
      port map(A => HIEFFPLA_NET_0_119288, B => 
        \U50_PATTERNS/ELINK_DOUTA_16[0]\, C => 
        HIEFFPLA_NET_0_118765, Y => HIEFFPLA_NET_0_118820);
    
    HIEFFPLA_INST_0_42983 : NAND3C
      port map(A => HIEFFPLA_NET_0_119631, B => 
        HIEFFPLA_NET_0_119374, C => HIEFFPLA_NET_0_119409, Y => 
        HIEFFPLA_NET_0_119410);
    
    \U_ELK16_CH/U_ELK1_CMD_TX/SER_OUT_FDEL\ : DFN1C0
      port map(D => \U_ELK16_CH/U_ELK1_CMD_TX/SER_OUT_FI_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_1, Q
         => \U_ELK16_CH/ELK_OUT_F\);
    
    HIEFFPLA_INST_0_54951 : AND3A
      port map(A => HIEFFPLA_NET_0_117245, B => 
        HIEFFPLA_NET_0_117242, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_3[6]_net_1\, Y => 
        HIEFFPLA_NET_0_117160);
    
    HIEFFPLA_INST_0_41467 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_7[1]\, B => 
        HIEFFPLA_NET_0_119576, S => HIEFFPLA_NET_0_119289, Y => 
        HIEFFPLA_NET_0_119734);
    
    \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[13]\ : DFN1C0
      port map(D => 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[13]_net_1\);
    
    HIEFFPLA_INST_0_54884 : AO1B
      port map(A => HIEFFPLA_NET_0_117365, B => 
        HIEFFPLA_NET_0_117106, C => HIEFFPLA_NET_0_117179, Y => 
        HIEFFPLA_NET_0_117182);
    
    HIEFFPLA_INST_0_39416 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_2[6]\, B => 
        HIEFFPLA_NET_0_119517, S => HIEFFPLA_NET_0_119278, Y => 
        HIEFFPLA_NET_0_119993);
    
    HIEFFPLA_INST_0_57140 : XA1B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_2[3]\, B => 
        HIEFFPLA_NET_0_116746, C => HIEFFPLA_NET_0_117179, Y => 
        HIEFFPLA_NET_0_116732);
    
    \U_ELK15_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]\ : DFN1C0
      port map(D => \U_ELK15_CH/U_SLAVE_1ELK/Q[13]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]_net_1\);
    
    \U_ELK19_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL\ : DFN1C0
      port map(D => \U_ELK19_CH/ELK_IN_F_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL_net_1\);
    
    \U_ELK11_CH/U_SLAVE_1ELK/RECD_SER_WORD[3]\ : DFN1C0
      port map(D => \U_ELK11_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[3]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_11[3]\);
    
    \U50_PATTERNS/ELINK_ADDRA_2[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119993, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_21, Q => 
        \U50_PATTERNS/ELINK_ADDRA_2[6]\);
    
    \U_ELK11_CH/U_SLAVE_1ELK/RECD_SER_WORD[6]\ : DFN1C0
      port map(D => \U_ELK11_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[6]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_11[6]\);
    
    HIEFFPLA_INST_0_56146 : NAND2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/MAX_CNT[0]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/MAX_CNT[1]\, Y => 
        HIEFFPLA_NET_0_116944);
    
    HIEFFPLA_INST_0_50626 : MX2
      port map(A => HIEFFPLA_NET_0_117910, B => 
        HIEFFPLA_NET_0_117908, S => \BIT_OS_SEL_4[1]\, Y => 
        HIEFFPLA_NET_0_117914);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_15[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116228, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_4, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_15[2]\);
    
    HIEFFPLA_INST_0_63036 : NAND3A
      port map(A => HIEFFPLA_NET_0_115920, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[6]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[5]\, Y => 
        HIEFFPLA_NET_0_115907);
    
    \U_ELK16_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL\ : DFN1C0
      port map(D => \U_ELK16_CH/ELK_IN_R_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL_net_1\);
    
    \U50_PATTERNS/ELINKS_STRT_ADDR[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120106, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_17, Q => 
        \U50_PATTERNS/ELINKS_STRT_ADDR[5]\);
    
    HIEFFPLA_INST_0_56241 : AND2A
      port map(A => DCB_SALT_SEL_c, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/RECD_SER_WORD[3]_net_1\, 
        Y => \TFC_RX_SER_WORD[3]\);
    
    \U_ELK15_CH/U_SLAVE_1ELK/Q[11]\ : DFN1C0
      port map(D => \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/Q[11]_net_1\);
    
    \U50_PATTERNS/ELINK_DINA_5[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119750, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_14, Q => 
        \U50_PATTERNS/ELINK_DINA_5[1]\);
    
    HIEFFPLA_INST_0_42816 : OA1A
      port map(A => \U50_PATTERNS/REG_STATE_0[2]_net_1\, B => 
        \U50_PATTERNS/REG_STATE_0[1]_net_1\, C => 
        \U50_PATTERNS/REG_STATE[3]_net_1\, Y => 
        HIEFFPLA_NET_0_119457);
    
    \U_ELK17_CH/U_SLAVE_1ELK/RECD_SER_WORD[6]\ : DFN1C0
      port map(D => \U_ELK17_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[6]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_17[6]\);
    
    HIEFFPLA_INST_0_50863 : NAND2B
      port map(A => \OP_MODE_c_0[1]\, B => \PATT_ELK_DAT_8[7]\, Y
         => HIEFFPLA_NET_0_117871);
    
    \U_ELK14_CH/U_SLAVE_1ELK/Q[1]\ : DFN1C0
      port map(D => \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/Q[1]_net_1\);
    
    \U50_PATTERNS/ELINK_ADDRA_1[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120005, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_20, Q => 
        \U50_PATTERNS/ELINK_ADDRA_1[2]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_SEL_5[1]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_BIT_OS_VAL[1]\, CLK
         => CLK_40M_GL, CLR => P_MASTER_POR_B_c_27_0, Q => 
        \BIT_OS_SEL_5[1]\);
    
    \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[2]\ : DFN1C0
      port map(D => 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[2]_net_1\);
    
    \U_ELK5_CH/U_SLAVE_1ELK/Q[11]\ : DFN1C0
      port map(D => \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/Q[11]_net_1\);
    
    HIEFFPLA_INST_0_47041 : MX2
      port map(A => HIEFFPLA_NET_0_118583, B => 
        HIEFFPLA_NET_0_118580, S => \BIT_OS_SEL[0]\, Y => 
        \U_ELK11_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[6]\);
    
    HIEFFPLA_INST_0_61139 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_1[2]\, 
        B => HIEFFPLA_NET_0_117181, S => HIEFFPLA_NET_0_117149, Y
         => HIEFFPLA_NET_0_116168);
    
    HIEFFPLA_INST_0_41941 : AND3C
      port map(A => HIEFFPLA_NET_0_119245, B => 
        HIEFFPLA_NET_0_119262, C => \U50_PATTERNS/SM_BANK_SEL[7]\, 
        Y => HIEFFPLA_NET_0_119653);
    
    \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117621, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_22, Q => 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM[0]_net_1\);
    
    \U50_PATTERNS/U4A_REGCROSS/SAMP_ONE[1]\ : DFN1C0
      port map(D => \U50_PATTERNS/TFC_STRT_ADDR[1]\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_32, Q => 
        \U50_PATTERNS/U4A_REGCROSS/SAMP_ONE[1]_net_1\);
    
    HIEFFPLA_INST_0_57107 : NAND3C
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_2[6]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_2[8]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_2[7]\, Y => 
        HIEFFPLA_NET_0_116741);
    
    HIEFFPLA_INST_0_56772 : NAND2A
      port map(A => HIEFFPLA_NET_0_116805, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_0[5]\, Y => 
        HIEFFPLA_NET_0_116801);
    
    HIEFFPLA_INST_0_51347 : MX2
      port map(A => HIEFFPLA_NET_0_117776, B => 
        \U_EXEC_MASTER/DEL_CNT[2]\, S => HIEFFPLA_NET_0_117796, Y
         => HIEFFPLA_NET_0_117793);
    
    \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[7]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117055, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_27, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[7]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/BEST_SEQCNT[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117440, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_8, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_SEQCNT[2]\);
    
    \U_ELK19_CH/U_SLAVE_1ELK/Q[12]\ : DFN1C0
      port map(D => \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/Q[12]_net_1\);
    
    HIEFFPLA_INST_0_45534 : NOR2A
      port map(A => \U50_PATTERNS/ELINKS_STRT_ADDR[2]\, B => 
        HIEFFPLA_NET_0_119428, Y => HIEFFPLA_NET_0_118895);
    
    HIEFFPLA_INST_0_39164 : MX2
      port map(A => HIEFFPLA_NET_0_119522, B => 
        \U50_PATTERNS/ELINK_ADDRA_18[2]\, S => 
        HIEFFPLA_NET_0_119264, Y => HIEFFPLA_NET_0_120021);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_7[6]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116597, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_14, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_7[6]\);
    
    HIEFFPLA_INST_0_54964 : AO1C
      port map(A => HIEFFPLA_NET_0_117341, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_3[6]_net_1\, C => 
        HIEFFPLA_NET_0_117115, Y => HIEFFPLA_NET_0_117154);
    
    \U_ELK5_CH/U_SLAVE_1ELK/Q[1]\ : DFN1C0
      port map(D => \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/Q[1]_net_1\);
    
    HIEFFPLA_INST_0_42467 : MX2
      port map(A => \U50_PATTERNS/REG_ADDR[3]\, B => 
        HIEFFPLA_NET_0_119506, S => HIEFFPLA_NET_0_119007, Y => 
        HIEFFPLA_NET_0_119530);
    
    HIEFFPLA_INST_0_62678 : AO13
      port map(A => HIEFFPLA_NET_0_115960, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_CLKPHASE[1]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_SEQCNT[2]\, Y => 
        HIEFFPLA_NET_0_115958);
    
    \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[14]\ : DFN1C0
      port map(D => 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[14]_net_1\);
    
    \U_ELK14_CH/U_ELK1_SERDAT_SOURCE/SERDAT[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118460, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_6, Q => 
        \U_ELK14_CH/ELK_TX_DAT[3]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_29[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116377, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_4, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_29[1]\);
    
    \U50_PATTERNS/ELINK_ADDRA_15[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120046, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_6, Q => 
        \U50_PATTERNS/ELINK_ADDRA_15[1]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_18[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116188, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_8, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_18[2]\);
    
    \U_ELK1_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118195, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_4, Q => 
        \U_ELK1_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]_net_1\);
    
    HIEFFPLA_INST_0_42667 : NAND3C
      port map(A => HIEFFPLA_NET_0_119490, B => 
        HIEFFPLA_NET_0_119404, C => HIEFFPLA_NET_0_119487, Y => 
        HIEFFPLA_NET_0_119488);
    
    \U_ELK2_CH/U_SLAVE_1ELK/Q[0]\ : DFN1C0
      port map(D => \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/Q[0]_net_1\);
    
    \P_USB_MASTER_EN_pad/U0/U0\ : IOPAD_TRI_U
      port map(D => \P_USB_MASTER_EN_pad/U0/NET1\, E => 
        \P_USB_MASTER_EN_pad/U0/NET2\, PAD => P_USB_MASTER_EN);
    
    HIEFFPLA_INST_0_38386 : MX2
      port map(A => \U50_PATTERNS/ELINKS_STRT_ADDR[2]\, B => 
        \U50_PATTERNS/ELINKS_STRT_ADDR_T[2]\, S => 
        HIEFFPLA_NET_0_119472, Y => HIEFFPLA_NET_0_120109);
    
    HIEFFPLA_INST_0_37301 : AND3B
      port map(A => \U200A_TFC/GP_PG_SM[2]_net_1\, B => 
        HIEFFPLA_NET_0_120299, C => \U200A_TFC/GP_PG_SM[3]_net_1\, 
        Y => HIEFFPLA_NET_0_120300);
    
    HIEFFPLA_INST_0_47372 : NAND2B
      port map(A => \OP_MODE_c[1]\, B => \PATT_ELK_DAT_13[2]\, Y
         => HIEFFPLA_NET_0_118506);
    
    HIEFFPLA_INST_0_161273 : DFN1C0
      port map(D => \U_ELK15_CH/ELK_TX_DAT[4]\, CLK => 
        CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_9, Q => 
        HIEFFPLA_NET_0_161282);
    
    HIEFFPLA_INST_0_57703 : AXOI4
      port map(A => HIEFFPLA_NET_0_117085, B => 
        HIEFFPLA_NET_0_117599, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_6[0]\, Y => 
        HIEFFPLA_NET_0_116632);
    
    HIEFFPLA_INST_0_44110 : MX2
      port map(A => \U50_PATTERNS/TFC_STRT_ADDR[0]\, B => 
        \U50_PATTERNS/TFC_STRT_ADDR_T[0]\, S => 
        HIEFFPLA_NET_0_119472, Y => HIEFFPLA_NET_0_119172);
    
    \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117619, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_22, Q => 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM[2]_net_1\);
    
    HIEFFPLA_INST_0_47698 : MX2
      port map(A => \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\, 
        B => \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[11]_net_1\, S => 
        \BIT_OS_SEL_2[2]\, Y => HIEFFPLA_NET_0_118445);
    
    \U_ELK19_CH/U_ELK1_SERDAT_SOURCE/SERDAT[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118235, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_15, Q => 
        \U_ELK19_CH/ELK_TX_DAT[3]\);
    
    HIEFFPLA_INST_0_54026 : AND3A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[1]_net_1\, B
         => \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[0]_net_1\, 
        C => \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_2[3]_net_1\, 
        Y => HIEFFPLA_NET_0_117318);
    
    \U_MASTER_DES/U13C_MASTER_DESER/ARB_WRD_40M_FIXED[9]\ : 
        DFN1C0
      port map(D => \U_MASTER_DES/U13C_MASTER_DESER/Q[9]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_26, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_WRD_40M_FIXED[9]_net_1\);
    
    \U_ELK2_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]\ : DFN1C0
      port map(D => \U_ELK2_CH/U_SLAVE_1ELK/Q[4]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]_net_1\);
    
    \U_ELK19_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U1\ : IOBI_ID_OD_EB
      port map(DR => \U_ELK19_CH/ELK_OUT_R\, DF => 
        \U_ELK19_CH/ELK_OUT_F\, CLR => \GND\, E => 
        \AFLSDF_INV_32\, ICLK => CCC_160M_ADJ, OCLK => 
        CCC_160M_FXD, YIN => 
        \U_ELK19_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\, DOUT => 
        \U_ELK19_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, EOUT => 
        \U_ELK19_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET2\, YR => 
        \U_ELK19_CH/ELK_IN_DDR_R\, YF => 
        \U_ELK19_CH/ELK_IN_DDR_F\);
    
    HIEFFPLA_INST_0_42422 : AND2
      port map(A => HIEFFPLA_NET_0_119473, B => 
        \U50_PATTERNS/RD_XFER_TYPE[1]_net_1\, Y => 
        HIEFFPLA_NET_0_119540);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_20[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116158, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_2, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_20[2]\);
    
    HIEFFPLA_INST_0_49925 : MX2
      port map(A => HIEFFPLA_NET_0_118044, B => 
        HIEFFPLA_NET_0_118040, S => \BIT_OS_SEL_6[1]\, Y => 
        HIEFFPLA_NET_0_118042);
    
    HIEFFPLA_INST_0_59737 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_30[1]\, B => 
        HIEFFPLA_NET_0_116349, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_1[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116355);
    
    \U50_PATTERNS/ELINK_DINA_12[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119845, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_12, Q => 
        \U50_PATTERNS/ELINK_DINA_12[2]\);
    
    HIEFFPLA_INST_0_59056 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_23[1]\, B => 
        HIEFFPLA_NET_0_116437, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_1[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116441);
    
    HIEFFPLA_INST_0_48700 : MX2
      port map(A => HIEFFPLA_NET_0_118273, B => 
        HIEFFPLA_NET_0_118271, S => \BIT_OS_SEL_0[1]\, Y => 
        HIEFFPLA_NET_0_118264);
    
    \U50_PATTERNS/ELINK_DINA_12[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119844, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_12, Q => 
        \U50_PATTERNS/ELINK_DINA_12[3]\);
    
    \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[9]\ : DFN1C0
      port map(D => \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\);
    
    HIEFFPLA_INST_0_57037 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_2[3]\, B => 
        HIEFFPLA_NET_0_116732, S => HIEFFPLA_NET_0_117601, Y => 
        HIEFFPLA_NET_0_116752);
    
    HIEFFPLA_INST_0_161274 : DFN1C0
      port map(D => \U_ELK15_CH/U_ELK1_CMD_TX/START_RISE_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_9, Q
         => HIEFFPLA_NET_0_161281);
    
    \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[4]\ : DFN1C0
      port map(D => \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\);
    
    \U50_PATTERNS/U4C_REGCROSS/LOCAL_REG_VAL[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119107, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_21, Q => \ELKS_STRT_ADDR[5]\);
    
    \U_ELK17_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118335, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_17, Q => 
        \U_ELK17_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]_net_1\);
    
    HIEFFPLA_INST_0_56455 : AOI1D
      port map(A => HIEFFPLA_NET_0_117432, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_SEL[3]_net_1\, C
         => \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[1]_net_1\, Y
         => HIEFFPLA_NET_0_116863);
    
    HIEFFPLA_INST_0_52542 : MX2
      port map(A => HIEFFPLA_NET_0_117490, B => 
        HIEFFPLA_NET_0_117486, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_2[3]\, Y => 
        HIEFFPLA_NET_0_117550);
    
    \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[5]\ : DFN1C0
      port map(D => \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\);
    
    \U_ELK13_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]\ : DFN1C0
      port map(D => \U_ELK13_CH/U_SLAVE_1ELK/Q[9]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]_net_1\);
    
    \U_ELK19_CH/U_SLAVE_1ELK/Q[3]\ : DFN1C0
      port map(D => \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/Q[3]_net_1\);
    
    \U50_PATTERNS/TFC_DINA[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119197, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_4, Q => \U50_PATTERNS/TFC_DINA[0]\);
    
    HIEFFPLA_INST_0_49154 : MX2
      port map(A => \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[2]_net_1\, B
         => \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\, S => 
        \BIT_OS_SEL[2]\, Y => HIEFFPLA_NET_0_118181);
    
    AFLSDF_INV_29 : INV
      port map(A => DCB_SALT_SEL_c, Y => \AFLSDF_INV_29\);
    
    \U50_PATTERNS/ELINK_ADDRA_2[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119992, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_21, Q => 
        \U50_PATTERNS/ELINK_ADDRA_2[7]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_2[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116364, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_18, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_2[3]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_20[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116465, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_13, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_20[2]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/RECD_SER_WORD[7]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_116897, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_30, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/RECD_SER_WORD[7]_net_1\);
    
    HIEFFPLA_INST_0_46738 : MX2
      port map(A => \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[3]_net_1\, 
        B => \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\, S => 
        \BIT_OS_SEL_5[2]\, Y => HIEFFPLA_NET_0_118620);
    
    HIEFFPLA_INST_0_61718 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_9[0]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_25[0]\, S
         => \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_3[4]_net_1\, 
        Y => HIEFFPLA_NET_0_116088);
    
    HIEFFPLA_INST_0_47925 : MX2
      port map(A => \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\, 
        B => \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\, S => 
        \BIT_OS_SEL_1[2]\, Y => HIEFFPLA_NET_0_118403);
    
    \U_ELK6_CH/U_SLAVE_1ELK/Q[9]\ : DFN1C0
      port map(D => \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/Q[9]_net_1\);
    
    \U0_200M_BUF/\\\\INBUF_LVDS[0]\\\\/U0/U2\ : IOPADN_IN
      port map(PAD => CLK200_N, N2POUT => 
        \U0_200M_BUF/\\\\INBUF_LVDS[0]\\\\/U0/U2_N2P\);
    
    HIEFFPLA_INST_0_49893 : MX2
      port map(A => \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[2]_net_1\, B
         => \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\, S => 
        \BIT_OS_SEL_6[2]\, Y => HIEFFPLA_NET_0_118047);
    
    \U50_PATTERNS/ELINK_ADDRA_16[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120036, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_8, Q => 
        \U50_PATTERNS/ELINK_ADDRA_16[3]\);
    
    HIEFFPLA_INST_0_53951 : AND3B
      port map(A => HIEFFPLA_NET_0_117237, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[0]_net_1\, C
         => \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_2[3]_net_1\, 
        Y => HIEFFPLA_NET_0_117328);
    
    HIEFFPLA_INST_0_55460 : MX2
      port map(A => HIEFFPLA_NET_0_116111, B => 
        HIEFFPLA_NET_0_116015, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[3]\, Y => 
        HIEFFPLA_NET_0_117034);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_7[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116603, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_14, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_7[0]\);
    
    HIEFFPLA_INST_0_56273 : NAND3C
      port map(A => HIEFFPLA_NET_0_116878, B => 
        HIEFFPLA_NET_0_116886, C => HIEFFPLA_NET_0_116894, Y => 
        HIEFFPLA_NET_0_116902);
    
    \U_ELK6_CH/U_SLAVE_1ELK/RECD_SER_WORD[5]\ : DFN1C0
      port map(D => \U_ELK6_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[5]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_6[5]\);
    
    \U_ELK5_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118017, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_2, Q => 
        \U_ELK5_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]_net_1\);
    
    HIEFFPLA_INST_0_42690 : NAND3B
      port map(A => \U50_PATTERNS/REG_ADDR[5]\, B => 
        \U50_PATTERNS/REG_ADDR[3]\, C => 
        \U50_PATTERNS/REG_STATE_0[5]_net_1\, Y => 
        HIEFFPLA_NET_0_119482);
    
    \U_ELK18_CH/U_ELK1_SERDAT_SOURCE/SERDAT[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118281, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_13, Q => 
        \U_ELK18_CH/ELK_TX_DAT[2]\);
    
    \U50_PATTERNS/ELINK_DINA_2[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119773, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_9, Q => 
        \U50_PATTERNS/ELINK_DINA_2[2]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[1]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_WRD_40M_FIXED[1]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_27, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[1]_net_1\);
    
    \U_ELK11_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL\ : DFN1C0
      port map(D => 
        \U_ELK11_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL_net_1\);
    
    HIEFFPLA_INST_0_53749 : AND2B
      port map(A => HIEFFPLA_NET_0_117391, B => 
        HIEFFPLA_NET_0_117392, Y => HIEFFPLA_NET_0_117359);
    
    \U50_PATTERNS/ELINK_ADDRA_8[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119946, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_8, Q => 
        \U50_PATTERNS/ELINK_ADDRA_8[5]\);
    
    \U_ELK7_CH/U_ELK1_SERDAT_SOURCE/SERDAT[5]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117918, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_3, Q => 
        \U_ELK7_CH/ELK_TX_DAT[5]\);
    
    AFLSDF_INV_27 : INV
      port map(A => DCB_SALT_SEL_c, Y => \AFLSDF_INV_27\);
    
    \U_ELK8_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117885, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]_net_1\);
    
    \U_ELK2_CH/U_SLAVE_1ELK/RECD_SER_WORD[2]\ : DFN1C0
      port map(D => \U_ELK2_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[2]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_2[2]\);
    
    HIEFFPLA_INST_0_56524 : AND3A
      port map(A => HIEFFPLA_NET_0_117430, B => \BIT_OS_SEL_1[2]\, 
        C => \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[8]_net_1\, 
        Y => HIEFFPLA_NET_0_116846);
    
    \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[47]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117725, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_18, Q => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[47]\);
    
    HIEFFPLA_INST_0_60711 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_15[0]\, B => 
        HIEFFPLA_NET_0_117190, S => HIEFFPLA_NET_0_117356, Y => 
        HIEFFPLA_NET_0_116230);
    
    HIEFFPLA_INST_0_45027 : NAND2A
      port map(A => \U50_PATTERNS/USB_TXE_B\, B => 
        \U50_PATTERNS/REG_STATE[4]_net_1\, Y => 
        HIEFFPLA_NET_0_118996);
    
    HIEFFPLA_INST_0_45947 : NAND3C
      port map(A => HIEFFPLA_NET_0_118950, B => 
        HIEFFPLA_NET_0_118958, C => HIEFFPLA_NET_0_118703, Y => 
        HIEFFPLA_NET_0_118804);
    
    HIEFFPLA_INST_0_41278 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_4[4]\, B => 
        HIEFFPLA_NET_0_119570, S => HIEFFPLA_NET_0_119284, Y => 
        HIEFFPLA_NET_0_119755);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_18[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116189, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_8, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_18[1]\);
    
    \U_ELK10_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]\ : DFN1C0
      port map(D => \U_ELK10_CH/U_SLAVE_1ELK/Q[11]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]_net_1\);
    
    \U_ELK6_CH/U_ELK1_SERDAT_SOURCE/SERDAT[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117965, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_1, Q => 
        \U_ELK6_CH/ELK_TX_DAT[3]\);
    
    \U_ELK18_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]\ : DFN1C0
      port map(D => \U_ELK18_CH/U_SLAVE_1ELK/Q[11]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]_net_1\);
    
    HIEFFPLA_INST_0_57264 : NAND3
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_3[3]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_3[2]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_3[1]\, Y => 
        HIEFFPLA_NET_0_116713);
    
    HIEFFPLA_INST_0_48365 : AND2
      port map(A => CLK_40M_GL, B => 
        \U_ELK17_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0_net_1\, Y => 
        HIEFFPLA_NET_0_118329);
    
    \U_ELK19_CH/U_SLAVE_1ELK/Q[1]\ : DFN1C0
      port map(D => \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/Q[1]_net_1\);
    
    \U50_PATTERNS/U4E_REGCROSS/DELCNT[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119046, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_25, Q => 
        \U50_PATTERNS/U4E_REGCROSS/DELCNT[1]_net_1\);
    
    HIEFFPLA_INST_0_52478 : MX2
      port map(A => HIEFFPLA_NET_0_117506, B => 
        HIEFFPLA_NET_0_117502, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[3]\, Y => 
        HIEFFPLA_NET_0_117558);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_6[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_115985, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_16, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_6[0]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_26[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116078, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_12, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_26[2]\);
    
    \U50_PATTERNS/U4B_REGCROSS/SAMP_ONE[2]\ : DFN1C0
      port map(D => \U50_PATTERNS/TFC_STOP_ADDR[2]\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_25, Q => 
        \U50_PATTERNS/U4B_REGCROSS/SAMP_ONE[2]_net_1\);
    
    \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[4]\ : DFN1C0
      port map(D => \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\);
    
    \U_TFC_SERDAT_SOURCE/SERDAT[0]\ : DFN1C0
      port map(D => \U_TFC_SERDAT_SOURCE/N_SERDAT[0]\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \TFC_TX_DAT[0]\);
    
    \U_ELK19_CH/U_ELK1_CMD_TX/START_RISE\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118239, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_8, Q => 
        \U_ELK19_CH/U_ELK1_CMD_TX/START_RISE_net_1\);
    
    \U_ELK13_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL\ : DFN1C0
      port map(D => 
        \U_ELK13_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL_net_1\);
    
    \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[5]\ : DFN1C0
      port map(D => \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\);
    
    HIEFFPLA_INST_0_43097 : NAND2
      port map(A => \U50_PATTERNS/REG_STATE[1]_net_1\, B => 
        \U50_PATTERNS/REG_STATE[0]_net_1\, Y => 
        HIEFFPLA_NET_0_119380);
    
    \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[5]\ : DFN1C0
      port map(D => \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\);
    
    HIEFFPLA_INST_0_43282 : MX2
      port map(A => \U50_PATTERNS/SI_CNT[1]\, B => 
        HIEFFPLA_NET_0_119326, S => HIEFFPLA_NET_0_119439, Y => 
        HIEFFPLA_NET_0_119333);
    
    HIEFFPLA_INST_0_42715 : AO1A
      port map(A => HIEFFPLA_NET_0_119451, B => 
        HIEFFPLA_NET_0_119455, C => HIEFFPLA_NET_0_119474, Y => 
        HIEFFPLA_NET_0_119476);
    
    HIEFFPLA_INST_0_43070 : AO1E
      port map(A => \U50_PATTERNS/REG_STATE[0]_net_1\, B => 
        HIEFFPLA_NET_0_119430, C => 
        \U50_PATTERNS/REG_STATE[3]_net_1\, Y => 
        HIEFFPLA_NET_0_119388);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_12[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116255, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_21, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_12[0]\);
    
    \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[6]\ : DFN1C0
      port map(D => 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\);
    
    HIEFFPLA_INST_0_44022 : MX2
      port map(A => \U50_PATTERNS/TFC_STOP_ADDR[5]\, B => 
        \U50_PATTERNS/TFC_STOP_ADDR_T[5]\, S => 
        HIEFFPLA_NET_0_119472, Y => HIEFFPLA_NET_0_119183);
    
    HIEFFPLA_INST_0_42931 : AO1A
      port map(A => HIEFFPLA_NET_0_119368, B => 
        HIEFFPLA_NET_0_119014, C => HIEFFPLA_NET_0_119406, Y => 
        HIEFFPLA_NET_0_119421);
    
    HIEFFPLA_INST_0_40972 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_19[2]\, B => 
        HIEFFPLA_NET_0_119575, S => HIEFFPLA_NET_0_119293, Y => 
        HIEFFPLA_NET_0_119789);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_21[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116454, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_14, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_21[2]\);
    
    \U_ELK5_CH/U_ELK1_SERDAT_SOURCE/SERDAT[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118013, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_17, Q => 
        \U_ELK5_CH/ELK_TX_DAT[0]\);
    
    HIEFFPLA_INST_0_111270 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_30[1]\, B => 
        HIEFFPLA_NET_0_116677, S => HIEFFPLA_NET_0_117328, Y => 
        HIEFFPLA_NET_0_116349);
    
    HIEFFPLA_INST_0_51908 : MX2
      port map(A => HIEFFPLA_NET_0_117660, B => 
        HIEFFPLA_NET_0_117659, S => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[5]\, Y => 
        HIEFFPLA_NET_0_117668);
    
    HIEFFPLA_INST_0_56238 : AND2
      port map(A => DCB_SALT_SEL_c, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/RECD_SER_WORD[2]_net_1\, 
        Y => \ELK_RX_SER_WORD_0[2]\);
    
    HIEFFPLA_INST_0_54908 : AOI1C
      port map(A => HIEFFPLA_NET_0_117184, B => 
        HIEFFPLA_NET_0_117388, C => HIEFFPLA_NET_0_117212, Y => 
        HIEFFPLA_NET_0_117173);
    
    HIEFFPLA_INST_0_51329 : AXOI7
      port map(A => \U_EXEC_MASTER/CCC_1_LOCK_STAT_1D_net_1\, B
         => HIEFFPLA_NET_0_117796, C => 
        \U_EXEC_MASTER/DEL_CNT[0]\, Y => HIEFFPLA_NET_0_117795);
    
    AFLSDF_INV_1 : INV
      port map(A => P_USB_MASTER_EN_c_22, Y => \AFLSDF_INV_1\);
    
    HIEFFPLA_INST_0_46724 : MX2
      port map(A => HIEFFPLA_NET_0_118635, B => 
        HIEFFPLA_NET_0_118631, S => \BIT_OS_SEL_5[1]\, Y => 
        HIEFFPLA_NET_0_118622);
    
    HIEFFPLA_INST_0_40115 : AOI1D
      port map(A => HIEFFPLA_NET_0_119389, B => 
        HIEFFPLA_NET_0_119464, C => \U50_PATTERNS/SM_BANK_SEL[3]\, 
        Y => HIEFFPLA_NET_0_119901);
    
    \U_ELK18_CH/U_SLAVE_1ELK/Q[10]\ : DFN1C0
      port map(D => \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/Q[10]_net_1\);
    
    \U_EXEC_MASTER/MPOR_B_7\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117787, CLK => CLK_40M_GL, CLR
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_1\, Q => 
        P_MASTER_POR_B_c_7);
    
    HIEFFPLA_INST_0_37041 : AO1A
      port map(A => HIEFFPLA_NET_0_120340, B => 
        HIEFFPLA_NET_0_120325, C => HIEFFPLA_NET_0_120345, Y => 
        HIEFFPLA_NET_0_120361);
    
    \U_ELK15_CH/U_SLAVE_1ELK/RECD_SER_WORD[1]\ : DFN1C0
      port map(D => \U_ELK15_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[1]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_15[1]\);
    
    \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[5]\ : DFN1C0
      port map(D => \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\);
    
    \U_ELK2_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]\ : DFN1C0
      port map(D => \U_ELK2_CH/U_SLAVE_1ELK/Q[14]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]_net_1\);
    
    \U_ELK15_CH/U_SLAVE_1ELK/Q[5]\ : DFN1C0
      port map(D => \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/Q[5]_net_1\);
    
    HIEFFPLA_INST_0_57658 : AO1A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_5[3]\, B => 
        HIEFFPLA_NET_0_116650, C => HIEFFPLA_NET_0_117179, Y => 
        HIEFFPLA_NET_0_116641);
    
    HIEFFPLA_INST_0_40270 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_0[4]\, B => 
        HIEFFPLA_NET_0_119570, S => HIEFFPLA_NET_0_119272, Y => 
        HIEFFPLA_NET_0_119867);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_13[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116250, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_1, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_13[0]\);
    
    HIEFFPLA_INST_0_41188 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_3[2]\, B => 
        HIEFFPLA_NET_0_119575, S => HIEFFPLA_NET_0_119247, Y => 
        HIEFFPLA_NET_0_119765);
    
    HIEFFPLA_INST_0_42661 : AND3C
      port map(A => HIEFFPLA_NET_0_119379, B => 
        \U50_PATTERNS/REG_STATE_0[5]_net_1\, C => 
        HIEFFPLA_NET_0_119017, Y => HIEFFPLA_NET_0_119489);
    
    HIEFFPLA_INST_0_37489 : MX2
      port map(A => \U200A_TFC/LOC_STRT_ADDR[6]\, B => 
        \TFC_STRT_ADDR[6]\, S => \U200A_TFC/GP_PG_SM_0[10]_net_1\, 
        Y => HIEFFPLA_NET_0_120276);
    
    HIEFFPLA_INST_0_47371 : NAND2B
      port map(A => \OP_MODE_c[1]\, B => \PATT_ELK_DAT_13[1]\, Y
         => HIEFFPLA_NET_0_118507);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_10[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116275, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_18, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_10[0]\);
    
    HIEFFPLA_INST_0_60858 : AND2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[4]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_16[0]\, Y => 
        HIEFFPLA_NET_0_116210);
    
    \U50_PATTERNS/ELINK_ADDRA_15[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120044, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_6, Q => 
        \U50_PATTERNS/ELINK_ADDRA_15[3]\);
    
    AFLSDF_INV_58 : INV
      port map(A => \U200B_ELINKS/RX_SER_WORD_2DEL[7]_net_1\, Y
         => \AFLSDF_INV_58\);
    
    \U_ELK12_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U1\ : IOBI_ID_OD_EB
      port map(DR => \U_ELK12_CH/ELK_OUT_R\, DF => 
        \U_ELK12_CH/ELK_OUT_F\, CLR => \GND\, E => 
        \AFLSDF_INV_18\, ICLK => CCC_160M_ADJ, OCLK => 
        CCC_160M_FXD, YIN => 
        \U_ELK12_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\, DOUT => 
        \U_ELK12_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, EOUT => 
        \U_ELK12_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET2\, YR => 
        \U_ELK12_CH/ELK_IN_DDR_R\, YF => 
        \U_ELK12_CH/ELK_IN_DDR_F\);
    
    HIEFFPLA_INST_0_50875 : MX2
      port map(A => HIEFFPLA_NET_0_117858, B => 
        HIEFFPLA_NET_0_117856, S => \BIT_OS_SEL_3[1]\, Y => 
        HIEFFPLA_NET_0_117869);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_1[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116170, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_8, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_1[0]\);
    
    \U200B_ELINKS/RX_SER_WORD_3DEL[0]\ : DFN1C0
      port map(D => \U200B_ELINKS/RX_SER_WORD_2DEL[0]_net_1\, CLK
         => CLK_40M_GL, CLR => P_MASTER_POR_B_c_31_0, Q => 
        \U200B_ELINKS/RX_SER_WORD_3DEL[0]_net_1\);
    
    \U_ELK7_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117925, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_11, Q => 
        \U_ELK7_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]_net_1\);
    
    \U_ELK15_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL\ : DFN1C0
      port map(D => 
        \U_ELK15_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL_net_1\);
    
    HIEFFPLA_INST_0_41889 : AND2
      port map(A => HIEFFPLA_NET_0_119389, B => 
        \U50_PATTERNS/SM_BANK_SEL[14]\, Y => 
        HIEFFPLA_NET_0_119673);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_17[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116205, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_6, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_17[0]\);
    
    \U50_PATTERNS/ELINK_DINA_17[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119800, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_19, Q => 
        \U50_PATTERNS/ELINK_DINA_17[7]\);
    
    HIEFFPLA_INST_0_37169 : AO1A
      port map(A => \OP_MODE_c[2]\, B => 
        \U200A_TFC/GP_PG_SM[0]_net_1\, C => HIEFFPLA_NET_0_120331, 
        Y => HIEFFPLA_NET_0_120335);
    
    HIEFFPLA_INST_0_37117 : AND3B
      port map(A => \U200A_TFC/LOC_STRT_ADDR[4]\, B => 
        HIEFFPLA_NET_0_120293, C => HIEFFPLA_NET_0_120328, Y => 
        HIEFFPLA_NET_0_120344);
    
    \U_ELK13_CH/U_SLAVE_1ELK/RECD_SER_WORD[6]\ : DFN1C0
      port map(D => \U_ELK13_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[6]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_13[6]\);
    
    \U50_PATTERNS/U4E_REGCROSS/SYNC_SM[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119055, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c, Q => 
        \U50_PATTERNS/U4E_REGCROSS/SYNC_SM[0]_net_1\);
    
    HIEFFPLA_INST_0_45136 : MX2
      port map(A => HIEFFPLA_NET_0_118969, B => 
        \U50_PATTERNS/WR_USB_ADBUS[6]\, S => 
        HIEFFPLA_NET_0_119486, Y => HIEFFPLA_NET_0_118979);
    
    HIEFFPLA_INST_0_57793 : NAND3
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_6[3]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_6[2]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_6[1]\, Y => 
        HIEFFPLA_NET_0_116621);
    
    HIEFFPLA_INST_0_46613 : MX2
      port map(A => 
        \U_ELK10_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]_net_1\, B => 
        \U_ELK10_CH/ELK_TX_DAT[5]\, S => 
        \U_ELK10_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118646);
    
    \U_ELK19_CH/U_SLAVE_1ELK/RECD_SER_WORD[3]\ : DFN1C0
      port map(D => \U_ELK19_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[3]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_19[3]\);
    
    HIEFFPLA_INST_0_41863 : AOI1B
      port map(A => HIEFFPLA_NET_0_119389, B => 
        \U50_PATTERNS/SM_BANK_SEL[0]\, C => HIEFFPLA_NET_0_119650, 
        Y => HIEFFPLA_NET_0_119680);
    
    \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[0]\ : DFN1C0
      port map(D => 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[0]_net_1\);
    
    HIEFFPLA_INST_0_54365 : MX2
      port map(A => HIEFFPLA_NET_0_116514, B => 
        HIEFFPLA_NET_0_116297, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_2[3]_net_1\, Y
         => HIEFFPLA_NET_0_117275);
    
    \U_ELK10_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U3\ : IOBI_ID_OD_EB
      port map(DR => \U_ELK10_CH/ELK_OUT_R\, DF => 
        \U_ELK10_CH/ELK_OUT_F\, CLR => \GND\, E => 
        \AFLSDF_INV_15\, ICLK => CCC_160M_ADJ, OCLK => 
        CCC_160M_FXD, YIN => 
        \U_ELK10_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\, DOUT => 
        OPEN, EOUT => 
        \U_ELK10_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET3\, YR => OPEN, 
        YF => OPEN);
    
    \U50_PATTERNS/U4C_REGCROSS/SAMP_TWO[2]\ : DFN1C0
      port map(D => \U50_PATTERNS/U4C_REGCROSS/SAMP_ONE[2]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_22_0, Q => 
        \U50_PATTERNS/U4C_REGCROSS/SAMP_TWO[2]_net_1\);
    
    HIEFFPLA_INST_0_61823 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_10[2]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_26[2]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_4[4]_net_1\, Y
         => HIEFFPLA_NET_0_116073);
    
    HIEFFPLA_INST_0_57822 : AND2A
      port map(A => HIEFFPLA_NET_0_116612, B => 
        HIEFFPLA_NET_0_116617, Y => HIEFFPLA_NET_0_116613);
    
    HIEFFPLA_INST_0_51515 : AX1
      port map(A => HIEFFPLA_NET_0_117755, B => 
        \U_EXEC_MASTER/PRESCALE[0]\, C => 
        \U_EXEC_MASTER/PRESCALE[3]\, Y => HIEFFPLA_NET_0_117757);
    
    HIEFFPLA_INST_0_42688 : AND3C
      port map(A => \U50_PATTERNS/REG_ADDR[7]\, B => 
        \U50_PATTERNS/REG_ADDR[6]\, C => HIEFFPLA_NET_0_119482, Y
         => HIEFFPLA_NET_0_119483);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_2[7]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116748, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_5, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_2[7]\);
    
    \U_ELK17_CH/U_SLAVE_1ELK/Q[5]\ : DFN1C0
      port map(D => \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/Q[5]_net_1\);
    
    HIEFFPLA_INST_0_56161 : NAND3C
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/MAX_CNT[8]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/MAX_CNT[7]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/MAX_CNT[6]\, Y => 
        HIEFFPLA_NET_0_116939);
    
    HIEFFPLA_INST_0_54749 : AND3A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[2]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[4]_net_1\, C => 
        HIEFFPLA_NET_0_117242, Y => HIEFFPLA_NET_0_117208);
    
    HIEFFPLA_INST_0_46923 : MX2
      port map(A => \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\, 
        B => \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[11]_net_1\, S => 
        \BIT_OS_SEL_4[2]\, Y => HIEFFPLA_NET_0_118584);
    
    HIEFFPLA_INST_0_50270 : MX2
      port map(A => HIEFFPLA_NET_0_117996, B => 
        HIEFFPLA_NET_0_117990, S => \BIT_OS_SEL_0[0]\, Y => 
        \U_ELK5_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[5]\);
    
    HIEFFPLA_INST_0_37499 : NAND2A
      port map(A => \U200A_TFC/RX_SER_WORD_2DEL[6]_net_1\, B => 
        \U200A_TFC/RX_SER_WORD_2DEL[7]_net_1\, Y => 
        HIEFFPLA_NET_0_120274);
    
    \U50_PATTERNS/ELINK_ADDRA_17[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120029, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_10, Q => 
        \U50_PATTERNS/ELINK_ADDRA_17[2]\);
    
    HIEFFPLA_INST_0_53278 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_SEQCNT[2]\, B => 
        HIEFFPLA_NET_0_117435, S => HIEFFPLA_NET_0_117062, Y => 
        HIEFFPLA_NET_0_117440);
    
    \U_ELK4_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL\ : DFN1C0
      port map(D => \U_ELK4_CH/ELK_IN_R_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL_net_1\);
    
    \U_ELK17_CH/U_SLAVE_1ELK/Q[7]\ : DFN1C0
      port map(D => \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/Q[7]_net_1\);
    
    HIEFFPLA_INST_0_48822 : MX2
      port map(A => \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\, 
        B => \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[14]_net_1\, S => 
        \BIT_OS_SEL_1[2]\, Y => HIEFFPLA_NET_0_118248);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_10[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116274, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_18, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_10[1]\);
    
    HIEFFPLA_INST_0_43751 : AND3A
      port map(A => \U50_PATTERNS/RD_USB_ADBUS[3]\, B => 
        HIEFFPLA_NET_0_119593, C => 
        \U50_PATTERNS/RD_USB_ADBUS[2]\, Y => 
        HIEFFPLA_NET_0_119223);
    
    HIEFFPLA_INST_0_41404 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_6[2]\, B => 
        HIEFFPLA_NET_0_119575, S => HIEFFPLA_NET_0_119258, Y => 
        HIEFFPLA_NET_0_119741);
    
    HIEFFPLA_INST_0_53561 : NAND3C
      port map(A => HIEFFPLA_NET_0_117350, B => 
        HIEFFPLA_NET_0_117070, C => HIEFFPLA_NET_0_117071, Y => 
        HIEFFPLA_NET_0_117388);
    
    HIEFFPLA_INST_0_48302 : MX2
      port map(A => HIEFFPLA_NET_0_118339, B => 
        HIEFFPLA_NET_0_118364, S => \BIT_OS_SEL_1[1]\, Y => 
        HIEFFPLA_NET_0_118341);
    
    HIEFFPLA_INST_0_40107 : AOI1C
      port map(A => \U50_PATTERNS/ELINK_BLKA[15]\, B => 
        HIEFFPLA_NET_0_119654, C => HIEFFPLA_NET_0_119903, Y => 
        HIEFFPLA_NET_0_119904);
    
    HIEFFPLA_INST_0_42529 : OA1A
      port map(A => HIEFFPLA_NET_0_119433, B => 
        HIEFFPLA_NET_0_119010, C => \U50_PATTERNS/REG_ADDR[3]\, Y
         => HIEFFPLA_NET_0_119520);
    
    \U_ELK12_CH/U_ELK1_CMD_TX/START_RISE\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118554, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_0, Q => 
        \U_ELK12_CH/U_ELK1_CMD_TX/START_RISE_net_1\);
    
    HIEFFPLA_INST_0_61643 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_8[2]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_24[2]\, S
         => \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_4[4]_net_1\, 
        Y => HIEFFPLA_NET_0_116098);
    
    \U50_PATTERNS/ELINK_DINA_4[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119759, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_12, Q => 
        \U50_PATTERNS/ELINK_DINA_4[0]\);
    
    HIEFFPLA_INST_0_59023 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_6[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_22[1]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_2[4]_net_1\, Y
         => HIEFFPLA_NET_0_116446);
    
    \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[11]\ : DFN1C0
      port map(D => \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\);
    
    \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[7]\ : DFN1C0
      port map(D => 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\);
    
    HIEFFPLA_INST_0_40087 : AO1A
      port map(A => HIEFFPLA_NET_0_119878, B => 
        \U50_PATTERNS/ELINK_BLKA[11]\, C => HIEFFPLA_NET_0_119910, 
        Y => HIEFFPLA_NET_0_119911);
    
    \U50_PATTERNS/U4A_REGCROSS/LOCAL_REG_VAL[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119152, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_17, Q => \TFC_STRT_ADDR[2]\);
    
    HIEFFPLA_INST_0_44368 : MX2
      port map(A => \TFC_STOP_ADDR[3]\, B => 
        \U50_PATTERNS/U4B_REGCROSS/SAMP_TWO[3]_net_1\, S => 
        HIEFFPLA_NET_0_119135, Y => HIEFFPLA_NET_0_119130);
    
    \U50_PATTERNS/SI_CNT[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119331, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_5, Q => \U50_PATTERNS/SI_CNT[3]\);
    
    \U_ELK1_CH/U_ELK1_CMD_TX/SER_OUT_RDEL\ : DFN1P0
      port map(D => \U_ELK1_CH/U_ELK1_CMD_TX/SER_OUT_RI_i\, CLK
         => CCC_160M_FXD, PRE => MASTER_SALT_POR_B_i_0_i_16, Q
         => \U_ELK1_CH/ELK_OUT_R_i_0\);
    
    HIEFFPLA_INST_0_37594 : AND3C
      port map(A => HIEFFPLA_NET_0_120238, B => 
        HIEFFPLA_NET_0_120241, C => HIEFFPLA_NET_0_120244, Y => 
        HIEFFPLA_NET_0_120251);
    
    \U_ELK4_CH/U_ELK1_SERDAT_SOURCE/SERDAT[5]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118053, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_16, Q => 
        \U_ELK4_CH/ELK_TX_DAT[5]\);
    
    \U50_PATTERNS/SI_CNT[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119334, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_5, Q => \U50_PATTERNS/SI_CNT[0]\);
    
    HIEFFPLA_INST_0_62094 : MX2
      port map(A => HIEFFPLA_NET_0_116139, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_29[0]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_2[3]\, Y => 
        HIEFFPLA_NET_0_116036);
    
    \U_ELK5_CH/U_SLAVE_1ELK/Q[0]\ : DFN1C0
      port map(D => \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/Q[0]_net_1\);
    
    HIEFFPLA_INST_0_56385 : AO1
      port map(A => HIEFFPLA_NET_0_117431, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[9]_net_1\, C => 
        HIEFFPLA_NET_0_116857, Y => HIEFFPLA_NET_0_116881);
    
    HIEFFPLA_INST_0_48599 : MX2
      port map(A => 
        \U_ELK18_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]_net_1\, B => 
        \U_ELK18_CH/ELK_TX_DAT[3]\, S => 
        \U_ELK18_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118287);
    
    HIEFFPLA_INST_0_43862 : MX2
      port map(A => HIEFFPLA_NET_0_119518, B => 
        \U50_PATTERNS/TFC_ADDRA[5]\, S => HIEFFPLA_NET_0_119294, 
        Y => HIEFFPLA_NET_0_119202);
    
    \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_2S_19\ : DFN1C0
      port map(D => 
        \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_1S_0_net_1\, CLK
         => CLK60MHZ, CLR => \U_EXEC_MASTER/P_MASTER_POR_B_c_0\, 
        Q => P_USB_MASTER_EN_c_19);
    
    \U200A_TFC/R_BLKB/U1\ : DFN1P0
      port map(D => HIEFFPLA_NET_0_120266, CLK => CLK_40M_GL, PRE
         => P_MASTER_POR_B_c_9, Q => TFC_RAM_BLKB_EN);
    
    \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[1]\ : DFN1C0
      port map(D => 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[1]_net_1\);
    
    HIEFFPLA_INST_0_38903 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_14[5]\, B => 
        HIEFFPLA_NET_0_119518, S => HIEFFPLA_NET_0_119249, Y => 
        HIEFFPLA_NET_0_120050);
    
    HIEFFPLA_INST_0_50855 : AND2
      port map(A => CLK_40M_GL, B => 
        \U_ELK8_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0_net_1\, Y => 
        HIEFFPLA_NET_0_117879);
    
    \U50_PATTERNS/U4E_REGCROSS/LOCAL_REG_VAL_0[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119062, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_1, Q => \OP_MODE_c_0[1]\);
    
    HIEFFPLA_INST_0_46576 : AND2A
      port map(A => \OP_MODE_c_4[1]\, B => \PATT_ELK_DAT_0[0]\, Y
         => HIEFFPLA_NET_0_118660);
    
    HIEFFPLA_INST_0_57542 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_5[1]\, B => 
        HIEFFPLA_NET_0_116644, S => HIEFFPLA_NET_0_117121, Y => 
        HIEFFPLA_NET_0_116660);
    
    HIEFFPLA_INST_0_46527 : AOI1A
      port map(A => HIEFFPLA_NET_0_119571, B => 
        HIEFFPLA_NET_0_119587, C => 
        \U50_PATTERNS/WR_XFER_TYPE[0]_net_1\, Y => 
        HIEFFPLA_NET_0_118672);
    
    \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[6]\ : DFN1C0
      port map(D => 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\);
    
    \U_ELK12_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118558, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_12, Q => 
        \U_ELK12_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]_net_1\);
    
    \U50_PATTERNS/ELINK_ADDRA_5[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119968, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_3, Q => 
        \U50_PATTERNS/ELINK_ADDRA_5[7]\);
    
    HIEFFPLA_INST_0_44190 : MX2
      port map(A => \U50_PATTERNS/TFC_STRT_ADDR_T[2]\, B => 
        \U50_PATTERNS/RD_USB_ADBUS[2]\, S => 
        HIEFFPLA_NET_0_119491, Y => HIEFFPLA_NET_0_119162);
    
    \U50_PATTERNS/ELINK_ADDRA_9[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119937, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_10, Q => 
        \U50_PATTERNS/ELINK_ADDRA_9[6]\);
    
    \U50_PATTERNS/ELINK_ADDRA_5[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119974, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_3, Q => 
        \U50_PATTERNS/ELINK_ADDRA_5[1]\);
    
    HIEFFPLA_INST_0_53935 : MX2
      port map(A => HIEFFPLA_NET_0_116191, B => 
        HIEFFPLA_NET_0_116086, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[3]_net_1\, Y
         => HIEFFPLA_NET_0_117331);
    
    HIEFFPLA_INST_0_37502 : OR3B
      port map(A => \U200A_TFC/RX_SER_WORD_2DEL[3]_net_1\, B => 
        \U200A_TFC/RX_SER_WORD_2DEL[2]_net_1\, C => 
        HIEFFPLA_NET_0_120272, Y => HIEFFPLA_NET_0_120273);
    
    \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[4]\ : DFN1C0
      port map(D => 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\);
    
    HIEFFPLA_INST_0_53770 : AND2
      port map(A => HIEFFPLA_NET_0_117414, B => 
        HIEFFPLA_NET_0_117359, Y => HIEFFPLA_NET_0_117354);
    
    HIEFFPLA_INST_0_49352 : MX2
      port map(A => 
        \U_ELK2_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]_net_1\, B => 
        \U_ELK2_CH/ELK_TX_DAT[5]\, S => 
        \U_ELK2_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118151);
    
    HIEFFPLA_INST_0_44616 : MX2B
      port map(A => HIEFFPLA_NET_0_119082, B => 
        HIEFFPLA_NET_0_119093, S => 
        \U50_PATTERNS/U4D_REGCROSS/SYNC_SM[0]_net_1\, Y => 
        HIEFFPLA_NET_0_119083);
    
    \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[5]\ : DFN1C0
      port map(D => 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\);
    
    HIEFFPLA_INST_0_51025 : MX2
      port map(A => HIEFFPLA_NET_0_117869, B => 
        HIEFFPLA_NET_0_117867, S => \BIT_OS_SEL_5[0]\, Y => 
        \U_ELK8_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[6]\);
    
    HIEFFPLA_INST_0_44310 : NAND3C
      port map(A => HIEFFPLA_NET_0_119142, B => 
        HIEFFPLA_NET_0_119143, C => HIEFFPLA_NET_0_119144, Y => 
        HIEFFPLA_NET_0_119145);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_25[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116419, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_20, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_25[1]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[4]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_115935, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_24_0, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[4]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_5[5]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116656, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_11, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_5[5]\);
    
    HIEFFPLA_INST_0_46172 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/SM_BANK_SEL[18]\, C => 
        \U50_PATTERNS/ELINK_DOUTA_1[3]\, Y => 
        HIEFFPLA_NET_0_118750);
    
    \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[9]\ : DFN1C0
      port map(D => 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\);
    
    HIEFFPLA_INST_0_47690 : MX2
      port map(A => HIEFFPLA_NET_0_118448, B => 
        HIEFFPLA_NET_0_118444, S => \BIT_OS_SEL_2[1]\, Y => 
        HIEFFPLA_NET_0_118446);
    
    \U_ELK1_CH/U_SLAVE_1ELK/Q[7]\ : DFN1C0
      port map(D => \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/Q[7]_net_1\);
    
    \U_ELK14_CH/U_ELK1_SERDAT_SOURCE/SERDAT[6]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118457, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_6, Q => 
        \U_ELK14_CH/ELK_TX_DAT[6]\);
    
    \U50_PATTERNS/ELINKS_STRT_ADDR_T[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120096, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_21, Q => 
        \U50_PATTERNS/ELINKS_STRT_ADDR_T[7]\);
    
    HIEFFPLA_INST_0_56852 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_1[3]\, B => 
        HIEFFPLA_NET_0_116765, S => HIEFFPLA_NET_0_117600, Y => 
        HIEFFPLA_NET_0_116785);
    
    HIEFFPLA_INST_0_53174 : MX2
      port map(A => HIEFFPLA_NET_0_117532, B => 
        HIEFFPLA_NET_0_117524, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_2[3]\, Y => 
        HIEFFPLA_NET_0_117456);
    
    HIEFFPLA_INST_0_47314 : MX2
      port map(A => HIEFFPLA_NET_0_118535, B => 
        HIEFFPLA_NET_0_118518, S => \BIT_OS_SEL_6[1]\, Y => 
        HIEFFPLA_NET_0_118520);
    
    \U_ELK8_CH/U_ELK1_SERDAT_SOURCE/SERDAT[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117876, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_5, Q => 
        \U_ELK8_CH/ELK_TX_DAT[2]\);
    
    HIEFFPLA_INST_0_44264 : MX2
      port map(A => \TFC_STRT_ADDR[3]\, B => 
        \U50_PATTERNS/U4A_REGCROSS/SAMP_TWO[3]_net_1\, S => 
        HIEFFPLA_NET_0_119156, Y => HIEFFPLA_NET_0_119151);
    
    HIEFFPLA_INST_0_51539 : AOI1A
      port map(A => 
        \U_EXEC_MASTER/USB_MASTER_EN/TEST_SM[3]_net_1\, B => 
        \U_EXEC_MASTER/USB_MASTER_EN/TEST_SM_i_0[2]\, C => 
        \U_EXEC_MASTER/USB_MASTER_EN/TERMCNT_FG40M2S_net_1\, Y
         => HIEFFPLA_NET_0_117750);
    
    \U_EXEC_MASTER/MPOR_SALT_B_2\ : DFI1P0
      port map(D => HIEFFPLA_NET_0_117781, CLK => CLK_40M_GL, PRE
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_2\, QN => 
        MASTER_SALT_POR_B_i_0_i_2);
    
    HIEFFPLA_INST_0_46125 : AO1
      port map(A => HIEFFPLA_NET_0_119250, B => 
        \U50_PATTERNS/ELINK_DOUTA_5[2]\, C => 
        HIEFFPLA_NET_0_118935, Y => HIEFFPLA_NET_0_118760);
    
    \U_ELK15_CH/U_SLAVE_1ELK/RECD_SER_WORD[5]\ : DFN1C0
      port map(D => \U_ELK15_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[5]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_15[5]\);
    
    HIEFFPLA_INST_0_54990 : AOI1D
      port map(A => HIEFFPLA_NET_0_117416, B => 
        HIEFFPLA_NET_0_116814, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_3[6]_net_1\, Y => 
        HIEFFPLA_NET_0_117147);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_5[4]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_115991, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_15, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_5[4]\);
    
    \U_ELK18_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL\ : DFN1C0
      port map(D => 
        \U_ELK18_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL_net_1\);
    
    AFLSDF_INV_40 : INV
      port map(A => DCB_SALT_SEL_c, Y => \AFLSDF_INV_40\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_1[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_115937, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_24_0, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_1[3]_net_1\);
    
    HIEFFPLA_INST_0_54580 : NAND3C
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[3]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[0]_net_1\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[1]_net_1\, Y => 
        HIEFFPLA_NET_0_117241);
    
    HIEFFPLA_INST_0_43183 : OA1A
      port map(A => \U50_PATTERNS/USB_RXF_B\, B => 
        \U50_PATTERNS/REG_STATE_0[2]_net_1\, C => 
        HIEFFPLA_NET_0_119351, Y => HIEFFPLA_NET_0_119353);
    
    HIEFFPLA_INST_0_56360 : AO1
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[4]_net_1\, B => 
        HIEFFPLA_NET_0_117431, C => HIEFFPLA_NET_0_116862, Y => 
        HIEFFPLA_NET_0_116886);
    
    HIEFFPLA_INST_0_52926 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_31[0]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_0[0]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_3[0]\, Y => 
        HIEFFPLA_NET_0_117488);
    
    HIEFFPLA_INST_0_44439 : XO1
      port map(A => \U50_PATTERNS/U4B_REGCROSS/SAMP_TWO[6]_net_1\, 
        B => \TFC_STOP_ADDR[6]\, C => HIEFFPLA_NET_0_119116, Y
         => HIEFFPLA_NET_0_119117);
    
    \U_ELK18_CH/ELK_IN_F\ : DFN1C0
      port map(D => \U_ELK18_CH/ELK_IN_DDR_F\, CLK => 
        CCC_160M_ADJ, CLR => DEV_RST_B_c, Q => 
        \U_ELK18_CH/ELK_IN_F_net_1\);
    
    \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[2]\ : DFN1C0
      port map(D => \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\);
    
    \U_ELK11_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118600, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_7, Q => 
        \U_ELK11_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]_net_1\);
    
    HIEFFPLA_INST_0_55476 : MX2
      port map(A => HIEFFPLA_NET_0_116108, B => 
        HIEFFPLA_NET_0_116013, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[3]\, Y => 
        HIEFFPLA_NET_0_117032);
    
    HIEFFPLA_INST_0_49863 : NAND2B
      port map(A => \OP_MODE_c_1[1]\, B => \PATT_ELK_DAT_4[3]\, Y
         => HIEFFPLA_NET_0_118055);
    
    HIEFFPLA_INST_0_40423 : MX2
      port map(A => HIEFFPLA_NET_0_119567, B => 
        \U50_PATTERNS/ELINK_DINA_11[5]\, S => 
        HIEFFPLA_NET_0_119280, Y => HIEFFPLA_NET_0_119850);
    
    \U_ELK19_CH/U_ELK1_SERDAT_SOURCE/SERDAT[6]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118232, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_15, Q => 
        \U_ELK19_CH/ELK_TX_DAT[6]\);
    
    HIEFFPLA_INST_0_50708 : MX2
      port map(A => \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\, B
         => \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[12]_net_1\, S => 
        \BIT_OS_SEL_4[2]\, Y => HIEFFPLA_NET_0_117902);
    
    \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[0]\ : DFN1C0
      port map(D => 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[0]_net_1\);
    
    HIEFFPLA_INST_0_37289 : AOI1B
      port map(A => HIEFFPLA_NET_0_120268, B => 
        HIEFFPLA_NET_0_120273, C => \U200A_TFC/GP_PG_SM[7]_net_1\, 
        Y => HIEFFPLA_NET_0_120304);
    
    HIEFFPLA_INST_0_51109 : AND2A
      port map(A => \OP_MODE_c_3[1]\, B => \PATT_ELK_DAT_9[4]\, Y
         => HIEFFPLA_NET_0_117829);
    
    HIEFFPLA_INST_0_55542 : AO1
      port map(A => HIEFFPLA_NET_0_117087, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_1[0]\, C => 
        HIEFFPLA_NET_0_116997, Y => HIEFFPLA_NET_0_117023);
    
    HIEFFPLA_INST_0_54109 : MX2
      port map(A => HIEFFPLA_NET_0_116138, B => 
        HIEFFPLA_NET_0_116244, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_1[3]_net_1\, Y
         => HIEFFPLA_NET_0_117307);
    
    HIEFFPLA_INST_0_42440 : AXOI4
      port map(A => HIEFFPLA_NET_0_119452, B => 
        HIEFFPLA_NET_0_119007, C => \U50_PATTERNS/REG_ADDR[0]\, Y
         => HIEFFPLA_NET_0_119533);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_2[4]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116751, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_5, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_2[4]\);
    
    \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[9]\ : DFN1C0
      port map(D => \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\);
    
    HIEFFPLA_INST_0_41413 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_6[3]\, B => 
        HIEFFPLA_NET_0_119574, S => HIEFFPLA_NET_0_119258, Y => 
        HIEFFPLA_NET_0_119740);
    
    \U_ELK13_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]\ : DFN1C0
      port map(D => \U_ELK13_CH/U_SLAVE_1ELK/Q[4]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]_net_1\);
    
    \U_ELK15_CH/ELK_IN_F\ : DFN1C0
      port map(D => \U_ELK15_CH/ELK_IN_DDR_F\, CLK => 
        CCC_160M_ADJ, CLR => DEV_RST_B_c, Q => 
        \U_ELK15_CH/ELK_IN_F_net_1\);
    
    \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_2S_7\ : DFN1C0
      port map(D => 
        \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_1S_net_1\, CLK
         => CLK60MHZ, CLR => P_MASTER_POR_B_c_0_0, Q => 
        P_USB_MASTER_EN_c_7);
    
    \U_ELK13_CH/U_ELK1_CMD_TX/START_RISE\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118509, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_9, Q => 
        \U_ELK13_CH/U_ELK1_CMD_TX/START_RISE_net_1\);
    
    HIEFFPLA_INST_0_55239 : AO1
      port map(A => HIEFFPLA_NET_0_115906, B => 
        HIEFFPLA_NET_0_117064, C => HIEFFPLA_NET_0_117124, Y => 
        HIEFFPLA_NET_0_117078);
    
    HIEFFPLA_INST_0_49017 : MX2
      port map(A => HIEFFPLA_NET_0_118223, B => 
        HIEFFPLA_NET_0_118221, S => \BIT_OS_SEL_2[0]\, Y => 
        \U_ELK19_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[4]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_19[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116478, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_20, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_19[3]\);
    
    HIEFFPLA_INST_0_55148 : NAND2B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[8]_net_1\, B => 
        HIEFFPLA_NET_0_117099, Y => HIEFFPLA_NET_0_117112);
    
    \U_EXEC_MASTER/USB_MASTER_EN/CNT_EN_40M\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117754, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_23, Q => 
        \U_EXEC_MASTER/USB_MASTER_EN/CNT_EN_40M_net_1\);
    
    \U_ELK8_CH/U_SLAVE_1ELK/RECD_SER_WORD[1]\ : DFN1C0
      port map(D => \U_ELK8_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[1]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_8[1]\);
    
    HIEFFPLA_INST_0_61184 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_1[3]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_2[3]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_1[0]\, Y => 
        HIEFFPLA_NET_0_116162);
    
    HIEFFPLA_INST_0_45954 : NAND3C
      port map(A => HIEFFPLA_NET_0_118852, B => 
        HIEFFPLA_NET_0_118702, C => HIEFFPLA_NET_0_118802, Y => 
        HIEFFPLA_NET_0_118803);
    
    \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[8]\ : DFN1C0
      port map(D => 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\);
    
    HIEFFPLA_INST_0_46243 : AO1
      port map(A => HIEFFPLA_NET_0_119476, B => 
        \U50_PATTERNS/CHKSUM[0]\, C => HIEFFPLA_NET_0_118905, Y
         => HIEFFPLA_NET_0_118733);
    
    HIEFFPLA_INST_0_45055 : MX2
      port map(A => USB_WR_BI, B => HIEFFPLA_NET_0_119486, S => 
        HIEFFPLA_NET_0_118989, Y => HIEFFPLA_NET_0_118990);
    
    HIEFFPLA_INST_0_42367 : AND3
      port map(A => HIEFFPLA_NET_0_119584, B => 
        HIEFFPLA_NET_0_119554, C => HIEFFPLA_NET_0_119552, Y => 
        HIEFFPLA_NET_0_119553);
    
    \U_ELK14_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]\ : DFN1C0
      port map(D => \U_ELK14_CH/U_SLAVE_1ELK/Q[6]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]_net_1\);
    
    HIEFFPLA_INST_0_58996 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_22[1]\, B => 
        HIEFFPLA_NET_0_116677, S => HIEFFPLA_NET_0_117095, Y => 
        HIEFFPLA_NET_0_116449);
    
    HIEFFPLA_INST_0_63077 : XA1B
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[13]\, 
        B => HIEFFPLA_NET_0_115883, C => HIEFFPLA_NET_0_117078, Y
         => HIEFFPLA_NET_0_115894);
    
    HIEFFPLA_INST_0_47931 : MX2
      port map(A => HIEFFPLA_NET_0_118410, B => 
        HIEFFPLA_NET_0_118408, S => \BIT_OS_SEL_2[1]\, Y => 
        HIEFFPLA_NET_0_118402);
    
    HIEFFPLA_INST_0_59829 : NAND2B
      port map(A => HIEFFPLA_NET_0_116708, B => 
        HIEFFPLA_NET_0_116813, Y => HIEFFPLA_NET_0_116345);
    
    HIEFFPLA_INST_0_45742 : AO1
      port map(A => HIEFFPLA_NET_0_119250, B => 
        \U50_PATTERNS/ELINK_DOUTA_5[7]\, C => 
        HIEFFPLA_NET_0_118782, Y => HIEFFPLA_NET_0_118854);
    
    HIEFFPLA_INST_0_41985 : AND3C
      port map(A => HIEFFPLA_NET_0_119271, B => 
        HIEFFPLA_NET_0_119262, C => \U50_PATTERNS/SM_BANK_SEL[6]\, 
        Y => HIEFFPLA_NET_0_119637);
    
    \U_ELK14_CH/U_SLAVE_1ELK/RECD_SER_WORD[5]\ : DFN1C0
      port map(D => \U_ELK14_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[5]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_14[5]\);
    
    HIEFFPLA_INST_0_55275 : AO1
      port map(A => HIEFFPLA_NET_0_117129, B => 
        HIEFFPLA_NET_0_116814, C => HIEFFPLA_NET_0_117076, Y => 
        HIEFFPLA_NET_0_117072);
    
    HIEFFPLA_INST_0_47869 : NAND2B
      port map(A => \OP_MODE_c_6[1]\, B => \PATT_ELK_DAT_15[1]\, 
        Y => HIEFFPLA_NET_0_118417);
    
    HIEFFPLA_INST_0_39980 : MX2
      port map(A => HIEFFPLA_NET_0_119904, B => 
        \U50_PATTERNS/ELINK_BLKA[15]\, S => 
        \U50_PATTERNS/SM_BANK_SEL[20]\, Y => 
        HIEFFPLA_NET_0_119929);
    
    HIEFFPLA_INST_0_48559 : MX2
      port map(A => HIEFFPLA_NET_0_118309, B => 
        HIEFFPLA_NET_0_118293, S => \BIT_OS_SEL_2[1]\, Y => 
        HIEFFPLA_NET_0_118295);
    
    \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117059, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_26, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[2]_net_1\);
    
    HIEFFPLA_INST_0_51706 : NAND2B
      port map(A => 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM[4]_net_1\, B => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[10]_net_1\, Y => 
        HIEFFPLA_NET_0_117720);
    
    \U200A_TFC/GP_PG_SM[7]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120312, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_28, Q => 
        \U200A_TFC/GP_PG_SM[7]_net_1\);
    
    HIEFFPLA_INST_0_58467 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_15[2]\, B => 
        HIEFFPLA_NET_0_116687, S => HIEFFPLA_NET_0_117098, Y => 
        HIEFFPLA_NET_0_116518);
    
    HIEFFPLA_INST_0_55060 : AND2A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[8]_net_1\, B => 
        HIEFFPLA_NET_0_115867, Y => HIEFFPLA_NET_0_117131);
    
    HIEFFPLA_INST_0_48013 : MX2
      port map(A => HIEFFPLA_NET_0_118395, B => 
        HIEFFPLA_NET_0_118407, S => \BIT_OS_SEL_3[0]\, Y => 
        \U_ELK15_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[3]\);
    
    HIEFFPLA_INST_0_38516 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_0[2]\, B => 
        HIEFFPLA_NET_0_119522, S => HIEFFPLA_NET_0_119272, Y => 
        HIEFFPLA_NET_0_120093);
    
    HIEFFPLA_INST_0_40064 : MX2
      port map(A => HIEFFPLA_NET_0_119882, B => 
        \U50_PATTERNS/ELINK_BLKA[8]\, S => 
        \U50_PATTERNS/SM_BANK_SEL[20]\, Y => 
        HIEFFPLA_NET_0_119917);
    
    HIEFFPLA_INST_0_111910 : AND3B
      port map(A => HIEFFPLA_NET_0_115822, B => 
        HIEFFPLA_NET_0_115823, C => HIEFFPLA_NET_0_119446, Y => 
        HIEFFPLA_NET_0_119631);
    
    HIEFFPLA_INST_0_38362 : MX2
      port map(A => \U50_PATTERNS/ELINKS_STOP_ADDR_T[7]\, B => 
        \U50_PATTERNS/RD_USB_ADBUS[7]\, S => 
        HIEFFPLA_NET_0_119413, Y => HIEFFPLA_NET_0_120112);
    
    \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[14]\ : DFN1C0
      port map(D => 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]_net_1\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[14]_net_1\);
    
    HIEFFPLA_INST_0_48061 : MX2
      port map(A => HIEFFPLA_NET_0_118398, B => 
        HIEFFPLA_NET_0_118383, S => \BIT_OS_SEL_4[1]\, Y => 
        HIEFFPLA_NET_0_118385);
    
    \U_ELK15_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]\ : DFN1C0
      port map(D => \U_ELK15_CH/U_SLAVE_1ELK/Q[5]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]_net_1\);
    
    \U_ELK19_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0\ : DFN1C0
      port map(D => CLK_40M_GL, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_10, Q => 
        \U_ELK19_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0_net_1\);
    
    HIEFFPLA_INST_0_54450 : AO1E
      port map(A => HIEFFPLA_NET_0_116708, B => 
        HIEFFPLA_NET_0_116740, C => HIEFFPLA_NET_0_117208, Y => 
        HIEFFPLA_NET_0_117264);
    
    \U_ELK6_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]\ : DFN1C0
      port map(D => \U_ELK6_CH/U_SLAVE_1ELK/Q[1]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]_net_1\);
    
    \U50_PATTERNS/ELINK_ADDRA_19[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120012, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_13, Q => 
        \U50_PATTERNS/ELINK_ADDRA_19[3]\);
    
    HIEFFPLA_INST_0_51986 : AND2A
      port map(A => HIEFFPLA_NET_0_117647, B => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[6]\, Y => 
        HIEFFPLA_NET_0_117657);
    
    HIEFFPLA_INST_0_58163 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_10[2]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_26[2]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_2[4]_net_1\, Y
         => HIEFFPLA_NET_0_116556);
    
    HIEFFPLA_INST_0_53006 : MX2
      port map(A => HIEFFPLA_NET_0_117461, B => 
        HIEFFPLA_NET_0_117457, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[2]\, Y => 
        HIEFFPLA_NET_0_117477);
    
    HIEFFPLA_INST_0_55139 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[8]_net_1\, B => 
        HIEFFPLA_NET_0_117321, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[6]_net_1\, Y => 
        HIEFFPLA_NET_0_117115);
    
    HIEFFPLA_INST_0_52470 : MX2
      port map(A => HIEFFPLA_NET_0_117507, B => 
        HIEFFPLA_NET_0_117503, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[3]\, Y => 
        HIEFFPLA_NET_0_117559);
    
    HIEFFPLA_INST_0_40729 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_15[7]\, B => 
        HIEFFPLA_NET_0_119560, S => HIEFFPLA_NET_0_119297, Y => 
        HIEFFPLA_NET_0_119816);
    
    HIEFFPLA_INST_0_49899 : MX2
      port map(A => \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[3]_net_1\, B
         => \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\, S => 
        \BIT_OS_SEL_6[2]\, Y => HIEFFPLA_NET_0_118046);
    
    \U_ELK7_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117931, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_14, Q => 
        \U_ELK7_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]_net_1\);
    
    HIEFFPLA_INST_0_45370 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/SM_BANK_SEL[2]\, C => 
        \U50_PATTERNS/ELINK_DOUTA_17[1]\, Y => 
        HIEFFPLA_NET_0_118928);
    
    \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[13]\ : DFN1C0
      port map(D => 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[13]_net_1\);
    
    \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[12]\ : DFN1C0
      port map(D => \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\, 
        CLK => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\);
    
    HIEFFPLA_INST_0_40621 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_14[3]\, B => 
        HIEFFPLA_NET_0_119574, S => HIEFFPLA_NET_0_119249, Y => 
        HIEFFPLA_NET_0_119828);
    
    \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[7]\ : DFN1C0
      port map(D => \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_6[5]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116627, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_12, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_6[5]\);
    
    \U_ELK6_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]\ : DFN1C0
      port map(D => \U_ELK6_CH/U_SLAVE_1ELK/Q[11]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]_net_1\);
    
    \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[14]\ : DFN1C0
      port map(D => \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\, 
        CLK => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[14]_net_1\);
    
    \U_ELK12_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]\ : DFN1C0
      port map(D => \U_ELK12_CH/U_SLAVE_1ELK/Q[5]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]_net_1\);
    
    \U_ELK10_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]\ : DFN1C0
      port map(D => \U_ELK10_CH/U_SLAVE_1ELK/Q[3]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]_net_1\);
    
    HIEFFPLA_INST_0_54874 : NAND3C
      port map(A => HIEFFPLA_NET_0_117191, B => 
        HIEFFPLA_NET_0_117189, C => HIEFFPLA_NET_0_117067, Y => 
        HIEFFPLA_NET_0_117184);
    
    HIEFFPLA_INST_0_54546 : AND2A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[3]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[0]_net_1\, Y => 
        HIEFFPLA_NET_0_117251);
    
    HIEFFPLA_INST_0_51226 : MX2
      port map(A => HIEFFPLA_NET_0_117801, B => 
        HIEFFPLA_NET_0_117824, S => \BIT_OS_SEL_4[0]\, Y => 
        \U_ELK9_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[0]\);
    
    HIEFFPLA_INST_0_43104 : AND3C
      port map(A => \U50_PATTERNS/REG_STATE[2]_net_1\, B => 
        \U50_PATTERNS/REG_STATE[0]_net_1\, C => 
        \U50_PATTERNS/REG_STATE[1]_net_1\, Y => 
        HIEFFPLA_NET_0_119375);
    
    HIEFFPLA_INST_0_41611 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_9[1]\, B => 
        HIEFFPLA_NET_0_119576, S => HIEFFPLA_NET_0_119292, Y => 
        HIEFFPLA_NET_0_119718);
    
    \U_ELK7_CH/U_ELK1_CMD_TX/START_RISE\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117924, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_2, Q => 
        \U_ELK7_CH/U_ELK1_CMD_TX/START_RISE_net_1\);
    
    HIEFFPLA_INST_0_56890 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_1[7]\, B => 
        HIEFFPLA_NET_0_116760, S => HIEFFPLA_NET_0_117600, Y => 
        HIEFFPLA_NET_0_116781);
    
    HIEFFPLA_INST_0_49367 : AND2A
      port map(A => \OP_MODE_c_1[1]\, B => \PATT_ELK_DAT_2[5]\, Y
         => HIEFFPLA_NET_0_118143);
    
    HIEFFPLA_INST_0_44321 : XO1
      port map(A => \U50_PATTERNS/U4A_REGCROSS/SAMP_TWO[3]_net_1\, 
        B => \TFC_STRT_ADDR[3]\, C => HIEFFPLA_NET_0_119139, Y
         => HIEFFPLA_NET_0_119143);
    
    \U_TFC_CMD_TX/SER_CMD_WORD_F[3]\ : DFN1C0
      port map(D => \U_TFC_CMD_TX/N_SER_CMD_WORD_F[3]\, CLK => 
        CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_TFC_CMD_TX/SER_CMD_WORD_F[3]_net_1\);
    
    \U_ELK3_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL\ : DFN1C0
      port map(D => \U_ELK3_CH/ELK_IN_F_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL_net_1\);
    
    HIEFFPLA_INST_0_48955 : MX2
      port map(A => \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[2]_net_1\, 
        B => \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\, S => 
        \BIT_OS_SEL[2]\, Y => HIEFFPLA_NET_0_118219);
    
    HIEFFPLA_INST_0_59676 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_2[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_18[1]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_1[4]_net_1\, Y
         => HIEFFPLA_NET_0_116363);
    
    \U50_PATTERNS/U4D_REGCROSS/LOCAL_REG_VAL[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119086, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_3, Q => \ELKS_STOP_ADDR[5]\);
    
    HIEFFPLA_INST_0_59844 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_31[0]\, B => 
        HIEFFPLA_NET_0_116680, S => HIEFFPLA_NET_0_117097, Y => 
        HIEFFPLA_NET_0_116343);
    
    \U50_PATTERNS/ELINK_ADDRA_4[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119976, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_2_0, Q => 
        \U50_PATTERNS/ELINK_ADDRA_4[7]\);
    
    HIEFFPLA_INST_0_43724 : NAND2B
      port map(A => HIEFFPLA_NET_0_119230, B => 
        \U50_PATTERNS/SM_BANK_SEL[2]\, Y => HIEFFPLA_NET_0_119231);
    
    HIEFFPLA_INST_0_43585 : NAND3C
      port map(A => \U50_PATTERNS/SM_BANK_SEL[12]\, B => 
        \U50_PATTERNS/SM_BANK_SEL[13]\, C => 
        HIEFFPLA_NET_0_119287, Y => HIEFFPLA_NET_0_119279);
    
    \U_ELK11_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]\ : DFN1C0
      port map(D => \U_ELK11_CH/U_SLAVE_1ELK/Q[13]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_1[6]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117099, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_27_1, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_1[6]_net_1\);
    
    HIEFFPLA_INST_0_44742 : MX2
      port map(A => \OP_MODE_c_4[1]\, B => 
        \U50_PATTERNS/U4E_REGCROSS/SAMP_TWO[1]_net_1\, S => 
        HIEFFPLA_NET_0_119072, Y => HIEFFPLA_NET_0_119058);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_0[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116569, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_15, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_0[3]\);
    
    HIEFFPLA_INST_0_52794 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_11[2]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_12[2]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_1[0]\, Y => 
        HIEFFPLA_NET_0_117510);
    
    HIEFFPLA_INST_0_51082 : MX2
      port map(A => 
        \U_ELK9_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]_net_1\, B => 
        \U_ELK9_CH/ELK_TX_DAT[6]\, S => 
        \U_ELK9_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_117839);
    
    HIEFFPLA_INST_0_48967 : MX2
      port map(A => \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[3]_net_1\, 
        B => \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\, S => 
        \BIT_OS_SEL[2]\, Y => HIEFFPLA_NET_0_118217);
    
    HIEFFPLA_INST_0_42892 : AO1E
      port map(A => HIEFFPLA_NET_0_119454, B => 
        HIEFFPLA_NET_0_119389, C => HIEFFPLA_NET_0_119632, Y => 
        HIEFFPLA_NET_0_119433);
    
    \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[0]\ : DFN1C0
      port map(D => 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[0]_net_1\);
    
    \U_ELK2_CH/U_ELK1_SERDAT_SOURCE/SERDAT[5]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118143, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_13, Q => 
        \U_ELK2_CH/ELK_TX_DAT[5]\);
    
    HIEFFPLA_INST_0_56100 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/MAX_CNT[4]\, 
        B => HIEFFPLA_NET_0_116935, S => HIEFFPLA_NET_0_117084, Y
         => HIEFFPLA_NET_0_116950);
    
    HIEFFPLA_INST_0_42844 : NAND3B
      port map(A => \U50_PATTERNS/REG_STATE[1]_net_1\, B => 
        \U50_PATTERNS/REG_STATE[3]_net_1\, C => 
        \U50_PATTERNS/REG_STATE[2]_net_1\, Y => 
        HIEFFPLA_NET_0_119449);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_30[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116030, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_7, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_30[0]\);
    
    HIEFFPLA_INST_0_55655 : AND3B
      port map(A => HIEFFPLA_NET_0_117168, B => 
        HIEFFPLA_NET_0_117087, C => HIEFFPLA_NET_0_117027, Y => 
        HIEFFPLA_NET_0_117008);
    
    \U_ELK17_CH/U_ELK1_SERDAT_SOURCE/SERDAT[4]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118324, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_11, Q => 
        \U_ELK17_CH/ELK_TX_DAT[4]\);
    
    \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[2]\ : DFN1C0
      port map(D => 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[2]_net_1\);
    
    HIEFFPLA_INST_0_61748 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_25[4]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_26[4]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_4[0]\, Y => 
        HIEFFPLA_NET_0_116083);
    
    \U50_PATTERNS/TFC_STRT_ADDR_T[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119157, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_5, Q => 
        \U50_PATTERNS/TFC_STRT_ADDR_T[7]\);
    
    \U50_PATTERNS/ELINK_DINA_17[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119801, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_19, Q => 
        \U50_PATTERNS/ELINK_DINA_17[6]\);
    
    \U_EXEC_MASTER/MPOR_B_16_0\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117787, CLK => CLK_40M_GL, CLR
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_0\, Q => 
        P_MASTER_POR_B_c_16_0);
    
    HIEFFPLA_INST_0_37045 : AOI1A
      port map(A => \TFC_STRT_ADDR[4]\, B => 
        HIEFFPLA_NET_0_120349, C => HIEFFPLA_NET_0_120359, Y => 
        HIEFFPLA_NET_0_120360);
    
    HIEFFPLA_INST_0_111275 : NAND3C
      port map(A => HIEFFPLA_NET_0_116774, B => 
        HIEFFPLA_NET_0_116740, C => HIEFFPLA_NET_0_116345, Y => 
        HIEFFPLA_NET_0_115844);
    
    HIEFFPLA_INST_0_56737 : NAND3C
      port map(A => HIEFFPLA_NET_0_116768, B => 
        HIEFFPLA_NET_0_117370, C => HIEFFPLA_NET_0_116811, Y => 
        HIEFFPLA_NET_0_116812);
    
    \U50_PATTERNS/U4C_REGCROSS/SAMP_ONE[3]\ : DFN1C0
      port map(D => \U50_PATTERNS/ELINKS_STRT_ADDR[3]\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_33, Q => 
        \U50_PATTERNS/U4C_REGCROSS/SAMP_ONE[3]_net_1\);
    
    HIEFFPLA_INST_0_52142 : NAND2B
      port map(A => 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM[3]_net_1\, B => 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM[1]_net_1\, Y => 
        HIEFFPLA_NET_0_117627);
    
    \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[12]\ : DFN1C0
      port map(D => \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\, 
        CLK => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\);
    
    HIEFFPLA_INST_0_56748 : NAND2A
      port map(A => HIEFFPLA_NET_0_116802, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_0[0]\, Y => 
        HIEFFPLA_NET_0_116809);
    
    \U50_PATTERNS/WR_USB_ADBUS[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118979, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_15, Q => 
        \U50_PATTERNS/WR_USB_ADBUS[6]\);
    
    HIEFFPLA_INST_0_54496 : MX2
      port map(A => HIEFFPLA_NET_0_116470, B => 
        HIEFFPLA_NET_0_116280, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[3]_net_1\, Y => 
        HIEFFPLA_NET_0_117258);
    
    HIEFFPLA_INST_0_46628 : AND2A
      port map(A => \OP_MODE_c_3[1]\, B => \PATT_ELK_DAT_10[5]\, 
        Y => HIEFFPLA_NET_0_118638);
    
    \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[7]\ : DFN1C0
      port map(D => 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\);
    
    HIEFFPLA_INST_0_59835 : MX2B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_30[3]\, B => 
        HIEFFPLA_NET_0_116774, S => HIEFFPLA_NET_0_117328, Y => 
        HIEFFPLA_NET_0_116344);
    
    HIEFFPLA_INST_0_56407 : NAND3C
      port map(A => HIEFFPLA_NET_0_116826, B => 
        HIEFFPLA_NET_0_116842, C => HIEFFPLA_NET_0_116850, Y => 
        HIEFFPLA_NET_0_116874);
    
    HIEFFPLA_INST_0_43801 : AND3
      port map(A => HIEFFPLA_NET_0_119594, B => 
        \U50_PATTERNS/RD_USB_ADBUS[2]\, C => 
        \U50_PATTERNS/RD_USB_ADBUS[3]\, Y => 
        HIEFFPLA_NET_0_119211);
    
    \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[10]\ : DFN1C0
      port map(D => \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\);
    
    \U_ELK9_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]\ : DFN1C0
      port map(D => \U_ELK9_CH/U_SLAVE_1ELK/Q[12]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]_net_1\);
    
    HIEFFPLA_INST_0_40071 : MX2
      port map(A => HIEFFPLA_NET_0_119880, B => 
        \U50_PATTERNS/ELINK_BLKA[9]\, S => 
        \U50_PATTERNS/SM_BANK_SEL[20]\, Y => 
        HIEFFPLA_NET_0_119916);
    
    \U50_PATTERNS/ELINK_RWA[5]/U1\ : DFN1P0
      port map(D => HIEFFPLA_NET_0_119696, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_6, Q => \U50_PATTERNS/ELINK_RWA[5]\);
    
    HIEFFPLA_INST_0_51568 : AX1C
      port map(A => 
        \U_EXEC_MASTER/USB_MASTER_EN/T_CNT60M[0]_net_1\, B => 
        HIEFFPLA_NET_0_117753, C => HIEFFPLA_NET_0_117735, Y => 
        HIEFFPLA_NET_0_117742);
    
    \U_ELK16_CH/U_ELK1_SERDAT_SOURCE/SERDAT[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118371, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_9, Q => 
        \U_ELK16_CH/ELK_TX_DAT[2]\);
    
    \U_ELK13_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118511, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_16, Q => 
        \U_ELK13_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]_net_1\);
    
    \U50_PATTERNS/U4E_REGCROSS/LOCAL_REG_VAL[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119069, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_6, Q => \OP_MODE_c[1]\);
    
    HIEFFPLA_INST_0_45030 : AND3B
      port map(A => HIEFFPLA_NET_0_119379, B => 
        HIEFFPLA_NET_0_118996, C => HIEFFPLA_NET_0_119430, Y => 
        HIEFFPLA_NET_0_118994);
    
    HIEFFPLA_INST_0_44543 : XO1
      port map(A => \U50_PATTERNS/U4C_REGCROSS/SAMP_TWO[6]_net_1\, 
        B => \ELKS_STRT_ADDR[6]\, C => HIEFFPLA_NET_0_119095, Y
         => HIEFFPLA_NET_0_119096);
    
    HIEFFPLA_INST_0_40136 : AOI1D
      port map(A => HIEFFPLA_NET_0_119389, B => 
        HIEFFPLA_NET_0_119464, C => 
        \U50_PATTERNS/SM_BANK_SEL[18]\, Y => 
        HIEFFPLA_NET_0_119895);
    
    \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[2]\ : DFN1C0
      port map(D => 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[2]_net_1\);
    
    HIEFFPLA_INST_0_46001 : AND3B
      port map(A => HIEFFPLA_NET_0_119426, B => 
        HIEFFPLA_NET_0_119379, C => \U50_PATTERNS/OP_MODE[3]\, Y
         => HIEFFPLA_NET_0_118791);
    
    \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[7]\ : DFN1C0
      port map(D => 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\);
    
    \U_ELK10_CH/U_SLAVE_1ELK/RECD_SER_WORD[1]\ : DFN1C0
      port map(D => \U_ELK10_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[1]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_10[1]\);
    
    HIEFFPLA_INST_0_52394 : MX2
      port map(A => HIEFFPLA_NET_0_117525, B => 
        HIEFFPLA_NET_0_117481, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[1]\, Y => 
        HIEFFPLA_NET_0_117569);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_29[4]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116041, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_16_0, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_29[4]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[8]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_115922, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_9, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[8]\);
    
    \U_ELK15_CH/U_ELK1_CMD_TX/START_RISE\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118419, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_9, Q => 
        \U_ELK15_CH/U_ELK1_CMD_TX/START_RISE_net_1\);
    
    HIEFFPLA_INST_0_49483 : MX2
      port map(A => HIEFFPLA_NET_0_118116, B => 
        HIEFFPLA_NET_0_118126, S => \BIT_OS_SEL_1[0]\, Y => 
        \U_ELK2_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[0]\);
    
    \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[11]\ : DFN1C0
      port map(D => \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\);
    
    HIEFFPLA_INST_0_51882 : NAND2B
      port map(A => \U_MASTER_DES/AUX_MODE\, B => 
        HIEFFPLA_NET_0_117625, Y => HIEFFPLA_NET_0_117671);
    
    \U_ELK10_CH/U_ELK1_SERDAT_SOURCE/SERDAT[5]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118638, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_17, Q => 
        \U_ELK10_CH/ELK_TX_DAT[5]\);
    
    HIEFFPLA_INST_0_60048 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_5[0]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_21[0]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_5[4]_net_1\, Y
         => HIEFFPLA_NET_0_116317);
    
    AFLSDF_INV_67 : INV
      port map(A => \U200B_ELINKS/RX_SER_WORD_2DEL[2]_net_1\, Y
         => \AFLSDF_INV_67\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_22[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116447, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_15, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_22[3]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_30[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116029, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_7, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_30[1]\);
    
    \U_ELK1_CH/U_SLAVE_1ELK/Q[14]\ : DFN1C0
      port map(D => \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[14]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/Q[14]_net_1\);
    
    \U_ELK13_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118513, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_16, Q => 
        \U_ELK13_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]_net_1\);
    
    HIEFFPLA_INST_0_55421 : AO1
      port map(A => HIEFFPLA_NET_0_117087, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[0]\, C => 
        HIEFFPLA_NET_0_116997, Y => HIEFFPLA_NET_0_117040);
    
    HIEFFPLA_INST_0_51208 : MX2
      port map(A => \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\, B
         => \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\, S => 
        \BIT_OS_SEL_2[2]\, Y => HIEFFPLA_NET_0_117812);
    
    HIEFFPLA_INST_0_43461 : MX2
      port map(A => \U50_PATTERNS/SM_BANK_SEL[2]\, B => 
        HIEFFPLA_NET_0_119216, S => HIEFFPLA_NET_0_118691, Y => 
        HIEFFPLA_NET_0_119308);
    
    \U_ELK15_CH/U_ELK1_CMD_TX/SER_OUT_FDEL\ : DFN1C0
      port map(D => \U_ELK15_CH/U_ELK1_CMD_TX/SER_OUT_FI_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_8, Q
         => \U_ELK15_CH/ELK_OUT_F\);
    
    HIEFFPLA_INST_0_52752 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_21[3]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_22[3]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[0]\, Y => 
        HIEFFPLA_NET_0_117517);
    
    HIEFFPLA_INST_0_52636 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_13[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_14[1]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_2[0]\, Y => 
        HIEFFPLA_NET_0_117535);
    
    \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[12]\ : DFN1C0
      port map(D => 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]_net_1\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[12]_net_1\);
    
    \P_OP_MODE1_SPE_pad/U0/U1\ : IOTRI_OB_EB
      port map(D => \OP_MODE_c[1]\, E => \VCC\, DOUT => 
        \P_OP_MODE1_SPE_pad/U0/NET1\, EOUT => 
        \P_OP_MODE1_SPE_pad/U0/NET2\);
    
    HIEFFPLA_INST_0_45435 : NAND2A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_19[6]\, Y => 
        HIEFFPLA_NET_0_118915);
    
    HIEFFPLA_INST_0_41813 : AOI1
      port map(A => HIEFFPLA_NET_0_119389, B => 
        \U50_PATTERNS/SM_BANK_SEL[19]\, C => 
        HIEFFPLA_NET_0_119665, Y => HIEFFPLA_NET_0_119691);
    
    HIEFFPLA_INST_0_37435 : MX2
      port map(A => \U200A_TFC/LOC_STOP_ADDR[5]\, B => 
        \TFC_STOP_ADDR[5]\, S => \U200A_TFC/GP_PG_SM_0[10]_net_1\, 
        Y => HIEFFPLA_NET_0_120285);
    
    HIEFFPLA_INST_0_46487 : AND3B
      port map(A => HIEFFPLA_NET_0_119571, B => 
        \U50_PATTERNS/RD_USB_ADBUS[1]\, C => 
        HIEFFPLA_NET_0_119587, Y => HIEFFPLA_NET_0_118680);
    
    \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_115926, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_9, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[4]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_28[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116052, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_15, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_28[3]\);
    
    \U_ELK3_CH/U_ELK1_SERDAT_SOURCE/SERDAT[6]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118097, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_15, Q => 
        \U_ELK3_CH/ELK_TX_DAT[6]\);
    
    HIEFFPLA_INST_0_63002 : AND2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[0]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[1]\, Y => 
        HIEFFPLA_NET_0_115918);
    
    \U_ELK14_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]\ : DFN1C0
      port map(D => \U_ELK14_CH/U_SLAVE_1ELK/Q[8]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]_net_1\);
    
    HIEFFPLA_INST_0_44472 : MX2
      port map(A => \ELKS_STRT_ADDR[3]\, B => 
        \U50_PATTERNS/U4C_REGCROSS/SAMP_TWO[3]_net_1\, S => 
        HIEFFPLA_NET_0_119114, Y => HIEFFPLA_NET_0_119109);
    
    HIEFFPLA_INST_0_53608 : MX2
      port map(A => HIEFFPLA_NET_0_117291, B => 
        HIEFFPLA_NET_0_117419, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[2]_net_1\, Y
         => HIEFFPLA_NET_0_117383);
    
    \U_ELK13_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]\ : DFN1C0
      port map(D => \U_ELK13_CH/U_SLAVE_1ELK/Q[5]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]_net_1\);
    
    \U50_PATTERNS/ELINK_DINA_12[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119842, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_12, Q => 
        \U50_PATTERNS/ELINK_DINA_12[5]\);
    
    \U50_PATTERNS/ELINK_ADDRA_10[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120087, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_21, Q => 
        \U50_PATTERNS/ELINK_ADDRA_10[0]\);
    
    HIEFFPLA_INST_0_55191 : AND3B
      port map(A => HIEFFPLA_NET_0_116941, B => 
        HIEFFPLA_NET_0_116943, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[7]_net_1\, Y => 
        HIEFFPLA_NET_0_117099);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_26[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116403, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_21, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_26[3]\);
    
    \U_ELK0_CMD_TX/SER_CMD_WORD_F[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118666, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_17, Q => 
        \U_ELK0_CMD_TX/SER_CMD_WORD_F[3]_net_1\);
    
    HIEFFPLA_INST_0_53491 : MX2
      port map(A => HIEFFPLA_NET_0_117405, B => 
        HIEFFPLA_NET_0_117295, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[2]_net_1\, Y
         => HIEFFPLA_NET_0_117400);
    
    \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_1[4]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_115935, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_24_0, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_1[4]_net_1\);
    
    \U_ELK16_CH/U_SLAVE_1ELK/RECD_SER_WORD[0]\ : DFN1C0
      port map(D => \U_ELK16_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[0]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_16[0]\);
    
    \U50_PATTERNS/ELINK_DINA_19[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119784, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_1, Q => 
        \U50_PATTERNS/ELINK_DINA_19[7]\);
    
    HIEFFPLA_INST_0_52335 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_BIT_OS_VAL[1]\, B
         => HIEFFPLA_NET_0_117575, S => HIEFFPLA_NET_0_117111, Y
         => HIEFFPLA_NET_0_117579);
    
    HIEFFPLA_INST_0_48208 : MX2
      port map(A => \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\, 
        B => \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[13]_net_1\, S => 
        \BIT_OS_SEL_1[2]\, Y => HIEFFPLA_NET_0_118353);
    
    \U50_PATTERNS/REG_STATE_0[4]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119480, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_22_0, Q => 
        \U50_PATTERNS/REG_STATE_0[4]_net_1\);
    
    \U_ELK9_CH/U_SLAVE_1ELK/Q[8]\ : DFN1C0
      port map(D => \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/Q[8]_net_1\);
    
    HIEFFPLA_INST_0_56544 : AND3A
      port map(A => HIEFFPLA_NET_0_117430, B => \BIT_OS_SEL_1[2]\, 
        C => \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[12]_net_1\, 
        Y => HIEFFPLA_NET_0_116842);
    
    \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[4]\ : DFN1C0
      port map(D => 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\);
    
    HIEFFPLA_INST_0_53957 : MX2
      port map(A => HIEFFPLA_NET_0_116123, B => 
        HIEFFPLA_NET_0_116021, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[3]_net_1\, Y
         => HIEFFPLA_NET_0_117327);
    
    HIEFFPLA_INST_0_50150 : MX2
      port map(A => \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[2]_net_1\, B
         => \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\, S => 
        \BIT_OS_SEL_6[2]\, Y => HIEFFPLA_NET_0_118001);
    
    HIEFFPLA_INST_0_48897 : MX2
      port map(A => HIEFFPLA_NET_0_118217, B => 
        HIEFFPLA_NET_0_118229, S => \BIT_OS_SEL_0[1]\, Y => 
        HIEFFPLA_NET_0_118227);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_10[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116273, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_18, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_10[2]\);
    
    HIEFFPLA_INST_0_56634 : AXOI4
      port map(A => HIEFFPLA_NET_0_117085, B => 
        HIEFFPLA_NET_0_117602, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_0[0]\, Y => 
        HIEFFPLA_NET_0_116824);
    
    HIEFFPLA_INST_0_54055 : MX2
      port map(A => HIEFFPLA_NET_0_116462, B => 
        HIEFFPLA_NET_0_116382, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[3]_net_1\, Y
         => HIEFFPLA_NET_0_117314);
    
    HIEFFPLA_INST_0_49025 : MX2
      port map(A => HIEFFPLA_NET_0_118221, B => 
        HIEFFPLA_NET_0_118224, S => \BIT_OS_SEL_2[0]\, Y => 
        \U_ELK19_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[5]\);
    
    \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[10]\ : DFN1C0
      port map(D => 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]_net_1\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\);
    
    HIEFFPLA_INST_0_62941 : MX2
      port map(A => HIEFFPLA_NET_0_115890, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[4]\, S => 
        HIEFFPLA_NET_0_117073, Y => HIEFFPLA_NET_0_115926);
    
    HIEFFPLA_INST_0_45082 : MX2
      port map(A => HIEFFPLA_NET_0_118977, B => 
        \U50_PATTERNS/WR_USB_ADBUS[0]\, S => 
        HIEFFPLA_NET_0_119486, Y => HIEFFPLA_NET_0_118985);
    
    \U_ELK9_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]\ : DFN1C0
      port map(D => \U_ELK9_CH/U_SLAVE_1ELK/Q[9]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]_net_1\);
    
    HIEFFPLA_INST_0_57934 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_7[7]\, B => 
        HIEFFPLA_NET_0_116577, S => HIEFFPLA_NET_0_117113, Y => 
        HIEFFPLA_NET_0_116596);
    
    HIEFFPLA_INST_0_43564 : AND2A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/SM_BANK_SEL[2]\, Y => HIEFFPLA_NET_0_119290);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_4[5]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116691, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_9, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_4[5]\);
    
    \U_ELK5_CH/U_SLAVE_1ELK/Q[5]\ : DFN1C0
      port map(D => \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/Q[5]_net_1\);
    
    HIEFFPLA_INST_0_39488 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_3[6]\, B => 
        HIEFFPLA_NET_0_119517, S => HIEFFPLA_NET_0_119247, Y => 
        HIEFFPLA_NET_0_119985);
    
    \U_ELK13_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]\ : DFN1C0
      port map(D => \U_ELK13_CH/U_SLAVE_1ELK/Q[1]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]_net_1\);
    
    HIEFFPLA_INST_0_49274 : MX2
      port map(A => HIEFFPLA_NET_0_118176, B => 
        HIEFFPLA_NET_0_118170, S => \BIT_OS_SEL_2[0]\, Y => 
        \U_ELK1_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[5]\);
    
    HIEFFPLA_INST_0_55056 : AO1C
      port map(A => HIEFFPLA_NET_0_117211, B => 
        HIEFFPLA_NET_0_117083, C => HIEFFPLA_NET_0_117180, Y => 
        HIEFFPLA_NET_0_117132);
    
    HIEFFPLA_INST_0_42614 : AND2
      port map(A => \U50_PATTERNS/REG_ADDR[1]\, B => 
        \U50_PATTERNS/REG_ADDR[0]\, Y => HIEFFPLA_NET_0_119500);
    
    \U_ELK4_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118065, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_1, Q => 
        \U_ELK4_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]_net_1\);
    
    HIEFFPLA_INST_0_53616 : MX2
      port map(A => HIEFFPLA_NET_0_117342, B => 
        HIEFFPLA_NET_0_117420, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[1]_net_1\, Y
         => HIEFFPLA_NET_0_117382);
    
    HIEFFPLA_INST_0_47499 : MX2
      port map(A => HIEFFPLA_NET_0_118494, B => 
        HIEFFPLA_NET_0_118490, S => \BIT_OS_SEL_4[0]\, Y => 
        \U_ELK13_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[1]\);
    
    \U_ELK12_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]\ : DFN1C0
      port map(D => \U_ELK12_CH/U_SLAVE_1ELK/Q[4]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]_net_1\);
    
    \U_ELK16_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118379, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_14, Q => 
        \U_ELK16_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]_net_1\);
    
    \U_ELK13_CH/U_SLAVE_1ELK/RECD_SER_WORD[4]\ : DFN1C0
      port map(D => \U_ELK13_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[4]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_13[4]\);
    
    HIEFFPLA_INST_0_42338 : AND2A
      port map(A => HIEFFPLA_NET_0_119275, B => 
        \U50_PATTERNS/RD_USB_ADBUS[5]\, Y => 
        HIEFFPLA_NET_0_119567);
    
    HIEFFPLA_INST_0_61712 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_25[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_26[1]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_4[0]\, Y => 
        HIEFFPLA_NET_0_116089);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_29[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116376, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_4, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_29[2]\);
    
    \U_TFC_CMD_TX/SER_CMD_WORD_R[1]\ : DFN1C0
      port map(D => \U_TFC_CMD_TX/N_SER_CMD_WORD_R[1]\, CLK => 
        CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_TFC_CMD_TX/SER_CMD_WORD_R[1]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/PHASE_ADJ[1]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[1]_net_1\, CLK
         => CLK_40M_GL, CLR => P_MASTER_POR_B_c, Q => 
        \U_MASTER_DES/PHASE_ADJ_160_L[1]\);
    
    HIEFFPLA_INST_0_43440 : MX2
      port map(A => \U50_PATTERNS/SM_BANK_SEL[1]\, B => 
        HIEFFPLA_NET_0_119217, S => HIEFFPLA_NET_0_118691, Y => 
        HIEFFPLA_NET_0_119311);
    
    HIEFFPLA_INST_0_41887 : AOI1C
      port map(A => \U50_PATTERNS/ELINK_RWA[5]\, B => 
        HIEFFPLA_NET_0_119642, C => HIEFFPLA_NET_0_119673, Y => 
        HIEFFPLA_NET_0_119674);
    
    HIEFFPLA_INST_0_54700 : MX2
      port map(A => HIEFFPLA_NET_0_117285, B => 
        HIEFFPLA_NET_0_117277, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[2]_net_1\, Y => 
        HIEFFPLA_NET_0_117221);
    
    HIEFFPLA_INST_0_47258 : MX2
      port map(A => HIEFFPLA_NET_0_118538, B => 
        HIEFFPLA_NET_0_118534, S => \BIT_OS_SEL_5[0]\, Y => 
        \U_ELK12_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[2]\);
    
    HIEFFPLA_INST_0_47025 : MX2
      port map(A => HIEFFPLA_NET_0_118576, B => 
        HIEFFPLA_NET_0_118588, S => \BIT_OS_SEL[0]\, Y => 
        \U_ELK11_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[4]\);
    
    HIEFFPLA_INST_0_46744 : MX2
      port map(A => HIEFFPLA_NET_0_118611, B => 
        HIEFFPLA_NET_0_118632, S => \BIT_OS_SEL_0[0]\, Y => 
        \U_ELK10_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[0]\);
    
    HIEFFPLA_INST_0_42869 : AND2A
      port map(A => \U50_PATTERNS/REG_STATE[3]_net_1\, B => 
        \U50_PATTERNS/REG_STATE[2]_net_1\, Y => 
        HIEFFPLA_NET_0_119441);
    
    HIEFFPLA_INST_0_37843 : NAND3A
      port map(A => \U200B_ELINKS/GP_PG_SM[4]_net_1\, B => 
        \U200B_ELINKS/GP_PG_SM[5]_net_1\, C => 
        HIEFFPLA_NET_0_120222, Y => HIEFFPLA_NET_0_120193);
    
    HIEFFPLA_INST_0_59029 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_6[2]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_22[2]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_2[4]_net_1\, Y
         => HIEFFPLA_NET_0_116445);
    
    \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[41]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117711, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_33, Q => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[41]_net_1\);
    
    \U_ELK17_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]\ : DFN1C0
      port map(D => \U_ELK17_CH/U_SLAVE_1ELK/Q[8]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]_net_1\);
    
    \U50_PATTERNS/ELINK_DINA_6[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119742, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_16, Q => 
        \U50_PATTERNS/ELINK_DINA_6[1]\);
    
    HIEFFPLA_INST_0_51545 : AND3
      port map(A => 
        \U_EXEC_MASTER/USB_MASTER_EN/T_CNT60M[5]_net_1\, B => 
        \U_EXEC_MASTER/USB_MASTER_EN/T_CNT60M[4]_net_1\, C => 
        HIEFFPLA_NET_0_117747, Y => HIEFFPLA_NET_0_117748);
    
    HIEFFPLA_INST_0_51214 : MX2
      port map(A => \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\, B
         => \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[11]_net_1\, S => 
        \BIT_OS_SEL_2[2]\, Y => HIEFFPLA_NET_0_117811);
    
    HIEFFPLA_INST_0_53870 : NAND3C
      port map(A => HIEFFPLA_NET_0_117389, B => 
        HIEFFPLA_NET_0_117350, C => HIEFFPLA_NET_0_117071, Y => 
        HIEFFPLA_NET_0_117339);
    
    HIEFFPLA_INST_0_47152 : MX2
      port map(A => HIEFFPLA_NET_0_118541, B => 
        HIEFFPLA_NET_0_118537, S => \BIT_OS_SEL_4[1]\, Y => 
        HIEFFPLA_NET_0_118542);
    
    HIEFFPLA_INST_0_51104 : AND2
      port map(A => CLK_40M_GL, B => 
        \U_ELK9_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0_net_1\, Y => 
        HIEFFPLA_NET_0_117834);
    
    HIEFFPLA_INST_0_49258 : MX2
      port map(A => HIEFFPLA_NET_0_118183, B => 
        HIEFFPLA_NET_0_118177, S => \BIT_OS_SEL_2[0]\, Y => 
        \U_ELK1_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[3]\);
    
    \U50_PATTERNS/U4B_REGCROSS/SAMP_TWO[2]\ : DFN1C0
      port map(D => \U50_PATTERNS/U4B_REGCROSS/SAMP_ONE[2]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_29, Q => 
        \U50_PATTERNS/U4B_REGCROSS/SAMP_TWO[2]_net_1\);
    
    HIEFFPLA_INST_0_60675 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_14[1]\, B => 
        HIEFFPLA_NET_0_117167, S => HIEFFPLA_NET_0_117228, Y => 
        HIEFFPLA_NET_0_116234);
    
    HIEFFPLA_INST_0_56977 : XA1C
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_1[6]\, B => 
        HIEFFPLA_NET_0_116777, C => HIEFFPLA_NET_0_117179, Y => 
        HIEFFPLA_NET_0_116761);
    
    HIEFFPLA_INST_0_49148 : MX2
      port map(A => \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[1]_net_1\, B
         => \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\, S => 
        \BIT_OS_SEL[2]\, Y => HIEFFPLA_NET_0_118182);
    
    HIEFFPLA_INST_0_56127 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/MAX_CNT[7]\, 
        B => HIEFFPLA_NET_0_116932, S => HIEFFPLA_NET_0_117084, Y
         => HIEFFPLA_NET_0_116947);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_9[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_115964, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_20, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_9[1]\);
    
    HIEFFPLA_INST_0_43125 : AND3B
      port map(A => \U50_PATTERNS/REG_STATE[0]_net_1\, B => 
        \U50_PATTERNS/REG_STATE[3]_net_1\, C => 
        \U50_PATTERNS/REG_STATE[1]_net_1\, Y => 
        HIEFFPLA_NET_0_119367);
    
    \U_ELK8_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117881, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_15, Q => 
        \U_ELK8_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]_net_1\);
    
    \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[5]\ : DFN1C0
      port map(D => 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\);
    
    HIEFFPLA_INST_0_63198 : AND2
      port map(A => \TFC_TX_DAT[0]\, B => 
        \U_TFC_CMD_TX/START_RISE_net_1\, Y => 
        \U_TFC_CMD_TX/N_SER_CMD_WORD_F[0]\);
    
    HIEFFPLA_INST_0_44769 : NAND3C
      port map(A => HIEFFPLA_NET_0_119052, B => 
        HIEFFPLA_NET_0_119050, C => HIEFFPLA_NET_0_119053, Y => 
        HIEFFPLA_NET_0_119054);
    
    HIEFFPLA_INST_0_39110 : MX2
      port map(A => HIEFFPLA_NET_0_119519, B => 
        \U50_PATTERNS/ELINK_ADDRA_17[4]\, S => 
        HIEFFPLA_NET_0_119260, Y => HIEFFPLA_NET_0_120027);
    
    HIEFFPLA_INST_0_61499 : MX2
      port map(A => HIEFFPLA_NET_0_117181, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_23[2]\, S => 
        HIEFFPLA_NET_0_117151, Y => HIEFFPLA_NET_0_116118);
    
    HIEFFPLA_INST_0_46343 : AO1
      port map(A => HIEFFPLA_NET_0_119277, B => 
        \U50_PATTERNS/ELINK_DOUTA_11[2]\, C => 
        HIEFFPLA_NET_0_118851, Y => HIEFFPLA_NET_0_118712);
    
    HIEFFPLA_INST_0_45716 : AO1
      port map(A => HIEFFPLA_NET_0_119288, B => 
        \U50_PATTERNS/ELINK_DOUTA_16[1]\, C => 
        HIEFFPLA_NET_0_118786, Y => HIEFFPLA_NET_0_118859);
    
    HIEFFPLA_INST_0_41179 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_3[1]\, B => 
        HIEFFPLA_NET_0_119576, S => HIEFFPLA_NET_0_119247, Y => 
        HIEFFPLA_NET_0_119766);
    
    \U50_PATTERNS/U4E_REGCROSS/LOCAL_REG_VAL_5[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119057, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_1, Q => \OP_MODE_c_5[1]\);
    
    \U_ELK13_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118510, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_16, Q => 
        \U_ELK13_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]_net_1\);
    
    HIEFFPLA_INST_0_57379 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_4[4]\, B => 
        HIEFFPLA_NET_0_116667, S => HIEFFPLA_NET_0_117122, Y => 
        HIEFFPLA_NET_0_116692);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_16[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116213, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_5, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_16[2]\);
    
    \U200B_ELINKS/ADDR_POINTER[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120255, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_31_0, Q => \ELKS_ADDRB[0]\);
    
    HIEFFPLA_INST_0_39200 : MX2
      port map(A => HIEFFPLA_NET_0_119517, B => 
        \U50_PATTERNS/ELINK_ADDRA_18[6]\, S => 
        HIEFFPLA_NET_0_119264, Y => HIEFFPLA_NET_0_120017);
    
    HIEFFPLA_INST_0_54014 : MX2
      port map(A => HIEFFPLA_NET_0_117422, B => 
        HIEFFPLA_NET_0_117255, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[1]_net_1\, Y
         => HIEFFPLA_NET_0_117320);
    
    HIEFFPLA_INST_0_50364 : AND2A
      port map(A => \OP_MODE_c_1[1]\, B => \PATT_ELK_DAT_6[6]\, Y
         => HIEFFPLA_NET_0_117962);
    
    HIEFFPLA_INST_0_38678 : MX2
      port map(A => HIEFFPLA_NET_0_119519, B => 
        \U50_PATTERNS/ELINK_ADDRA_11[4]\, S => 
        HIEFFPLA_NET_0_119280, Y => HIEFFPLA_NET_0_120075);
    
    \U_ELK14_CH/U_SLAVE_1ELK/Q[10]\ : DFN1C0
      port map(D => \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/Q[10]_net_1\);
    
    HIEFFPLA_INST_0_51861 : NAND2B
      port map(A => HIEFFPLA_NET_0_117629, B => 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM_0[4]_net_1\, Y => 
        HIEFFPLA_NET_0_117674);
    
    \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[10]\ : DFN1C0
      port map(D => 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\);
    
    \U_ELK15_CH/U_SLAVE_1ELK/RECD_SER_WORD[6]\ : DFN1C0
      port map(D => \U_ELK15_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[6]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_15[6]\);
    
    HIEFFPLA_INST_0_63139 : AX1C
      port map(A => HIEFFPLA_NET_0_115875, B => 
        HIEFFPLA_NET_0_115876, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[4]_net_1\, Y => 
        HIEFFPLA_NET_0_115878);
    
    HIEFFPLA_INST_0_50453 : MX2
      port map(A => \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\, B
         => \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[11]_net_1\, S => 
        \BIT_OS_SEL_5[2]\, Y => HIEFFPLA_NET_0_117948);
    
    \U_ELK2_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]\ : DFN1C0
      port map(D => \U_ELK2_CH/U_SLAVE_1ELK/Q[3]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]_net_1\);
    
    HIEFFPLA_INST_0_42351 : AND2A
      port map(A => HIEFFPLA_NET_0_119275, B => 
        \U50_PATTERNS/RD_USB_ADBUS[7]\, Y => 
        HIEFFPLA_NET_0_119560);
    
    HIEFFPLA_INST_0_58899 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_4[2]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_20[2]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_2[4]_net_1\, Y
         => HIEFFPLA_NET_0_116461);
    
    HIEFFPLA_INST_0_42948 : AO1
      port map(A => HIEFFPLA_NET_0_119367, B => 
        HIEFFPLA_NET_0_119569, C => HIEFFPLA_NET_0_119396, Y => 
        HIEFFPLA_NET_0_119417);
    
    HIEFFPLA_INST_0_42326 : AND2A
      port map(A => HIEFFPLA_NET_0_119275, B => 
        \U50_PATTERNS/RD_USB_ADBUS[4]\, Y => 
        HIEFFPLA_NET_0_119570);
    
    HIEFFPLA_INST_0_61007 : MX2
      port map(A => HIEFFPLA_NET_0_117166, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_18[4]\, S => 
        HIEFFPLA_NET_0_117134, Y => HIEFFPLA_NET_0_116186);
    
    HIEFFPLA_INST_0_60162 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_7[1]\, B => 
        HIEFFPLA_NET_0_116677, S => HIEFFPLA_NET_0_117157, Y => 
        HIEFFPLA_NET_0_116302);
    
    \U_ELK4_CH/U_SLAVE_1ELK/RECD_SER_WORD[4]\ : DFN1C0
      port map(D => \U_ELK4_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[4]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_4[4]\);
    
    \U50_PATTERNS/ELINK_DINA_11[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119854, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_11, Q => 
        \U50_PATTERNS/ELINK_DINA_11[1]\);
    
    \U_ELK16_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL\ : DFN1C0
      port map(D => \U_ELK16_CH/ELK_IN_F_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL_net_1\);
    
    \U_ELK10_CH/U_SLAVE_1ELK/Q[5]\ : DFN1C0
      port map(D => \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/Q[5]_net_1\);
    
    HIEFFPLA_INST_0_41647 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_9[5]\, B => 
        HIEFFPLA_NET_0_119567, S => HIEFFPLA_NET_0_119292, Y => 
        HIEFFPLA_NET_0_119714);
    
    HIEFFPLA_INST_0_111810 : OR3B
      port map(A => HIEFFPLA_NET_0_117629, B => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[1]\, C => 
        HIEFFPLA_NET_0_117682, Y => HIEFFPLA_NET_0_115830);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_16[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116510, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_16_0, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_16[2]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_3[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116725, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_7, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_3[0]\);
    
    HIEFFPLA_INST_0_51551 : AND3
      port map(A => 
        \U_EXEC_MASTER/USB_MASTER_EN/T_CNT60M[0]_net_1\, B => 
        \U_EXEC_MASTER/USB_MASTER_EN/T_CNT60M[1]_net_1\, C => 
        \U_EXEC_MASTER/USB_MASTER_EN/T_CNT60M[2]_net_1\, Y => 
        HIEFFPLA_NET_0_117746);
    
    \U_ELK17_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]\ : DFN1C0
      port map(D => \U_ELK17_CH/U_SLAVE_1ELK/Q[10]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]_net_1\);
    
    \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[8]\ : DFN1C0
      port map(D => 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\);
    
    HIEFFPLA_INST_0_45820 : NAND2A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_12[5]\, Y => 
        HIEFFPLA_NET_0_118832);
    
    HIEFFPLA_INST_0_56616 : AND3
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[12]_net_1\, B
         => HIEFFPLA_NET_0_117424, C => HIEFFPLA_NET_0_117427, Y
         => HIEFFPLA_NET_0_116827);
    
    HIEFFPLA_INST_0_37417 : MX2
      port map(A => \U200A_TFC/LOC_STOP_ADDR[2]\, B => 
        \TFC_STOP_ADDR[2]\, S => \U200A_TFC/GP_PG_SM_0[10]_net_1\, 
        Y => HIEFFPLA_NET_0_120288);
    
    AFLSDF_INV_4 : INV
      port map(A => P_USB_MASTER_EN_c_22, Y => \AFLSDF_INV_4\);
    
    \U_ELK17_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118331, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_14, Q => 
        \U_ELK17_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]_net_1\);
    
    \U50_PATTERNS/U4C_REGCROSS/SAMP_TWO[5]\ : DFN1C0
      port map(D => \U50_PATTERNS/U4C_REGCROSS/SAMP_ONE[5]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_22_0, Q => 
        \U50_PATTERNS/U4C_REGCROSS/SAMP_TWO[5]_net_1\);
    
    HIEFFPLA_INST_0_46086 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/SM_BANK_SEL[13]\, C => 
        \U50_PATTERNS/ELINK_DOUTA_6[6]\, Y => 
        HIEFFPLA_NET_0_118770);
    
    HIEFFPLA_INST_0_59005 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_22[2]\, B => 
        HIEFFPLA_NET_0_116687, S => HIEFFPLA_NET_0_117095, Y => 
        HIEFFPLA_NET_0_116448);
    
    HIEFFPLA_INST_0_52276 : AND2B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[5]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[4]_net_1\, Y => 
        HIEFFPLA_NET_0_117593);
    
    HIEFFPLA_INST_0_48619 : AND2A
      port map(A => \OP_MODE_c_2[1]\, B => \PATT_ELK_DAT_18[4]\, 
        Y => HIEFFPLA_NET_0_118279);
    
    HIEFFPLA_INST_0_43777 : AND3A
      port map(A => HIEFFPLA_NET_0_119585, B => 
        HIEFFPLA_NET_0_119563, C => HIEFFPLA_NET_0_119597, Y => 
        HIEFFPLA_NET_0_119216);
    
    \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_SEL_4[2]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_BIT_OS_VAL[2]\, CLK
         => CLK_40M_GL, CLR => P_MASTER_POR_B_c_27_0, Q => 
        \BIT_OS_SEL_4[2]\);
    
    HIEFFPLA_INST_0_61475 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_6[0]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_22[0]\, S
         => \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_5[4]_net_1\, 
        Y => HIEFFPLA_NET_0_116121);
    
    HIEFFPLA_INST_0_60232 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_8[0]\, B => 
        HIEFFPLA_NET_0_116680, S => HIEFFPLA_NET_0_117160, Y => 
        HIEFFPLA_NET_0_116293);
    
    HIEFFPLA_INST_0_51070 : MX2
      port map(A => 
        \U_ELK9_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]_net_1\, B => 
        \U_ELK9_CH/ELK_TX_DAT[2]\, S => 
        \U_ELK9_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_117841);
    
    HIEFFPLA_INST_0_62475 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_6[1]\, 
        B => HIEFFPLA_NET_0_117114, S => HIEFFPLA_NET_0_117132, Y
         => HIEFFPLA_NET_0_115984);
    
    HIEFFPLA_INST_0_43844 : MX2
      port map(A => HIEFFPLA_NET_0_119520, B => 
        \U50_PATTERNS/TFC_ADDRA[3]\, S => HIEFFPLA_NET_0_119294, 
        Y => HIEFFPLA_NET_0_119204);
    
    \U50_PATTERNS/ELINK_DINA_10[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119858, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_9, Q => 
        \U50_PATTERNS/ELINK_DINA_10[5]\);
    
    HIEFFPLA_INST_0_61277 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_4[1]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_20[1]\, S
         => \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_5[4]_net_1\, 
        Y => HIEFFPLA_NET_0_116149);
    
    HIEFFPLA_INST_0_56315 : AO1
      port map(A => HIEFFPLA_NET_0_117429, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[2]_net_1\, C => 
        HIEFFPLA_NET_0_116871, Y => HIEFFPLA_NET_0_116895);
    
    \U50_PATTERNS/ELINK_ADDRA_3[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119990, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_1, Q => 
        \U50_PATTERNS/ELINK_ADDRA_3[1]\);
    
    HIEFFPLA_INST_0_46578 : NAND2B
      port map(A => \OP_MODE_c_4[1]\, B => \PATT_ELK_DAT_0[2]\, Y
         => HIEFFPLA_NET_0_118658);
    
    HIEFFPLA_INST_0_45382 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/SM_BANK_SEL[2]\, C => 
        \U50_PATTERNS/ELINK_DOUTA_17[5]\, Y => 
        HIEFFPLA_NET_0_118925);
    
    \U50_PATTERNS/ELINK_RWA[10]/U1\ : DFN1P0
      port map(D => HIEFFPLA_NET_0_119710, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_11, Q => 
        \U50_PATTERNS/ELINK_RWA[10]\);
    
    HIEFFPLA_INST_0_41965 : AND3C
      port map(A => HIEFFPLA_NET_0_119255, B => 
        HIEFFPLA_NET_0_119262, C => 
        \U50_PATTERNS/SM_BANK_SEL[16]\, Y => 
        HIEFFPLA_NET_0_119643);
    
    \U50_PATTERNS/ELINK_ADDRA_0[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120094, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_18, Q => 
        \U50_PATTERNS/ELINK_ADDRA_0[1]\);
    
    HIEFFPLA_INST_0_62658 : MX2
      port map(A => HIEFFPLA_NET_0_117075, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_9[3]\, S => 
        HIEFFPLA_NET_0_117183, Y => HIEFFPLA_NET_0_115962);
    
    HIEFFPLA_INST_0_53142 : MX2
      port map(A => HIEFFPLA_NET_0_117540, B => 
        HIEFFPLA_NET_0_117536, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_1[3]\, Y => 
        HIEFFPLA_NET_0_117460);
    
    \EXT_INT_REF_SEL_pad/U0/U1\ : IOIN_IB
      port map(YIN => \EXT_INT_REF_SEL_pad/U0/NET1\, Y => 
        EXT_INT_REF_SEL_c);
    
    HIEFFPLA_INST_0_38068 : NAND3B
      port map(A => \U200B_ELINKS/RX_SER_WORD_2DEL[6]_net_1\, B
         => \U200B_ELINKS/RX_SER_WORD_2DEL[4]_net_1\, C => 
        \U200B_ELINKS/RX_SER_WORD_2DEL[7]_net_1\, Y => 
        HIEFFPLA_NET_0_120161);
    
    HIEFFPLA_INST_0_63116 : AND2A
      port map(A => HIEFFPLA_NET_0_115916, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[9]\, Y => 
        HIEFFPLA_NET_0_115884);
    
    HIEFFPLA_INST_0_59465 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_27[3]\, B => 
        HIEFFPLA_NET_0_116815, S => HIEFFPLA_NET_0_117162, Y => 
        HIEFFPLA_NET_0_116391);
    
    HIEFFPLA_INST_0_49477 : MX2
      port map(A => \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[1]_net_1\, B
         => \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\, S => 
        \BIT_OS_SEL_7[2]\, Y => HIEFFPLA_NET_0_118125);
    
    HIEFFPLA_INST_0_41386 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_6[0]\, B => 
        HIEFFPLA_NET_0_119578, S => HIEFFPLA_NET_0_119258, Y => 
        HIEFFPLA_NET_0_119743);
    
    \U_ELK5_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2\ : IOPADN_BI
      port map(DB => \U_ELK5_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, 
        E => \U_ELK5_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET3\, PAD => 
        ELK5_DAT_N, N2POUT => 
        \U_ELK5_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2_N2P\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_6[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_115983, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_16, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_6[2]\);
    
    \U_ELK12_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0\ : DFN1C0
      port map(D => CLK_40M_GL, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_6, Q => 
        \U_ELK12_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0_net_1\);
    
    \U50_PATTERNS/REG_ADDR[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119527, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_10, Q => \U50_PATTERNS/REG_ADDR[6]\);
    
    HIEFFPLA_INST_0_46547 : MX2
      port map(A => HIEFFPLA_NET_0_161280, B => 
        HIEFFPLA_NET_0_161279, S => HIEFFPLA_NET_0_161278, Y => 
        HIEFFPLA_NET_0_118667);
    
    HIEFFPLA_INST_0_43679 : AND2A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/SM_BANK_SEL[17]\, Y => 
        HIEFFPLA_NET_0_119244);
    
    \U_ELK10_CH/U_ELK1_SERDAT_SOURCE/SERDAT[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118642, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_17, Q => 
        \U_ELK10_CH/ELK_TX_DAT[1]\);
    
    HIEFFPLA_INST_0_48835 : MX2
      port map(A => 
        \U_ELK19_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]_net_1\, B => 
        \U_ELK19_CH/ELK_TX_DAT[4]\, S => 
        \U_ELK19_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118245);
    
    HIEFFPLA_INST_0_42802 : AND3C
      port map(A => \U50_PATTERNS/REG_STATE[1]_net_1\, B => 
        HIEFFPLA_NET_0_119432, C => HIEFFPLA_NET_0_118996, Y => 
        HIEFFPLA_NET_0_119460);
    
    \U_ELK19_CH/ELK_IN_F\ : DFN1C0
      port map(D => \U_ELK19_CH/ELK_IN_DDR_F\, CLK => 
        CCC_160M_ADJ, CLR => DEV_RST_B_c, Q => 
        \U_ELK19_CH/ELK_IN_F_net_1\);
    
    \U_ELK7_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0\ : DFN1C0
      port map(D => CLK_40M_GL, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_11, Q => 
        \U_ELK7_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0_net_1\);
    
    \U_ELK11_CH/ELK_IN_F\ : DFN1C0
      port map(D => \U_ELK11_CH/ELK_IN_DDR_F\, CLK => 
        CCC_160M_ADJ, CLR => DEV_RST_B_c, Q => 
        \U_ELK11_CH/ELK_IN_F_net_1\);
    
    HIEFFPLA_INST_0_50736 : MX2
      port map(A => HIEFFPLA_NET_0_117900, B => 
        HIEFFPLA_NET_0_117914, S => \BIT_OS_SEL_5[0]\, Y => 
        \U_ELK7_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[1]\);
    
    \U_ELK5_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U3\ : IOBI_ID_OD_EB
      port map(DR => \U_ELK5_CH/ELK_OUT_R\, DF => 
        \U_ELK5_CH/ELK_OUT_F\, CLR => \GND\, E => \AFLSDF_INV_43\, 
        ICLK => CCC_160M_ADJ, OCLK => CCC_160M_FXD, YIN => 
        \U_ELK5_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\, DOUT => OPEN, 
        EOUT => \U_ELK5_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET3\, YR
         => OPEN, YF => OPEN);
    
    \U_ELK7_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]\ : DFN1C0
      port map(D => \U_ELK7_CH/U_SLAVE_1ELK/Q[11]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]_net_1\);
    
    \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[2]\ : DFN1C0
      port map(D => \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\);
    
    HIEFFPLA_INST_0_49716 : MX2
      port map(A => HIEFFPLA_NET_0_118094, B => 
        HIEFFPLA_NET_0_118091, S => \BIT_OS_SEL_6[1]\, Y => 
        HIEFFPLA_NET_0_118081);
    
    \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[2]\ : DFN1C0
      port map(D => \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\);
    
    HIEFFPLA_INST_0_41269 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_4[3]\, B => 
        HIEFFPLA_NET_0_119574, S => HIEFFPLA_NET_0_119284, Y => 
        HIEFFPLA_NET_0_119756);
    
    HIEFFPLA_INST_0_37589 : AOI1A
      port map(A => HIEFFPLA_NET_0_120245, B => 
        HIEFFPLA_NET_0_120220, C => HIEFFPLA_NET_0_120252, Y => 
        HIEFFPLA_NET_0_120253);
    
    \U_ELK18_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]\ : DFN1C0
      port map(D => \U_ELK18_CH/U_SLAVE_1ELK/Q[8]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]_net_1\);
    
    HIEFFPLA_INST_0_47401 : MX2
      port map(A => \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\, 
        B => \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\, S => 
        \BIT_OS_SEL_3[2]\, Y => HIEFFPLA_NET_0_118497);
    
    \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_SEL_1[0]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_BIT_OS_VAL[0]\, CLK
         => CLK_40M_GL, CLR => P_MASTER_POR_B_c_27_0, Q => 
        \BIT_OS_SEL_1[0]\);
    
    \U50_PATTERNS/U4A_REGCROSS/LOCAL_REG_VAL[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119150, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_17, Q => \TFC_STRT_ADDR[4]\);
    
    HIEFFPLA_INST_0_43159 : AOI1A
      port map(A => \U50_PATTERNS/REG_STATE_0[5]_net_1\, B => 
        \U50_PATTERNS/REG_STATE[3]_net_1\, C => 
        \U50_PATTERNS/REG_STATE_0[2]_net_1\, Y => 
        HIEFFPLA_NET_0_119358);
    
    \U_REFCLKBUF/\\\\BIBUF_LVDS[0]\\\\/U0/U0\ : IOPADP_BI
      port map(N2PIN => 
        \U_REFCLKBUF/\\\\BIBUF_LVDS[0]\\\\/U0/U2_N2P\, D => 
        \U_REFCLKBUF/\\\\BIBUF_LVDS[0]\\\\/U0/NET1\, E => 
        \U_REFCLKBUF/\\\\BIBUF_LVDS[0]\\\\/U0/NET2\, PAD => 
        REF_CLK_0P, Y => 
        \U_REFCLKBUF/\\\\BIBUF_LVDS[0]\\\\/U0/NET4\);
    
    \U_ELK4_CH/U_SLAVE_1ELK/Q[1]\ : DFN1C0
      port map(D => \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/Q[1]_net_1\);
    
    HIEFFPLA_INST_0_62164 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_30[2]\, B => 
        HIEFFPLA_NET_0_117181, S => HIEFFPLA_NET_0_117330, Y => 
        HIEFFPLA_NET_0_116028);
    
    HIEFFPLA_INST_0_49109 : MX2
      port map(A => 
        \U_ELK1_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]_net_1\, B => 
        \U_ELK1_CH/ELK_TX_DAT[7]\, S => 
        \U_ELK1_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118195);
    
    HIEFFPLA_INST_0_46231 : AO1
      port map(A => HIEFFPLA_NET_0_119263, B => 
        \U50_PATTERNS/ELINK_DOUTA_8[6]\, C => 
        HIEFFPLA_NET_0_118735, Y => HIEFFPLA_NET_0_118736);
    
    HIEFFPLA_INST_0_46145 : AO1
      port map(A => HIEFFPLA_NET_0_119290, B => 
        \U50_PATTERNS/ELINK_DOUTA_17[6]\, C => 
        HIEFFPLA_NET_0_118931, Y => HIEFFPLA_NET_0_118756);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_20[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116467, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_13, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_20[0]\);
    
    \U_ELK18_CH/U_ELK1_SERDAT_SOURCE/SERDAT[5]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118278, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_13, Q => 
        \U_ELK18_CH/ELK_TX_DAT[5]\);
    
    HIEFFPLA_INST_0_47867 : AND2
      port map(A => CLK_40M_GL, B => 
        \U_ELK15_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0_net_1\, Y => 
        HIEFFPLA_NET_0_118419);
    
    HIEFFPLA_INST_0_52304 : AND3B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[0]_net_1\, B => 
        HIEFFPLA_NET_0_117585, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[4]_net_1\, Y => 
        HIEFFPLA_NET_0_117586);
    
    HIEFFPLA_INST_0_115780 : NAND2A
      port map(A => \TFC_ADDRB[0]\, B => 
        \U200A_TFC/LOC_STOP_ADDR[0]\, Y => HIEFFPLA_NET_0_115805);
    
    \U50_PATTERNS/ELINK_DINA_0[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119869, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_5, Q => 
        \U50_PATTERNS/ELINK_DINA_0[2]\);
    
    HIEFFPLA_INST_0_49387 : MX2
      port map(A => \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[2]_net_1\, B
         => \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\, S => 
        \BIT_OS_SEL_7[2]\, Y => HIEFFPLA_NET_0_118138);
    
    HIEFFPLA_INST_0_61775 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_26[1]\, B => 
        HIEFFPLA_NET_0_117114, S => HIEFFPLA_NET_0_117138, Y => 
        HIEFFPLA_NET_0_116079);
    
    \U_MASTER_DES/U13A_ADJ_160M/BITCNT[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117692, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_14, Q => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[6]\);
    
    \U_ELK1_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]\ : DFN1C0
      port map(D => \U_ELK1_CH/U_SLAVE_1ELK/Q[12]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]_net_1\);
    
    HIEFFPLA_INST_0_52446 : MX2
      port map(A => HIEFFPLA_NET_0_117514, B => 
        HIEFFPLA_NET_0_117510, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[3]\, Y => 
        HIEFFPLA_NET_0_117562);
    
    HIEFFPLA_INST_0_46883 : MX2
      port map(A => \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[3]_net_1\, 
        B => \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\, S => 
        \BIT_OS_SEL_4[2]\, Y => HIEFFPLA_NET_0_118590);
    
    HIEFFPLA_INST_0_50572 : MX2
      port map(A => 
        \U_ELK7_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]_net_1\, B => 
        \U_ELK7_CH/ELK_TX_DAT[2]\, S => 
        \U_ELK7_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_117931);
    
    HIEFFPLA_INST_0_49569 : MX2
      port map(A => \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\, 
        B => \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[14]_net_1\, S => 
        \BIT_OS_SEL_0[2]\, Y => HIEFFPLA_NET_0_118113);
    
    HIEFFPLA_INST_0_161260 : DFN1C0
      port map(D => DCB_SALT_SEL_c, CLK => CCC_160M_ADJ, CLR => 
        P_MASTER_POR_B_c_26, Q => HIEFFPLA_NET_0_161295);
    
    HIEFFPLA_INST_0_60310 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_9[2]\, B => 
        HIEFFPLA_NET_0_116277, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_0[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116283);
    
    HIEFFPLA_INST_0_56502 : AO1
      port map(A => HIEFFPLA_NET_0_117428, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[10]_net_1\, C
         => HIEFFPLA_NET_0_116834, Y => HIEFFPLA_NET_0_116850);
    
    \U_EXEC_MASTER/MPOR_B_26\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117787, CLK => CLK_40M_GL, CLR
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_0\, Q => 
        P_MASTER_POR_B_c_26);
    
    HIEFFPLA_INST_0_48356 : MX2
      port map(A => 
        \U_ELK17_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]_net_1\, B => 
        \U_ELK17_CH/ELK_TX_DAT[5]\, S => 
        \U_ELK17_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118331);
    
    \U_ELK9_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117837, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_0, Q => 
        \U_ELK9_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]_net_1\);
    
    \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[14]\ : DFN1C0
      port map(D => 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[14]_net_1\);
    
    HIEFFPLA_INST_0_49124 : MX2
      port map(A => HIEFFPLA_NET_0_118181, B => 
        HIEFFPLA_NET_0_118179, S => \BIT_OS_SEL_0[1]\, Y => 
        HIEFFPLA_NET_0_118185);
    
    \U_ELK9_CH/ELK_IN_F\ : DFN1C0
      port map(D => \U_ELK9_CH/ELK_IN_DDR_F\, CLK => CCC_160M_ADJ, 
        CLR => DEV_RST_B_c, Q => \U_ELK9_CH/ELK_IN_F_net_1\);
    
    HIEFFPLA_INST_0_38474 : MX2
      port map(A => \U50_PATTERNS/ELINKS_STRT_ADDR_T[5]\, B => 
        \U50_PATTERNS/RD_USB_ADBUS[5]\, S => 
        HIEFFPLA_NET_0_119493, Y => HIEFFPLA_NET_0_120098);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_27[4]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116066, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_13, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_27[4]\);
    
    \U_ELK18_CH/U_SLAVE_1ELK/Q[0]\ : DFN1C0
      port map(D => \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/Q[0]_net_1\);
    
    HIEFFPLA_INST_0_60042 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_5[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_21[1]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_5[4]_net_1\, Y
         => HIEFFPLA_NET_0_116318);
    
    HIEFFPLA_INST_0_52271 : NOR3B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[7]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[3]_net_1\, C => 
        HIEFFPLA_NET_0_117595, Y => HIEFFPLA_NET_0_117596);
    
    \U_MASTER_DES/U13C_MASTER_DESER/TUNE_CLKPHASE[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_115945, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_13, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/TUNE_CLKPHASE[4]\);
    
    HIEFFPLA_INST_0_40738 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_16[0]\, B => 
        HIEFFPLA_NET_0_119578, S => HIEFFPLA_NET_0_119257, Y => 
        HIEFFPLA_NET_0_119815);
    
    HIEFFPLA_INST_0_50648 : MX2
      port map(A => HIEFFPLA_NET_0_117909, B => 
        HIEFFPLA_NET_0_117907, S => \BIT_OS_SEL_4[1]\, Y => 
        HIEFFPLA_NET_0_117911);
    
    HIEFFPLA_INST_0_53515 : NAND2
      port map(A => HIEFFPLA_NET_0_117337, B => 
        HIEFFPLA_NET_0_116593, Y => HIEFFPLA_NET_0_117397);
    
    HIEFFPLA_INST_0_52966 : MX2
      port map(A => HIEFFPLA_NET_0_117470, B => 
        HIEFFPLA_NET_0_117466, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[4]\, Y => 
        HIEFFPLA_NET_0_117482);
    
    \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[2]\ : DFN1C0
      port map(D => \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\);
    
    HIEFFPLA_INST_0_37994 : MX2
      port map(A => \U200B_ELINKS/LOC_STRT_ADDR[2]\, B => 
        \ELKS_STRT_ADDR[2]\, S => 
        \U200B_ELINKS/GP_PG_SM_0[10]_net_1\, Y => 
        HIEFFPLA_NET_0_120177);
    
    \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[10]\ : DFN1C0
      port map(D => \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\);
    
    HIEFFPLA_INST_0_49945 : MX2
      port map(A => \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\, B
         => \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[12]_net_1\, S => 
        \BIT_OS_SEL_6[2]\, Y => HIEFFPLA_NET_0_118039);
    
    HIEFFPLA_INST_0_47140 : MX2
      port map(A => \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[3]_net_1\, 
        B => \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\, S => 
        \BIT_OS_SEL_3[2]\, Y => HIEFFPLA_NET_0_118544);
    
    HIEFFPLA_INST_0_111820 : MX2B
      port map(A => 
        \U_EXEC_MASTER/USB_MASTER_EN/CNT_EN_60M2S_net_1\, B => 
        HIEFFPLA_NET_0_115829, S => HIEFFPLA_NET_0_117753, Y => 
        HIEFFPLA_NET_0_117736);
    
    \U50_PATTERNS/ELINK_DINA_13[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119833, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_14, Q => 
        \U50_PATTERNS/ELINK_DINA_13[6]\);
    
    HIEFFPLA_INST_0_52402 : MX2
      port map(A => HIEFFPLA_NET_0_117520, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_29[0]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[3]\, Y => 
        HIEFFPLA_NET_0_117568);
    
    HIEFFPLA_INST_0_60140 : AND2
      port map(A => HIEFFPLA_NET_0_117211, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_6[0]\, Y => 
        HIEFFPLA_NET_0_116305);
    
    HIEFFPLA_INST_0_59540 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_12[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_28[1]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[4]_net_1\, Y
         => HIEFFPLA_NET_0_116381);
    
    HIEFFPLA_INST_0_40128 : AO1A
      port map(A => HIEFFPLA_NET_0_119874, B => 
        \U50_PATTERNS/ELINK_BLKA[19]\, C => HIEFFPLA_NET_0_119897, 
        Y => HIEFFPLA_NET_0_119898);
    
    \U_ELK14_CH/U_SLAVE_1ELK/RECD_SER_WORD[3]\ : DFN1C0
      port map(D => \U_ELK14_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[3]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_14[3]\);
    
    \U_ELK6_CH/U_SLAVE_1ELK/Q[13]\ : DFN1C0
      port map(D => \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[13]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/Q[13]_net_1\);
    
    \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[14]\ : DFN1C0
      port map(D => 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]_net_1\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[14]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_22[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116128, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_5, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_22[2]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/BEST_SEQCNT[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117438, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_9, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_SEQCNT[4]\);
    
    HIEFFPLA_INST_0_47124 : NAND2B
      port map(A => \OP_MODE_c_3[1]\, B => \PATT_ELK_DAT_12[3]\, 
        Y => HIEFFPLA_NET_0_118550);
    
    \U_ELK12_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]\ : DFN1C0
      port map(D => \U_ELK12_CH/U_SLAVE_1ELK/Q[2]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]_net_1\);
    
    HIEFFPLA_INST_0_58115 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_10[0]\, B => 
        HIEFFPLA_NET_0_116680, S => HIEFFPLA_NET_0_117165, Y => 
        HIEFFPLA_NET_0_116562);
    
    HIEFFPLA_INST_0_61631 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_8[0]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_24[0]\, S
         => \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_4[4]_net_1\, 
        Y => HIEFFPLA_NET_0_116100);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_30[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116028, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_7, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_30[2]\);
    
    \U50_PATTERNS/WR_USB_ADBUS[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118982, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_15, Q => 
        \U50_PATTERNS/WR_USB_ADBUS[3]\);
    
    \U50_PATTERNS/ELINK_DINA_12[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119843, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_12, Q => 
        \U50_PATTERNS/ELINK_DINA_12[4]\);
    
    HIEFFPLA_INST_0_51707 : NAND2B
      port map(A => 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM[4]_net_1\, B => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[11]_net_1\, Y => 
        HIEFFPLA_NET_0_117719);
    
    HIEFFPLA_INST_0_57017 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_2[1]\, B => 
        HIEFFPLA_NET_0_116734, S => HIEFFPLA_NET_0_117601, Y => 
        HIEFFPLA_NET_0_116754);
    
    HIEFFPLA_INST_0_52878 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_27[0]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_28[0]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_1[0]\, Y => 
        HIEFFPLA_NET_0_117496);
    
    AFLSDF_INV_24 : INV
      port map(A => DCB_SALT_SEL_c, Y => \AFLSDF_INV_24\);
    
    HIEFFPLA_INST_0_49965 : MX2
      port map(A => HIEFFPLA_NET_0_118041, B => 
        HIEFFPLA_NET_0_118039, S => \BIT_OS_SEL_6[1]\, Y => 
        HIEFFPLA_NET_0_118036);
    
    \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[6]\ : DFN1C0
      port map(D => 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\);
    
    HIEFFPLA_INST_0_49821 : AND2
      port map(A => \U_ELK4_CH/ELK_TX_DAT[0]\, B => 
        \U_ELK4_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118067);
    
    \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[8]\ : DFN1C0
      port map(D => \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\);
    
    \U50_PATTERNS/USB_TRIEN_B/U1\ : DFI1P0
      port map(D => HIEFFPLA_NET_0_119012, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_16, QN => \U50_PATTERNS/TrienAux\);
    
    HIEFFPLA_INST_0_58907 : MX2
      port map(A => HIEFFPLA_NET_0_116677, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_20[1]\, S => 
        HIEFFPLA_NET_0_117203, Y => HIEFFPLA_NET_0_116459);
    
    HIEFFPLA_INST_0_46503 : AOI1
      port map(A => HIEFFPLA_NET_0_119583, B => 
        HIEFFPLA_NET_0_119596, C => HIEFFPLA_NET_0_119571, Y => 
        HIEFFPLA_NET_0_118677);
    
    HIEFFPLA_INST_0_42340 : AND2A
      port map(A => HIEFFPLA_NET_0_119275, B => 
        \U50_PATTERNS/RD_USB_ADBUS[6]\, Y => 
        HIEFFPLA_NET_0_119566);
    
    \U_EXEC_MASTER/PRESCALE[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117766, CLK => CLK_40M_GL, CLR
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i\, Q => 
        \U_EXEC_MASTER/PRESCALE[2]\);
    
    \U200B_ELINKS/RX_SER_WORD_1DEL[6]\ : DFN1C0
      port map(D => \ELK_RX_SER_WORD_0[6]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_23, Q => 
        \U200B_ELINKS/RX_SER_WORD_1DEL[6]_net_1\);
    
    HIEFFPLA_INST_0_57617 : NAND3A
      port map(A => HIEFFPLA_NET_0_116645, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_5[7]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_5[6]\, Y => 
        HIEFFPLA_NET_0_116651);
    
    \U_ELK15_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]\ : DFN1C0
      port map(D => \U_ELK15_CH/U_SLAVE_1ELK/Q[2]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]_net_1\);
    
    \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[2]\ : DFN1C0
      port map(D => \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\);
    
    \U_ELK12_CH/U_SLAVE_1ELK/RECD_SER_WORD[2]\ : DFN1C0
      port map(D => \U_ELK12_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[2]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_12[2]\);
    
    HIEFFPLA_INST_0_55981 : MX2
      port map(A => HIEFFPLA_NET_0_116151, B => 
        HIEFFPLA_NET_0_116056, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[3]\, Y => 
        HIEFFPLA_NET_0_116965);
    
    \U_ELK8_CH/U_ELK1_SERDAT_SOURCE/SERDAT[5]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117873, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_5, Q => 
        \U_ELK8_CH/ELK_TX_DAT[5]\);
    
    AFLSDF_INV_50 : INV
      port map(A => DCB_SALT_SEL_c, Y => \AFLSDF_INV_50\);
    
    \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[5]\ : DFN1C0
      port map(D => 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\);
    
    HIEFFPLA_INST_0_161266 : DFN1C0
      port map(D => \U_ELK9_CH/U_ELK1_CMD_TX/START_RISE_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_0, Q
         => HIEFFPLA_NET_0_161289);
    
    \U_ELK18_CH/U_ELK1_CMD_TX/SER_OUT_RI\ : DFN1C0
      port map(D => 
        \U_ELK18_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_9, Q => 
        \U_ELK18_CH/U_ELK1_CMD_TX/SER_OUT_RI_net_1\);
    
    HIEFFPLA_INST_0_57869 : AXOI4
      port map(A => HIEFFPLA_NET_0_117085, B => 
        HIEFFPLA_NET_0_117113, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_7[0]\, Y => 
        HIEFFPLA_NET_0_116603);
    
    \U_ELK19_CH/U_SLAVE_1ELK/Q[2]\ : DFN1C0
      port map(D => \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/Q[2]_net_1\);
    
    HIEFFPLA_INST_0_50238 : MX2
      port map(A => HIEFFPLA_NET_0_117991, B => 
        HIEFFPLA_NET_0_118005, S => \BIT_OS_SEL_0[0]\, Y => 
        \U_ELK5_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[1]\);
    
    HIEFFPLA_INST_0_46067 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_7[7]\, C => 
        \U50_PATTERNS/SM_BANK_SEL[12]\, Y => 
        HIEFFPLA_NET_0_118774);
    
    HIEFFPLA_INST_0_40675 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_15[1]\, B => 
        HIEFFPLA_NET_0_119576, S => HIEFFPLA_NET_0_119297, Y => 
        HIEFFPLA_NET_0_119822);
    
    \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[14]\ : DFN1C0
      port map(D => 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]_net_1\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[14]_net_1\);
    
    \U50_PATTERNS/REG_ADDR[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119532, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_10, Q => \U50_PATTERNS/REG_ADDR[1]\);
    
    HIEFFPLA_INST_0_45868 : NAND2A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_4[4]\, Y => 
        HIEFFPLA_NET_0_118824);
    
    HIEFFPLA_INST_0_40097 : AOI1C
      port map(A => \U50_PATTERNS/ELINK_BLKA[13]\, B => 
        HIEFFPLA_NET_0_119657, C => HIEFFPLA_NET_0_119906, Y => 
        HIEFFPLA_NET_0_119907);
    
    \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_115924, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_9, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[6]\);
    
    HIEFFPLA_INST_0_57989 : XA1B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_7[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_7[0]\, C => 
        HIEFFPLA_NET_0_117179, Y => HIEFFPLA_NET_0_116583);
    
    HIEFFPLA_INST_0_57359 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_4[2]\, B => 
        HIEFFPLA_NET_0_116669, S => HIEFFPLA_NET_0_117122, Y => 
        HIEFFPLA_NET_0_116694);
    
    HIEFFPLA_INST_0_161277 : DFN1C0
      port map(D => \U_ELK0_CMD_TX/START_RISE_net_1\, CLK => 
        CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_17, Q => 
        HIEFFPLA_NET_0_161278);
    
    \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[2]\ : DFN1C0
      port map(D => 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[2]_net_1\);
    
    HIEFFPLA_INST_0_54800 : MX2
      port map(A => HIEFFPLA_NET_0_116335, B => 
        HIEFFPLA_NET_0_116390, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[3]_net_1\, Y => 
        HIEFFPLA_NET_0_117198);
    
    HIEFFPLA_INST_0_50425 : MX2
      port map(A => \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\, B
         => \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\, S => 
        \BIT_OS_SEL_5[2]\, Y => HIEFFPLA_NET_0_117952);
    
    \U50_PATTERNS/ELINK_DINA_6[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119736, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_16, Q => 
        \U50_PATTERNS/ELINK_DINA_6[7]\);
    
    \U_ELK17_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118332, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_14, Q => 
        \U_ELK17_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]_net_1\);
    
    \U50_PATTERNS/ELINK_DINA_8[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119720, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_18, Q => 
        \U50_PATTERNS/ELINK_DINA_8[7]\);
    
    HIEFFPLA_INST_0_46024 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/SM_BANK_SEL[3]\, C => 
        \U50_PATTERNS/ELINK_DOUTA_16[5]\, Y => 
        HIEFFPLA_NET_0_118784);
    
    HIEFFPLA_INST_0_57957 : NAND3
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_7[0]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_7[1]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_7[2]\, Y => 
        HIEFFPLA_NET_0_116592);
    
    HIEFFPLA_INST_0_47366 : MX2
      port map(A => 
        \U_ELK13_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]_net_1\, B => 
        \U_ELK13_CH/ELK_TX_DAT[7]\, S => 
        \U_ELK13_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118510);
    
    HIEFFPLA_INST_0_37282 : NAND3B
      port map(A => \U200A_TFC/GP_PG_SM[6]_net_1\, B => 
        \U200A_TFC/GP_PG_SM[7]_net_1\, C => 
        \U200A_TFC/GP_PG_SM[8]_net_1\, Y => HIEFFPLA_NET_0_120307);
    
    \U_ELK7_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]\ : DFN1C0
      port map(D => \U_ELK7_CH/U_SLAVE_1ELK/Q[2]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]_net_1\);
    
    HIEFFPLA_INST_0_56056 : AND3A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_0[8]_net_1\, B => 
        HIEFFPLA_NET_0_115873, C => HIEFFPLA_NET_0_117027, Y => 
        HIEFFPLA_NET_0_116955);
    
    HIEFFPLA_INST_0_62182 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_30[4]\, B => 
        HIEFFPLA_NET_0_117166, S => HIEFFPLA_NET_0_117330, Y => 
        HIEFFPLA_NET_0_116026);
    
    HIEFFPLA_INST_0_43359 : MX2
      port map(A => \U50_PATTERNS/SM_BANK_SEL[11]\, B => 
        HIEFFPLA_NET_0_119226, S => HIEFFPLA_NET_0_118691, Y => 
        HIEFFPLA_NET_0_119320);
    
    \U_ELK1_CH/U_SLAVE_1ELK/Q[2]\ : DFN1C0
      port map(D => \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/Q[2]_net_1\);
    
    HIEFFPLA_INST_0_53269 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_SEQCNT[1]\, B => 
        HIEFFPLA_NET_0_117436, S => HIEFFPLA_NET_0_117062, Y => 
        HIEFFPLA_NET_0_117441);
    
    HIEFFPLA_INST_0_41843 : AOI1B
      port map(A => HIEFFPLA_NET_0_119389, B => 
        \U50_PATTERNS/SM_BANK_SEL[4]\, C => HIEFFPLA_NET_0_119655, 
        Y => HIEFFPLA_NET_0_119685);
    
    HIEFFPLA_INST_0_51063 : MX2
      port map(A => \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\, 
        B => \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[14]_net_1\, S => 
        \BIT_OS_SEL_6[2]\, Y => HIEFFPLA_NET_0_117843);
    
    HIEFFPLA_INST_0_50511 : MX2
      port map(A => HIEFFPLA_NET_0_117951, B => 
        HIEFFPLA_NET_0_117950, S => \BIT_OS_SEL[0]\, Y => 
        \U_ELK6_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[4]\);
    
    \U_ELK17_CH/U_SLAVE_1ELK/RECD_SER_WORD[0]\ : DFN1C0
      port map(D => \U_ELK17_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[0]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_17[0]\);
    
    \U50_PATTERNS/U4A_REGCROSS/SAMP_TWO[1]\ : DFN1C0
      port map(D => \U50_PATTERNS/U4A_REGCROSS/SAMP_ONE[1]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_22, Q => 
        \U50_PATTERNS/U4A_REGCROSS/SAMP_TWO[1]_net_1\);
    
    HIEFFPLA_INST_0_47584 : MX2
      port map(A => 
        \U_ELK14_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]_net_1\, B => 
        \U_ELK14_CH/ELK_TX_DAT[2]\, S => 
        \U_ELK14_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118471);
    
    HIEFFPLA_INST_0_47491 : MX2
      port map(A => HIEFFPLA_NET_0_118476, B => 
        HIEFFPLA_NET_0_118494, S => \BIT_OS_SEL_4[0]\, Y => 
        \U_ELK13_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[0]\);
    
    HIEFFPLA_INST_0_46648 : MX2
      port map(A => \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\, 
        B => \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\, S => 
        \BIT_OS_SEL_5[2]\, Y => HIEFFPLA_NET_0_118633);
    
    HIEFFPLA_INST_0_53251 : AND2A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[8]_net_1\, B => 
        HIEFFPLA_NET_0_115871, Y => HIEFFPLA_NET_0_117445);
    
    \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[11]\ : DFN1C0
      port map(D => \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\);
    
    \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[7]\\\\/U0/U0\ : 
        IOPAD_BI_U
      port map(D => 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[7]\\\\/U0/NET1\, 
        E => 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[7]\\\\/U0/NET2\, 
        Y => 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[7]\\\\/U0/NET3\, 
        PAD => BIDIR_USB_ADBUS(7));
    
    HIEFFPLA_INST_0_40342 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_10[4]\, B => 
        HIEFFPLA_NET_0_119570, S => HIEFFPLA_NET_0_119239, Y => 
        HIEFFPLA_NET_0_119859);
    
    HIEFFPLA_INST_0_37575 : AND2
      port map(A => \TFC_ADDRB[1]\, B => HIEFFPLA_NET_0_120262, Y
         => HIEFFPLA_NET_0_120257);
    
    HIEFFPLA_INST_0_51089 : MX2
      port map(A => 
        \U_ELK9_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]_net_1\, B => 
        \U_ELK9_CH/ELK_TX_DAT[3]\, S => 
        \U_ELK9_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_117837);
    
    \U50_PATTERNS/ELINKS_STOP_ADDR_T[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120118, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_7, Q => 
        \U50_PATTERNS/ELINKS_STOP_ADDR_T[1]\);
    
    HIEFFPLA_INST_0_49314 : MX2
      port map(A => \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[0]_net_1\, B
         => \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\, S => 
        \BIT_OS_SEL[2]\, Y => HIEFFPLA_NET_0_118159);
    
    HIEFFPLA_INST_0_38714 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_12[0]\, B => 
        HIEFFPLA_NET_0_119524, S => HIEFFPLA_NET_0_119295, Y => 
        HIEFFPLA_NET_0_120071);
    
    \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[9]\ : DFN1C0
      port map(D => 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\);
    
    HIEFFPLA_INST_0_44552 : MX2
      port map(A => \ELKS_STOP_ADDR[0]\, B => 
        \U50_PATTERNS/U4D_REGCROSS/SAMP_TWO[0]_net_1\, S => 
        HIEFFPLA_NET_0_119093, Y => HIEFFPLA_NET_0_119091);
    
    HIEFFPLA_INST_0_39623 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_5[5]\, B => 
        HIEFFPLA_NET_0_119518, S => HIEFFPLA_NET_0_119251, Y => 
        HIEFFPLA_NET_0_119970);
    
    HIEFFPLA_INST_0_53723 : AND3C
      port map(A => HIEFFPLA_NET_0_117110, B => 
        HIEFFPLA_NET_0_117370, C => HIEFFPLA_NET_0_117364, Y => 
        HIEFFPLA_NET_0_117365);
    
    HIEFFPLA_INST_0_63208 : MX2
      port map(A => \U_TFC_CMD_TX/SER_CMD_WORD_F[1]_net_1\, B => 
        \TFC_TX_DAT[4]\, S => \U_TFC_CMD_TX/START_RISE_net_1\, Y
         => \U_TFC_CMD_TX/N_SER_CMD_WORD_F[2]\);
    
    \U50_PATTERNS/U4E_REGCROSS/LOCAL_REG_VAL[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119070, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_6, Q => \OP_MODE[0]\);
    
    HIEFFPLA_INST_0_43413 : MX2
      port map(A => \U50_PATTERNS/SM_BANK_SEL[17]\, B => 
        HIEFFPLA_NET_0_119220, S => HIEFFPLA_NET_0_118691, Y => 
        HIEFFPLA_NET_0_119314);
    
    HIEFFPLA_INST_0_41828 : AOI1B
      port map(A => HIEFFPLA_NET_0_119389, B => 
        \U50_PATTERNS/SM_BANK_SEL[7]\, C => HIEFFPLA_NET_0_119660, 
        Y => HIEFFPLA_NET_0_119688);
    
    \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[5]\ : DFN1C0
      port map(D => \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\);
    
    \U_ELK16_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]\ : DFN1C0
      port map(D => \U_ELK16_CH/U_SLAVE_1ELK/Q[6]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]_net_1\);
    
    \U_ELK3_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118108, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_12, Q => 
        \U_ELK3_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]_net_1\);
    
    HIEFFPLA_INST_0_56843 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_1[2]\, B => 
        HIEFFPLA_NET_0_116766, S => HIEFFPLA_NET_0_117600, Y => 
        HIEFFPLA_NET_0_116786);
    
    HIEFFPLA_INST_0_61358 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_5[0]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_21[0]\, S
         => \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_1[4]_net_1\, 
        Y => HIEFFPLA_NET_0_116138);
    
    HIEFFPLA_INST_0_52998 : MX2
      port map(A => HIEFFPLA_NET_0_117462, B => 
        HIEFFPLA_NET_0_117458, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[2]\, Y => 
        HIEFFPLA_NET_0_117478);
    
    HIEFFPLA_INST_0_50714 : MX2
      port map(A => \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\, B
         => \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[13]_net_1\, S => 
        \BIT_OS_SEL_5[2]\, Y => HIEFFPLA_NET_0_117901);
    
    HIEFFPLA_INST_0_43506 : MX2
      port map(A => \U50_PATTERNS/SM_BANK_SEL[7]\, B => 
        HIEFFPLA_NET_0_119211, S => HIEFFPLA_NET_0_118691, Y => 
        HIEFFPLA_NET_0_119303);
    
    \U50_PATTERNS/ELINKS_STRT_ADDR_T[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120097, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_21, Q => 
        \U50_PATTERNS/ELINKS_STRT_ADDR_T[6]\);
    
    HIEFFPLA_INST_0_37292 : AND3B
      port map(A => HIEFFPLA_NET_0_120291, B => 
        \U200A_TFC/GP_PG_SM[9]_net_1\, C => \OP_MODE_c[2]\, Y => 
        HIEFFPLA_NET_0_120302);
    
    HIEFFPLA_INST_0_161269 : DFN1C0
      port map(D => 
        \U_ELK16_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_10, Q
         => HIEFFPLA_NET_0_161286);
    
    \U_ELK16_CH/U_SLAVE_1ELK/Q[8]\ : DFN1C0
      port map(D => \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/Q[8]_net_1\);
    
    HIEFFPLA_INST_0_50821 : MX2
      port map(A => 
        \U_ELK8_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]_net_1\, B => 
        \U_ELK8_CH/ELK_TX_DAT[2]\, S => 
        \U_ELK8_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_117886);
    
    HIEFFPLA_INST_0_39461 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_3[3]\, B => 
        HIEFFPLA_NET_0_119520, S => HIEFFPLA_NET_0_119247, Y => 
        HIEFFPLA_NET_0_119988);
    
    HIEFFPLA_INST_0_37649 : NAND2B
      port map(A => \U200B_ELINKS/LOC_STRT_ADDR[5]\, B => 
        HIEFFPLA_NET_0_120190, Y => HIEFFPLA_NET_0_120240);
    
    HIEFFPLA_INST_0_53398 : AND2B
      port map(A => HIEFFPLA_NET_0_117325, B => 
        HIEFFPLA_NET_0_117390, Y => HIEFFPLA_NET_0_117414);
    
    \U_MASTER_DES/U13C_MASTER_DESER/ARB_WRD_40M_FIXED[0]\ : 
        DFN1C0
      port map(D => \U_MASTER_DES/U13C_MASTER_DESER/Q[0]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_26, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_WRD_40M_FIXED[0]_net_1\);
    
    HIEFFPLA_INST_0_42036 : AND3
      port map(A => \U50_PATTERNS/TFC_DOUTA[1]\, B => 
        HIEFFPLA_NET_0_118997, C => HIEFFPLA_NET_0_119365, Y => 
        HIEFFPLA_NET_0_119626);
    
    HIEFFPLA_INST_0_38482 : MX2
      port map(A => \U50_PATTERNS/ELINKS_STRT_ADDR_T[6]\, B => 
        \U50_PATTERNS/RD_USB_ADBUS[6]\, S => 
        HIEFFPLA_NET_0_119493, Y => HIEFFPLA_NET_0_120097);
    
    HIEFFPLA_INST_0_111369 : MX2B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_16[3]\, B => 
        HIEFFPLA_NET_0_115839, S => HIEFFPLA_NET_0_117215, Y => 
        HIEFFPLA_NET_0_116505);
    
    \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[10]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_115933, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_21, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[10]\);
    
    HIEFFPLA_INST_0_59588 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_13[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_29[1]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[4]_net_1\, Y => 
        HIEFFPLA_NET_0_116374);
    
    \U_ELK16_CH/U_SLAVE_1ELK/Q[12]\ : DFN1C0
      port map(D => \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/Q[12]_net_1\);
    
    HIEFFPLA_INST_0_51811 : AND3A
      port map(A => HIEFFPLA_NET_0_117685, B => 
        HIEFFPLA_NET_0_117686, C => HIEFFPLA_NET_0_117681, Y => 
        HIEFFPLA_NET_0_117689);
    
    \U_ELK16_CH/U_SLAVE_1ELK/Q[5]\ : DFN1C0
      port map(D => \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/Q[5]_net_1\);
    
    HIEFFPLA_INST_0_61742 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_9[2]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_25[2]\, S
         => \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_3[4]_net_1\, 
        Y => HIEFFPLA_NET_0_116084);
    
    HIEFFPLA_INST_0_47242 : MX2
      port map(A => HIEFFPLA_NET_0_118521, B => 
        HIEFFPLA_NET_0_118540, S => \BIT_OS_SEL_5[0]\, Y => 
        \U_ELK12_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[0]\);
    
    HIEFFPLA_INST_0_37623 : AND3B
      port map(A => HIEFFPLA_NET_0_120149, B => 
        \U200B_ELINKS/GP_PG_SM[10]_net_1\, C => 
        HIEFFPLA_NET_0_120220, Y => HIEFFPLA_NET_0_120244);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_24[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116105, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_8, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_24[0]\);
    
    \U_ELK3_CH/U_ELK1_SERDAT_SOURCE/SERDAT[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118103, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_14, Q => 
        \U_ELK3_CH/ELK_TX_DAT[0]\);
    
    HIEFFPLA_INST_0_52063 : AND2A
      port map(A => \U_MASTER_DES/U13A_ADJ_160M/BITCNT[0]\, B => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[2]_net_1\, Y => 
        HIEFFPLA_NET_0_117643);
    
    \U_ELK2_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL\ : DFN1C0
      port map(D => 
        \U_ELK2_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL_net_1\);
    
    HIEFFPLA_INST_0_56176 : XA1C
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/MAX_CNT[3]\, 
        B => HIEFFPLA_NET_0_116942, C => HIEFFPLA_NET_0_117112, Y
         => HIEFFPLA_NET_0_116936);
    
    \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[4]\ : DFN1C0
      port map(D => 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\);
    
    HIEFFPLA_INST_0_43102 : NAND3
      port map(A => \U50_PATTERNS/REG_STATE[2]_net_1\, B => 
        \U50_PATTERNS/REG_STATE[0]_net_1\, C => 
        \U50_PATTERNS/REG_STATE[1]_net_1\, Y => 
        HIEFFPLA_NET_0_119376);
    
    HIEFFPLA_INST_0_111190 : AOI1B
      port map(A => HIEFFPLA_NET_0_115848, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[0]_net_1\, C => 
        HIEFFPLA_NET_0_117103, Y => HIEFFPLA_NET_0_117081);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_20[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116466, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_13, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_20[1]\);
    
    HIEFFPLA_INST_0_59862 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_31[2]\, B => 
        HIEFFPLA_NET_0_116687, S => HIEFFPLA_NET_0_117097, Y => 
        HIEFFPLA_NET_0_116341);
    
    HIEFFPLA_INST_0_44256 : MX2
      port map(A => \TFC_STRT_ADDR[2]\, B => 
        \U50_PATTERNS/U4A_REGCROSS/SAMP_TWO[2]_net_1\, S => 
        HIEFFPLA_NET_0_119156, Y => HIEFFPLA_NET_0_119152);
    
    HIEFFPLA_INST_0_55414 : MX2
      port map(A => HIEFFPLA_NET_0_116955, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[4]\, S => 
        HIEFFPLA_NET_0_117087, Y => HIEFFPLA_NET_0_117041);
    
    \U_DDR_ELK0/BIBUF_LVDS_0/U0/U1\ : IOBI_ID_OD_EB
      port map(DR => ELK0_OUT_R_i_0, DF => ELK0_OUT_F_i_0, CLR
         => \GND\, E => \AFLSDF_INV_12\, ICLK => CCC_160M_ADJ, 
        OCLK => CCC_160M_FXD, YIN => 
        \U_DDR_ELK0/BIBUF_LVDS_0/U0/NET4\, DOUT => 
        \U_DDR_ELK0/BIBUF_LVDS_0/U0/NET1\, EOUT => 
        \U_DDR_ELK0/BIBUF_LVDS_0/U0/NET2\, YR => 
        \U_DDR_ELK0/ELK0_IN_DDR_R\, YF => 
        \U_DDR_ELK0/ELK0_IN_DDR_F\);
    
    \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[0]\ : DFN1C0
      port map(D => 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[0]_net_1\);
    
    \U50_PATTERNS/U4C_REGCROSS/LOCAL_REG_VAL[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119106, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_21, Q => \ELKS_STRT_ADDR[6]\);
    
    \U_ELK18_CH/U_ELK1_SERDAT_SOURCE/SERDAT[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118282, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_13, Q => 
        \U_ELK18_CH/ELK_TX_DAT[1]\);
    
    HIEFFPLA_INST_0_54940 : AOI1D
      port map(A => HIEFFPLA_NET_0_117349, B => 
        HIEFFPLA_NET_0_117410, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_3[6]_net_1\, Y => 
        HIEFFPLA_NET_0_117164);
    
    HIEFFPLA_INST_0_43242 : AND3B
      port map(A => \U50_PATTERNS/REG_STATE_0[1]_net_1\, B => 
        \U50_PATTERNS/USB_TXE_B\, C => HIEFFPLA_NET_0_119424, Y
         => HIEFFPLA_NET_0_119340);
    
    HIEFFPLA_INST_0_58059 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_0[2]\, B => 
        HIEFFPLA_NET_0_116564, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_1[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116570);
    
    \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[4]\ : DFN1C0
      port map(D => \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\);
    
    HIEFFPLA_INST_0_57446 : NAND3C
      port map(A => HIEFFPLA_NET_0_116770, B => 
        HIEFFPLA_NET_0_116586, C => HIEFFPLA_NET_0_116676, Y => 
        HIEFFPLA_NET_0_116680);
    
    \U50_PATTERNS/TFC_STRT_ADDR_T[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119161, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_4, Q => 
        \U50_PATTERNS/TFC_STRT_ADDR_T[3]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_19[4]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116176, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_11, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_19[4]\);
    
    \U_ELK2_CH/U_SLAVE_1ELK/Q[13]\ : DFN1C0
      port map(D => \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[13]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/Q[13]_net_1\);
    
    \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[3]\ : DFN1C0
      port map(D => \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\);
    
    HIEFFPLA_INST_0_45781 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_9[1]\, C => 
        \U50_PATTERNS/SM_BANK_SEL[10]\, Y => 
        HIEFFPLA_NET_0_118844);
    
    \U50_PATTERNS/ELINK_ADDRA_18[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120019, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_12, Q => 
        \U50_PATTERNS/ELINK_ADDRA_18[4]\);
    
    HIEFFPLA_INST_0_54568 : NAND2B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[4]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[2]_net_1\, Y => 
        HIEFFPLA_NET_0_117245);
    
    HIEFFPLA_INST_0_43719 : AND2B
      port map(A => HIEFFPLA_NET_0_119230, B => 
        \U50_PATTERNS/SM_BANK_SEL[1]\, Y => HIEFFPLA_NET_0_119233);
    
    \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[3]\ : DFN1C0
      port map(D => \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\);
    
    HIEFFPLA_INST_0_44434 : XOR2
      port map(A => \TFC_STOP_ADDR[1]\, B => 
        \U50_PATTERNS/U4B_REGCROSS/SAMP_TWO[1]_net_1\, Y => 
        HIEFFPLA_NET_0_119118);
    
    HIEFFPLA_INST_0_38696 : MX2
      port map(A => HIEFFPLA_NET_0_119517, B => 
        \U50_PATTERNS/ELINK_ADDRA_11[6]\, S => 
        HIEFFPLA_NET_0_119280, Y => HIEFFPLA_NET_0_120073);
    
    \U200A_TFC/RX_SER_WORD_2DEL[7]\ : DFN1C0
      port map(D => \U200A_TFC/RX_SER_WORD_1DEL[7]_net_1\, CLK
         => CLK_40M_GL, CLR => P_MASTER_POR_B_c, Q => 
        \U200A_TFC/RX_SER_WORD_2DEL[7]_net_1\);
    
    HIEFFPLA_INST_0_58827 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_1[0]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_17[0]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[4]_net_1\, Y
         => HIEFFPLA_NET_0_116471);
    
    \U_ELK18_CH/U_ELK1_CMD_TX/START_RISE\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118284, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_17, Q => 
        \U_ELK18_CH/U_ELK1_CMD_TX/START_RISE_net_1\);
    
    HIEFFPLA_INST_0_53446 : AND3
      port map(A => HIEFFPLA_NET_0_116740, B => 
        HIEFFPLA_NET_0_117360, C => HIEFFPLA_NET_0_117414, Y => 
        HIEFFPLA_NET_0_117407);
    
    HIEFFPLA_INST_0_48728 : MX2
      port map(A => HIEFFPLA_NET_0_118272, B => 
        HIEFFPLA_NET_0_118270, S => \BIT_OS_SEL_0[1]\, Y => 
        HIEFFPLA_NET_0_118260);
    
    HIEFFPLA_INST_0_57271 : NAND3C
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_3[4]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_3[8]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_3[5]\, Y => 
        HIEFFPLA_NET_0_116710);
    
    \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[44]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117709, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_33, Q => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[44]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_3[6]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117099, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_27_1, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_3[6]_net_1\);
    
    HIEFFPLA_INST_0_45182 : NAND3C
      port map(A => HIEFFPLA_NET_0_118798, B => 
        HIEFFPLA_NET_0_118876, C => HIEFFPLA_NET_0_118961, Y => 
        HIEFFPLA_NET_0_118970);
    
    \U_ELK11_CH/U_SLAVE_1ELK/RECD_SER_WORD[0]\ : DFN1C0
      port map(D => \U_ELK11_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[0]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_11[0]\);
    
    HIEFFPLA_INST_0_46482 : AND3B
      port map(A => HIEFFPLA_NET_0_119571, B => 
        \U50_PATTERNS/RD_USB_ADBUS[0]\, C => 
        HIEFFPLA_NET_0_119587, Y => HIEFFPLA_NET_0_118681);
    
    \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[1]\ : DFN1C0
      port map(D => 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[1]_net_1\);
    
    \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[12]\ : DFN1C0
      port map(D => 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[12]_net_1\);
    
    HIEFFPLA_INST_0_42494 : MX2
      port map(A => \U50_PATTERNS/REG_ADDR[6]\, B => 
        HIEFFPLA_NET_0_119503, S => HIEFFPLA_NET_0_119007, Y => 
        HIEFFPLA_NET_0_119527);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_2[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116367, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_18, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_2[0]\);
    
    HIEFFPLA_INST_0_37568 : AX1C
      port map(A => \TFC_ADDRB[6]\, B => HIEFFPLA_NET_0_120256, C
         => \TFC_ADDRB[7]\, Y => HIEFFPLA_NET_0_120259);
    
    HIEFFPLA_INST_0_51510 : NOR3B
      port map(A => \U_EXEC_MASTER/CCC_1_LOCK_STAT_1D_net_1\, B
         => HIEFFPLA_NET_0_117764, C => HIEFFPLA_NET_0_117756, Y
         => HIEFFPLA_NET_0_117759);
    
    HIEFFPLA_INST_0_44900 : AO1A
      port map(A => \U50_PATTERNS/USB_RXF_B\, B => 
        \U50_PATTERNS/REG_STATE[3]_net_1\, C => 
        \U50_PATTERNS/REG_STATE[0]_net_1\, Y => 
        HIEFFPLA_NET_0_119025);
    
    \U_ELK1_CH/U_SLAVE_1ELK/RECD_SER_WORD[0]\ : DFN1C0
      port map(D => \U_ELK1_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[0]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_1[0]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_18[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116187, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_8, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_18[3]\);
    
    HIEFFPLA_INST_0_51622 : MX2
      port map(A => 
        \U_EXEC_MASTER/USB_MASTER_EN/CNT_EN_60M2S_net_1\, B => 
        \U_EXEC_MASTER/USB_MASTER_EN/T_CNT60M[3]_net_1\, S => 
        HIEFFPLA_NET_0_117753, Y => HIEFFPLA_NET_0_117734);
    
    HIEFFPLA_INST_0_56601 : AND3
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[9]_net_1\, B => 
        HIEFFPLA_NET_0_117424, C => HIEFFPLA_NET_0_117427, Y => 
        HIEFFPLA_NET_0_116830);
    
    HIEFFPLA_INST_0_55564 : MX2
      port map(A => HIEFFPLA_NET_0_116199, B => 
        HIEFFPLA_NET_0_116090, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_1[3]\, Y => 
        HIEFFPLA_NET_0_117020);
    
    HIEFFPLA_INST_0_59063 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_23[2]\, B => 
        HIEFFPLA_NET_0_116436, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_1[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116440);
    
    HIEFFPLA_INST_0_45737 : AO1
      port map(A => HIEFFPLA_NET_0_119250, B => 
        \U50_PATTERNS/ELINK_DOUTA_5[6]\, C => 
        HIEFFPLA_NET_0_118770, Y => HIEFFPLA_NET_0_118855);
    
    \U_ELK5_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL\ : DFN1C0
      port map(D => \U_ELK5_CH/ELK_IN_R_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL_net_1\);
    
    HIEFFPLA_INST_0_58655 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_18[3]\, B => 
        HIEFFPLA_NET_0_116488, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_2[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116492);
    
    HIEFFPLA_INST_0_44869 : AO1A
      port map(A => HIEFFPLA_NET_0_119025, B => 
        HIEFFPLA_NET_0_119429, C => HIEFFPLA_NET_0_119024, Y => 
        HIEFFPLA_NET_0_119032);
    
    HIEFFPLA_INST_0_47322 : MX2
      port map(A => \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[0]_net_1\, 
        B => \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\, S => 
        \BIT_OS_SEL_3[2]\, Y => HIEFFPLA_NET_0_118519);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_3[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116339, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_19, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_3[0]\);
    
    \U50_PATTERNS/ELINK_DINA_14[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119825, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_16, Q => 
        \U50_PATTERNS/ELINK_DINA_14[6]\);
    
    \U_ELK10_CH/U_ELK1_SERDAT_SOURCE/SERDAT[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118643, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_17, Q => 
        \U_ELK10_CH/ELK_TX_DAT[0]\);
    
    \U_EXEC_MASTER/MPOR_B_2\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117787, CLK => CLK_40M_GL, CLR
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_2\, Q => 
        P_MASTER_POR_B_c_2);
    
    \U_ELK9_CH/U_SLAVE_1ELK/RECD_SER_WORD[0]\ : DFN1C0
      port map(D => \U_ELK9_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[0]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_9[0]\);
    
    HIEFFPLA_INST_0_60825 : MX2
      port map(A => HIEFFPLA_NET_0_117167, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_16[1]\, S => 
        HIEFFPLA_NET_0_117142, Y => HIEFFPLA_NET_0_116214);
    
    HIEFFPLA_INST_0_57993 : XA1C
      port map(A => HIEFFPLA_NET_0_116584, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_7[2]\, C => 
        HIEFFPLA_NET_0_117179, Y => HIEFFPLA_NET_0_116582);
    
    \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[3]\ : DFN1C0
      port map(D => \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\);
    
    HIEFFPLA_INST_0_49867 : NAND2B
      port map(A => \OP_MODE_c_1[1]\, B => \PATT_ELK_DAT_4[7]\, Y
         => HIEFFPLA_NET_0_118051);
    
    HIEFFPLA_INST_0_57722 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_6[2]\, B => 
        HIEFFPLA_NET_0_116614, S => HIEFFPLA_NET_0_117599, Y => 
        HIEFFPLA_NET_0_116630);
    
    HIEFFPLA_INST_0_47065 : MX2
      port map(A => HIEFFPLA_NET_0_118581, B => 
        HIEFFPLA_NET_0_118563, S => \BIT_OS_SEL_6[1]\, Y => 
        HIEFFPLA_NET_0_118565);
    
    \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[10]\ : DFN1C0
      port map(D => \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\);
    
    HIEFFPLA_INST_0_43591 : NAND2A
      port map(A => \U50_PATTERNS/SM_BANK_SEL[21]\, B => 
        HIEFFPLA_NET_0_119389, Y => HIEFFPLA_NET_0_119275);
    
    \U_ELK18_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118288, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_0, Q => 
        \U_ELK18_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]_net_1\);
    
    \U_ELK18_CH/U_SLAVE_1ELK/RECD_SER_WORD[4]\ : DFN1C0
      port map(D => \U_ELK18_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[4]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_18[4]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_115940, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_24, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[0]_net_1\);
    
    HIEFFPLA_INST_0_38029 : AOI1A
      port map(A => \ELKS_STRT_ADDR[6]\, B => 
        HIEFFPLA_NET_0_120219, C => HIEFFPLA_NET_0_120170, Y => 
        HIEFFPLA_NET_0_120171);
    
    \U50_PATTERNS/U4C_REGCROSS/SAMP_ONE[2]\ : DFN1C0
      port map(D => \U50_PATTERNS/ELINKS_STRT_ADDR[2]\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_33, Q => 
        \U50_PATTERNS/U4C_REGCROSS/SAMP_ONE[2]_net_1\);
    
    HIEFFPLA_INST_0_48194 : MX2
      port map(A => \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\, 
        B => \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[12]_net_1\, S => 
        \BIT_OS_SEL_1[2]\, Y => HIEFFPLA_NET_0_118355);
    
    \U_ELK2_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U1\ : IOBI_ID_OD_EB
      port map(DR => \U_ELK2_CH/ELK_OUT_R\, DF => 
        \U_ELK2_CH/ELK_OUT_F\, CLR => \GND\, E => \AFLSDF_INV_36\, 
        ICLK => CCC_160M_ADJ, OCLK => CCC_160M_FXD, YIN => 
        \U_ELK2_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\, DOUT => 
        \U_ELK2_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, EOUT => 
        \U_ELK2_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET2\, YR => 
        \U_ELK2_CH/ELK_IN_DDR_R\, YF => \U_ELK2_CH/ELK_IN_DDR_F\);
    
    HIEFFPLA_INST_0_56190 : AND3B
      port map(A => HIEFFPLA_NET_0_117112, B => 
        HIEFFPLA_NET_0_116930, C => HIEFFPLA_NET_0_116945, Y => 
        HIEFFPLA_NET_0_116933);
    
    HIEFFPLA_INST_0_48864 : AND2A
      port map(A => \OP_MODE_c_5[1]\, B => \PATT_ELK_DAT_19[0]\, 
        Y => HIEFFPLA_NET_0_118238);
    
    HIEFFPLA_INST_0_40166 : AOI1D
      port map(A => HIEFFPLA_NET_0_119389, B => 
        HIEFFPLA_NET_0_119464, C => 
        \U50_PATTERNS/SM_BANK_SEL[12]\, Y => 
        HIEFFPLA_NET_0_119883);
    
    HIEFFPLA_INST_0_48933 : MX2
      port map(A => HIEFFPLA_NET_0_118225, B => 
        HIEFFPLA_NET_0_118216, S => \BIT_OS_SEL_0[1]\, Y => 
        HIEFFPLA_NET_0_118222);
    
    HIEFFPLA_INST_0_44949 : AO1D
      port map(A => \U50_PATTERNS/TrienAux\, B => 
        HIEFFPLA_NET_0_119392, C => HIEFFPLA_NET_0_119452, Y => 
        HIEFFPLA_NET_0_119012);
    
    \U_ELK15_CH/U_SLAVE_1ELK/Q[14]\ : DFN1C0
      port map(D => \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[14]_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/Q[14]_net_1\);
    
    HIEFFPLA_INST_0_52299 : AND3A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[4]_net_1\, B => 
        HIEFFPLA_NET_0_117594, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[5]_net_1\, Y => 
        HIEFFPLA_NET_0_117587);
    
    \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[2]\ : DFN1C0
      port map(D => \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\);
    
    \U_ELK9_CH/U_SLAVE_1ELK/Q[1]\ : DFN1C0
      port map(D => \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/Q[1]_net_1\);
    
    \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[11]\ : DFN1C0
      port map(D => \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\);
    
    \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[7]\ : DFN1C0
      port map(D => 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\);
    
    HIEFFPLA_INST_0_49732 : MX2
      port map(A => HIEFFPLA_NET_0_118071, B => 
        HIEFFPLA_NET_0_118084, S => \BIT_OS_SEL_1[0]\, Y => 
        \U_ELK3_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[0]\);
    
    HIEFFPLA_INST_0_56497 : AO1
      port map(A => HIEFFPLA_NET_0_117428, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[9]_net_1\, C => 
        HIEFFPLA_NET_0_116835, Y => HIEFFPLA_NET_0_116851);
    
    HIEFFPLA_INST_0_42821 : AXOI5
      port map(A => \U50_PATTERNS/REG_STATE_0[1]_net_1\, B => 
        \U50_PATTERNS/REG_STATE[3]_net_1\, C => 
        \U50_PATTERNS/REG_STATE_0[2]_net_1\, Y => 
        HIEFFPLA_NET_0_119456);
    
    \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[2]\ : DFN1C0
      port map(D => 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[2]_net_1\);
    
    HIEFFPLA_INST_0_53589 : MX2
      port map(A => HIEFFPLA_NET_0_116463, B => 
        HIEFFPLA_NET_0_116379, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[3]_net_1\, Y
         => HIEFFPLA_NET_0_117385);
    
    HIEFFPLA_INST_0_46889 : MX2
      port map(A => \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\, 
        B => \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\, S => 
        \BIT_OS_SEL_4[2]\, Y => HIEFFPLA_NET_0_118589);
    
    \U200B_ELINKS/LOC_STOP_ADDR[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120182, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_7, Q => 
        \U200B_ELINKS/LOC_STOP_ADDR[5]\);
    
    HIEFFPLA_INST_0_52359 : AND2A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[8]_net_1\, B => 
        HIEFFPLA_NET_0_117572, Y => HIEFFPLA_NET_0_117576);
    
    HIEFFPLA_INST_0_49206 : MX2
      port map(A => \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\, B
         => \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[12]_net_1\, S => 
        \BIT_OS_SEL[2]\, Y => HIEFFPLA_NET_0_118173);
    
    HIEFFPLA_INST_0_45556 : AO1A
      port map(A => HIEFFPLA_NET_0_119622, B => 
        \U50_PATTERNS/TFC_STOP_ADDR[6]\, C => 
        HIEFFPLA_NET_0_118783, Y => HIEFFPLA_NET_0_118891);
    
    HIEFFPLA_INST_0_43813 : NAND3B
      port map(A => \U50_PATTERNS/RD_USB_ADBUS[4]\, B => 
        HIEFFPLA_NET_0_119585, C => 
        \U50_PATTERNS/RD_USB_ADBUS[5]\, Y => 
        HIEFFPLA_NET_0_119208);
    
    HIEFFPLA_INST_0_111809 : XA1A
      port map(A => HIEFFPLA_NET_0_115830, B => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[3]\, C => 
        HIEFFPLA_NET_0_117631, Y => HIEFFPLA_NET_0_117695);
    
    \U50_PATTERNS/RD_XFER_TYPE[7]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119542, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c, Q => 
        \U50_PATTERNS/RD_XFER_TYPE[7]_net_1\);
    
    HIEFFPLA_INST_0_39038 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_16[4]\, B => 
        HIEFFPLA_NET_0_119519, S => HIEFFPLA_NET_0_119257, Y => 
        HIEFFPLA_NET_0_120035);
    
    HIEFFPLA_INST_0_46468 : AOI1C
      port map(A => \U50_PATTERNS/WR_XFER_TYPE[4]_net_1\, B => 
        HIEFFPLA_NET_0_119577, C => HIEFFPLA_NET_0_118677, Y => 
        HIEFFPLA_NET_0_118685);
    
    \P_CCC_160M_ADJ_pad/U0/U0\ : IOPAD_TRI_U
      port map(D => \P_CCC_160M_ADJ_pad/U0/NET1\, E => 
        \P_CCC_160M_ADJ_pad/U0/NET2\, PAD => P_CCC_160M_ADJ);
    
    HIEFFPLA_INST_0_45028 : AND2
      port map(A => \U50_PATTERNS/REG_STATE[4]_net_1\, B => 
        \U50_PATTERNS/USB_TXE_B\, Y => HIEFFPLA_NET_0_118995);
    
    HIEFFPLA_INST_0_46016 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/SM_BANK_SEL[19]\, C => 
        \U50_PATTERNS/ELINK_DOUTA_0[1]\, Y => 
        HIEFFPLA_NET_0_118786);
    
    HIEFFPLA_INST_0_45751 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_7[1]\, C => 
        \U50_PATTERNS/SM_BANK_SEL[12]\, Y => 
        HIEFFPLA_NET_0_118852);
    
    HIEFFPLA_INST_0_61433 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_22[3]\, B => 
        HIEFFPLA_NET_0_117186, S => HIEFFPLA_NET_0_117080, Y => 
        HIEFFPLA_NET_0_116127);
    
    \U_ELK14_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U3\ : IOBI_ID_OD_EB
      port map(DR => \U_ELK14_CH/ELK_OUT_R\, DF => 
        \U_ELK14_CH/ELK_OUT_F\, CLR => \GND\, E => 
        \AFLSDF_INV_23\, ICLK => CCC_160M_ADJ, OCLK => 
        CCC_160M_FXD, YIN => 
        \U_ELK14_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\, DOUT => 
        OPEN, EOUT => 
        \U_ELK14_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET3\, YR => OPEN, 
        YF => OPEN);
    
    HIEFFPLA_INST_0_52914 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_23[2]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_24[2]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_2[0]\, Y => 
        HIEFFPLA_NET_0_117490);
    
    HIEFFPLA_INST_0_46572 : MX2
      port map(A => \U_ELK0_CMD_TX/SER_CMD_WORD_R[2]_net_1\, B
         => \ELK0_TX_DAT[7]\, S => 
        \U_ELK0_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118662);
    
    HIEFFPLA_INST_0_62968 : MX2
      port map(A => HIEFFPLA_NET_0_115887, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[7]\, S => 
        HIEFFPLA_NET_0_117073, Y => HIEFFPLA_NET_0_115923);
    
    HIEFFPLA_INST_0_60648 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_13[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_14[1]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_3[0]\, Y => 
        HIEFFPLA_NET_0_116238);
    
    HIEFFPLA_INST_0_161259 : DFN1C0
      port map(D => \ELK0_IN_R\, CLK => CCC_160M_ADJ, CLR => 
        P_MASTER_POR_B_c_26, Q => HIEFFPLA_NET_0_161296);
    
    \U_ELK4_CH/U_SLAVE_1ELK/RECD_SER_WORD[6]\ : DFN1C0
      port map(D => \U_ELK4_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[6]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_4[6]\);
    
    HIEFFPLA_INST_0_45646 : AO1
      port map(A => HIEFFPLA_NET_0_119241, B => 
        \U50_PATTERNS/ELINK_DOUTA_1[6]\, C => 
        HIEFFPLA_NET_0_118707, Y => HIEFFPLA_NET_0_118873);
    
    HIEFFPLA_INST_0_45152 : NAND3C
      port map(A => HIEFFPLA_NET_0_118804, B => 
        HIEFFPLA_NET_0_118881, C => HIEFFPLA_NET_0_118966, Y => 
        HIEFFPLA_NET_0_118977);
    
    HIEFFPLA_INST_0_42584 : XA1C
      port map(A => HIEFFPLA_NET_0_119514, B => 
        \U50_PATTERNS/REG_ADDR[3]\, C => HIEFFPLA_NET_0_119452, Y
         => HIEFFPLA_NET_0_119506);
    
    HIEFFPLA_INST_0_43098 : NAND2A
      port map(A => \U50_PATTERNS/REG_STATE[0]_net_1\, B => 
        \U50_PATTERNS/REG_STATE[1]_net_1\, Y => 
        HIEFFPLA_NET_0_119379);
    
    \U_ELK4_CH/U_SLAVE_1ELK/Q[9]\ : DFN1C0
      port map(D => \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/Q[9]_net_1\);
    
    \U_ELK1_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]\ : DFN1C0
      port map(D => \U_ELK1_CH/U_SLAVE_1ELK/Q[2]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]_net_1\);
    
    HIEFFPLA_INST_0_44376 : MX2
      port map(A => \TFC_STOP_ADDR[4]\, B => 
        \U50_PATTERNS/U4B_REGCROSS/SAMP_TWO[4]_net_1\, S => 
        HIEFFPLA_NET_0_119135, Y => HIEFFPLA_NET_0_119129);
    
    \U_ELK9_CH/U_SLAVE_1ELK/RECD_SER_WORD[6]\ : DFN1C0
      port map(D => \U_ELK9_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[6]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_9[6]\);
    
    HIEFFPLA_INST_0_54896 : AOI1C
      port map(A => HIEFFPLA_NET_0_117184, B => 
        HIEFFPLA_NET_0_117388, C => HIEFFPLA_NET_0_117207, Y => 
        HIEFFPLA_NET_0_117177);
    
    HIEFFPLA_INST_0_47911 : MX2
      port map(A => \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\, 
        B => \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\, S => 
        \BIT_OS_SEL_1[2]\, Y => HIEFFPLA_NET_0_118405);
    
    HIEFFPLA_INST_0_57317 : AND3B
      port map(A => HIEFFPLA_NET_0_116697, B => 
        HIEFFPLA_NET_0_117179, C => HIEFFPLA_NET_0_116709, Y => 
        HIEFFPLA_NET_0_116700);
    
    HIEFFPLA_INST_0_112590 : AO13
      port map(A => HIEFFPLA_NET_0_115836, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_SEQCNT[2]\, C => 
        HIEFFPLA_NET_0_116977, Y => HIEFFPLA_NET_0_115814);
    
    HIEFFPLA_INST_0_62418 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_5[3]\, 
        B => HIEFFPLA_NET_0_117075, S => HIEFFPLA_NET_0_117172, Y
         => HIEFFPLA_NET_0_115992);
    
    HIEFFPLA_INST_0_46352 : AO1
      port map(A => HIEFFPLA_NET_0_119290, B => 
        \U50_PATTERNS/ELINK_DOUTA_17[4]\, C => 
        HIEFFPLA_NET_0_118709, Y => HIEFFPLA_NET_0_118710);
    
    \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[6]\ : DFN1C0
      port map(D => \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_4[4]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_115996, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_13, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_4[4]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_1[4]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116784, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_4, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_1[4]\);
    
    \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[6]\ : DFN1C0
      port map(D => \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\);
    
    HIEFFPLA_INST_0_55041 : AOI1D
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[6]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[8]_net_1\, C => 
        HIEFFPLA_NET_0_116649, Y => HIEFFPLA_NET_0_117135);
    
    HIEFFPLA_INST_0_51105 : AND2A
      port map(A => \OP_MODE_c_3[1]\, B => \PATT_ELK_DAT_9[0]\, Y
         => HIEFFPLA_NET_0_117833);
    
    HIEFFPLA_INST_0_40450 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_12[0]\, B => 
        HIEFFPLA_NET_0_119578, S => HIEFFPLA_NET_0_119295, Y => 
        HIEFFPLA_NET_0_119847);
    
    \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[14]\ : DFN1C0
      port map(D => \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[14]_net_1\);
    
    \U50_PATTERNS/ELINK_DINA_11[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119848, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_11, Q => 
        \U50_PATTERNS/ELINK_DINA_11[7]\);
    
    HIEFFPLA_INST_0_38507 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_0[1]\, B => 
        HIEFFPLA_NET_0_119523, S => HIEFFPLA_NET_0_119272, Y => 
        HIEFFPLA_NET_0_120094);
    
    HIEFFPLA_INST_0_49346 : MX2
      port map(A => 
        \U_ELK2_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]_net_1\, B => 
        \U_ELK2_CH/ELK_TX_DAT[3]\, S => 
        \U_ELK2_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118152);
    
    \U_ELK5_CH/U_ELK1_CMD_TX/START_RISE\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118014, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_3, Q => 
        \U_ELK5_CH/U_ELK1_CMD_TX/START_RISE_net_1\);
    
    \U_ELK16_CH/U_ELK1_SERDAT_SOURCE/SERDAT[5]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118368, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_9, Q => 
        \U_ELK16_CH/ELK_TX_DAT[5]\);
    
    HIEFFPLA_INST_0_57665 : AND3B
      port map(A => HIEFFPLA_NET_0_117179, B => 
        HIEFFPLA_NET_0_116634, C => HIEFFPLA_NET_0_116645, Y => 
        HIEFFPLA_NET_0_116639);
    
    \U_ELK4_CH/U_SLAVE_1ELK/Q[0]\ : DFN1C0
      port map(D => \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/Q[0]_net_1\);
    
    \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[0]\ : DFN1C0
      port map(D => 
        \U_ELK13_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\);
    
    HIEFFPLA_INST_0_57998 : XA1C
      port map(A => HIEFFPLA_NET_0_116592, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_7[3]\, C => 
        HIEFFPLA_NET_0_117179, Y => HIEFFPLA_NET_0_116581);
    
    \U_ELK3_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]\ : DFN1C0
      port map(D => \U_ELK3_CH/U_SLAVE_1ELK/Q[7]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]_net_1\);
    
    HIEFFPLA_INST_0_62613 : MX2
      port map(A => HIEFFPLA_NET_0_117075, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_8[3]\, S => 
        HIEFFPLA_NET_0_117153, Y => HIEFFPLA_NET_0_115967);
    
    HIEFFPLA_INST_0_61508 : MX2
      port map(A => HIEFFPLA_NET_0_117186, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_23[3]\, S => 
        HIEFFPLA_NET_0_117151, Y => HIEFFPLA_NET_0_116117);
    
    HIEFFPLA_INST_0_46276 : NAND3B
      port map(A => HIEFFPLA_NET_0_118891, B => 
        HIEFFPLA_NET_0_118883, C => HIEFFPLA_NET_0_119427, Y => 
        HIEFFPLA_NET_0_118727);
    
    \U_ELK18_CH/U_SLAVE_1ELK/Q[13]\ : DFN1C0
      port map(D => \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[13]_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/Q[13]_net_1\);
    
    \U50_PATTERNS/REG_STATE_0[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119468, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_22_0, Q => 
        \U50_PATTERNS/REG_STATE_0[1]_net_1\);
    
    \U200B_ELINKS/RX_SER_WORD_3DEL[5]\ : DFN1C0
      port map(D => \U200B_ELINKS/RX_SER_WORD_2DEL[5]_net_1\, CLK
         => CLK_40M_GL, CLR => P_MASTER_POR_B_c_31_0, Q => 
        \U200B_ELINKS/RX_SER_WORD_3DEL[5]_net_1\);
    
    HIEFFPLA_INST_0_62853 : MX2
      port map(A => HIEFFPLA_NET_0_115879, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/TUNE_CLKPHASE[1]\, S => 
        HIEFFPLA_NET_0_117102, Y => HIEFFPLA_NET_0_115936);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_17[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116499, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_18, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_17[2]\);
    
    HIEFFPLA_INST_0_54245 : MX2
      port map(A => HIEFFPLA_NET_0_116565, B => 
        HIEFFPLA_NET_0_116287, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_1[3]_net_1\, Y
         => HIEFFPLA_NET_0_117290);
    
    HIEFFPLA_INST_0_58323 : AND3A
      port map(A => HIEFFPLA_NET_0_116532, B => 
        HIEFFPLA_NET_0_116530, C => HIEFFPLA_NET_0_117367, Y => 
        HIEFFPLA_NET_0_116534);
    
    HIEFFPLA_INST_0_43143 : AO1
      port map(A => HIEFFPLA_NET_0_119584, B => 
        HIEFFPLA_NET_0_119348, C => HIEFFPLA_NET_0_119346, Y => 
        HIEFFPLA_NET_0_119361);
    
    HIEFFPLA_INST_0_58124 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_10[1]\, B => 
        HIEFFPLA_NET_0_116677, S => HIEFFPLA_NET_0_117165, Y => 
        HIEFFPLA_NET_0_116561);
    
    HIEFFPLA_INST_0_41323 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_5[1]\, B => 
        HIEFFPLA_NET_0_119576, S => HIEFFPLA_NET_0_119251, Y => 
        HIEFFPLA_NET_0_119750);
    
    \U_ELK8_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL\ : DFN1C0
      port map(D => 
        \U_ELK8_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL_net_1\);
    
    \U_EXEC_MASTER/MPOR_B_22_0\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117787, CLK => CLK_40M_GL, CLR
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_0\, Q => 
        P_MASTER_POR_B_c_22_0);
    
    \U_ELK18_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]\ : DFN1C0
      port map(D => \U_ELK18_CH/U_SLAVE_1ELK/Q[4]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]_net_1\);
    
    HIEFFPLA_INST_0_111799 : OR3B
      port map(A => \U_MASTER_DES/U13A_ADJ_160M/BITCNT[3]\, B => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[1]\, C => 
        HIEFFPLA_NET_0_117682, Y => HIEFFPLA_NET_0_115831);
    
    \U_ELK17_CH/U_ELK1_CMD_TX/SER_OUT_FDEL\ : DFN1C0
      port map(D => \U_ELK17_CH/U_ELK1_CMD_TX/SER_OUT_FI_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_12, Q
         => \U_ELK17_CH/ELK_OUT_F\);
    
    \U50_PATTERNS/ELINK_ADDRA_16[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120033, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_9, Q => 
        \U50_PATTERNS/ELINK_ADDRA_16[6]\);
    
    HIEFFPLA_INST_0_53942 : AO1C
      port map(A => HIEFFPLA_NET_0_117107, B => 
        HIEFFPLA_NET_0_117328, C => HIEFFPLA_NET_0_117086, Y => 
        HIEFFPLA_NET_0_117330);
    
    HIEFFPLA_INST_0_46640 : MX2
      port map(A => HIEFFPLA_NET_0_118633, B => 
        HIEFFPLA_NET_0_118628, S => \BIT_OS_SEL_5[1]\, Y => 
        HIEFFPLA_NET_0_118634);
    
    HIEFFPLA_INST_0_40936 : MX2
      port map(A => HIEFFPLA_NET_0_119566, B => 
        \U50_PATTERNS/ELINK_DINA_18[6]\, S => 
        HIEFFPLA_NET_0_119264, Y => HIEFFPLA_NET_0_119793);
    
    \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[14]\ : DFN1C0
      port map(D => \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[14]_net_1\);
    
    HIEFFPLA_INST_0_51548 : AND2
      port map(A => HIEFFPLA_NET_0_117746, B => 
        \U_EXEC_MASTER/USB_MASTER_EN/T_CNT60M[3]_net_1\, Y => 
        HIEFFPLA_NET_0_117747);
    
    HIEFFPLA_INST_0_49366 : AND2A
      port map(A => \OP_MODE_c_1[1]\, B => \PATT_ELK_DAT_2[4]\, Y
         => HIEFFPLA_NET_0_118144);
    
    HIEFFPLA_INST_0_45007 : AND3A
      port map(A => \U50_PATTERNS/REG_STATE_0[2]_net_1\, B => 
        \U50_PATTERNS/USB_TXE_B\, C => 
        \U50_PATTERNS/REG_STATE_0[1]_net_1\, Y => 
        HIEFFPLA_NET_0_119001);
    
    HIEFFPLA_INST_0_37642 : AND3B
      port map(A => \U200B_ELINKS/LOC_STRT_ADDR[3]\, B => 
        HIEFFPLA_NET_0_120190, C => HIEFFPLA_NET_0_120234, Y => 
        HIEFFPLA_NET_0_120241);
    
    \U50_PATTERNS/ELINK_DINA_7[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119734, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_17, Q => 
        \U50_PATTERNS/ELINK_DINA_7[1]\);
    
    HIEFFPLA_INST_0_56799 : XA1C
      port map(A => HIEFFPLA_NET_0_116801, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_0[6]\, C => 
        HIEFFPLA_NET_0_117179, Y => HIEFFPLA_NET_0_116794);
    
    \U_ELK12_CH/U_SLAVE_1ELK/Q[11]\ : DFN1C0
      port map(D => \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/Q[11]_net_1\);
    
    \U_ELK3_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118105, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_12, Q => 
        \U_ELK3_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]_net_1\);
    
    HIEFFPLA_INST_0_55322 : AND2A
      port map(A => HIEFFPLA_NET_0_117027, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[4]_net_1\, Y => 
        HIEFFPLA_NET_0_117060);
    
    \U200B_ELINKS/RX_SER_WORD_3DEL[3]\ : DFN1P0
      port map(D => \AFLSDF_INV_60\, CLK => CLK_40M_GL, PRE => 
        P_MASTER_POR_B_c_31_0, Q => 
        \U200B_ELINKS/RX_SER_WORD_3DEL_i_0[3]\);
    
    HIEFFPLA_INST_0_55027 : AO1B
      port map(A => HIEFFPLA_NET_0_117337, B => 
        HIEFFPLA_NET_0_117147, C => HIEFFPLA_NET_0_117086, Y => 
        HIEFFPLA_NET_0_117138);
    
    HIEFFPLA_INST_0_50919 : MX2
      port map(A => \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[3]_net_1\, B
         => \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\, S => 
        \BIT_OS_SEL_3[2]\, Y => HIEFFPLA_NET_0_117863);
    
    HIEFFPLA_INST_0_43317 : AND2A
      port map(A => HIEFFPLA_NET_0_119328, B => 
        HIEFFPLA_NET_0_119443, Y => HIEFFPLA_NET_0_119327);
    
    HIEFFPLA_INST_0_48160 : MX2
      port map(A => \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\, 
        B => \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\, S => 
        \BIT_OS_SEL_1[2]\, Y => HIEFFPLA_NET_0_118360);
    
    HIEFFPLA_INST_0_46031 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_9[7]\, C => 
        \U50_PATTERNS/SM_BANK_SEL[10]\, Y => 
        HIEFFPLA_NET_0_118782);
    
    HIEFFPLA_INST_0_44030 : MX2
      port map(A => \U50_PATTERNS/TFC_STOP_ADDR[6]\, B => 
        \U50_PATTERNS/TFC_STOP_ADDR_T[6]\, S => 
        HIEFFPLA_NET_0_119472, Y => HIEFFPLA_NET_0_119182);
    
    \U200A_TFC/GP_PG_SM[10]\ : DFN1P0
      port map(D => HIEFFPLA_NET_0_120335, CLK => CLK_40M_GL, PRE
         => P_MASTER_POR_B_c_27_1, Q => 
        \U200A_TFC/GP_PG_SM[10]_net_1\);
    
    HIEFFPLA_INST_0_37557 : AND2
      port map(A => \TFC_ADDRB[4]\, B => HIEFFPLA_NET_0_120258, Y
         => HIEFFPLA_NET_0_120260);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_1[7]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116781, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_4, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_1[7]\);
    
    \U200B_ELINKS/RX_SER_WORD_3DEL[1]\ : DFN1P0
      port map(D => \AFLSDF_INV_61\, CLK => CLK_40M_GL, PRE => 
        P_MASTER_POR_B_c_31_0, Q => 
        \U200B_ELINKS/RX_SER_WORD_3DEL_i_0[1]\);
    
    HIEFFPLA_INST_0_58106 : MX2
      port map(A => HIEFFPLA_NET_0_116815, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_0[3]\, S => 
        HIEFFPLA_NET_0_117201, Y => HIEFFPLA_NET_0_116563);
    
    HIEFFPLA_INST_0_59986 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_4[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_20[1]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_2[4]_net_1\, Y
         => HIEFFPLA_NET_0_116325);
    
    HIEFFPLA_INST_0_44340 : AND2A
      port map(A => \U50_PATTERNS/U4B_REGCROSS/DELCNT[0]_net_1\, 
        B => \U50_PATTERNS/U4B_REGCROSS/SYNC_SM[0]_net_1\, Y => 
        HIEFFPLA_NET_0_119134);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_7[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_115978, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_17_0, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_7[2]\);
    
    \U200A_TFC/RX_SER_WORD_1DEL[5]\ : DFN1C0
      port map(D => \TFC_RX_SER_WORD[5]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_31, Q => 
        \U200A_TFC/RX_SER_WORD_1DEL[5]_net_1\);
    
    HIEFFPLA_INST_0_63024 : NAND2B
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[13]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[11]\, Y => 
        HIEFFPLA_NET_0_115911);
    
    HIEFFPLA_INST_0_54837 : AO1C
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_0[8]_net_1\, B => 
        HIEFFPLA_NET_0_117192, C => HIEFFPLA_NET_0_117104, Y => 
        HIEFFPLA_NET_0_117193);
    
    HIEFFPLA_INST_0_53363 : MX2
      port map(A => HIEFFPLA_NET_0_117262, B => 
        HIEFFPLA_NET_0_117387, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[2]_net_1\, Y
         => HIEFFPLA_NET_0_117420);
    
    AFLSDF_INV_5 : INV
      port map(A => P_USB_MASTER_EN_c_22, Y => \AFLSDF_INV_5\);
    
    HIEFFPLA_INST_0_61082 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_19[4]\, B => 
        HIEFFPLA_NET_0_117100, S => HIEFFPLA_NET_0_117170, Y => 
        HIEFFPLA_NET_0_116176);
    
    \U_EXEC_MASTER/DEL_CNT[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117793, CLK => CLK_40M_GL, CLR
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i\, Q => 
        \U_EXEC_MASTER/DEL_CNT[2]\);
    
    HIEFFPLA_INST_0_52908 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_23[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_24[1]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_2[0]\, Y => 
        HIEFFPLA_NET_0_117491);
    
    HIEFFPLA_INST_0_113977 : AO18
      port map(A => HIEFFPLA_NET_0_115807, B => \TFC_ADDRB[2]\, C
         => \U200A_TFC/LOC_STOP_ADDR[2]\, Y => 
        HIEFFPLA_NET_0_115811);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_5[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_115995, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_15, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_5[0]\);
    
    \U_ELK1_CH/U_ELK1_SERDAT_SOURCE/SERDAT[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118191, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_11, Q => 
        \U_ELK1_CH/ELK_TX_DAT[2]\);
    
    HIEFFPLA_INST_0_48029 : MX2
      port map(A => HIEFFPLA_NET_0_118404, B => 
        HIEFFPLA_NET_0_118400, S => \BIT_OS_SEL_3[0]\, Y => 
        \U_ELK15_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[5]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_0[5]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116819, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_3, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_0[5]\);
    
    \U50_PATTERNS/RD_XFER_TYPE[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119549, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c, Q => 
        \U50_PATTERNS/RD_XFER_TYPE[0]_net_1\);
    
    HIEFFPLA_INST_0_53392 : AND2
      port map(A => HIEFFPLA_NET_0_117334, B => 
        HIEFFPLA_NET_0_117380, Y => HIEFFPLA_NET_0_117416);
    
    HIEFFPLA_INST_0_44902 : AND3B
      port map(A => HIEFFPLA_NET_0_119449, B => 
        \U50_PATTERNS/REG_STATE_0[5]_net_1\, C => 
        \U50_PATTERNS/REG_STATE[0]_net_1\, Y => 
        HIEFFPLA_NET_0_119024);
    
    \U_ELK6_CH/U_SLAVE_1ELK/Q[12]\ : DFN1C0
      port map(D => \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/Q[12]_net_1\);
    
    \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[13]\ : DFN1C0
      port map(D => 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[13]_net_1\);
    
    HIEFFPLA_INST_0_41849 : AND2
      port map(A => HIEFFPLA_NET_0_119389, B => 
        \U50_PATTERNS/SM_BANK_SEL[3]\, Y => HIEFFPLA_NET_0_119683);
    
    HIEFFPLA_INST_0_37748 : AO1
      port map(A => \OP_MODE_c[6]\, B => 
        \U200B_ELINKS/GP_PG_SM[0]_net_1\, C => 
        \U200B_ELINKS/GP_PG_SM[1]_net_1\, Y => 
        HIEFFPLA_NET_0_120217);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_0[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116823, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_2, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_0[1]\);
    
    \U_ELK16_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U1\ : IOBI_ID_OD_EB
      port map(DR => \U_ELK16_CH/ELK_OUT_R\, DF => 
        \U_ELK16_CH/ELK_OUT_F\, CLR => \GND\, E => 
        \AFLSDF_INV_26\, ICLK => CCC_160M_ADJ, OCLK => 
        CCC_160M_FXD, YIN => 
        \U_ELK16_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\, DOUT => 
        \U_ELK16_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, EOUT => 
        \U_ELK16_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET2\, YR => 
        \U_ELK16_CH/ELK_IN_DDR_R\, YF => 
        \U_ELK16_CH/ELK_IN_DDR_F\);
    
    HIEFFPLA_INST_0_60654 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_13[2]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_14[2]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_3[0]\, Y => 
        HIEFFPLA_NET_0_116237);
    
    \U50_PATTERNS/U4D_REGCROSS/SAMP_TWO[1]\ : DFN1C0
      port map(D => \U50_PATTERNS/U4D_REGCROSS/SAMP_ONE[1]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_30, Q => 
        \U50_PATTERNS/U4D_REGCROSS/SAMP_TWO[1]_net_1\);
    
    \U50_PATTERNS/U4B_REGCROSS/SAMP_TWO[6]\ : DFN1C0
      port map(D => \U50_PATTERNS/U4B_REGCROSS/SAMP_ONE[6]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_29, Q => 
        \U50_PATTERNS/U4B_REGCROSS/SAMP_TWO[6]_net_1\);
    
    HIEFFPLA_INST_0_37727 : XO1
      port map(A => HIEFFPLA_NET_0_120144, B => \ELKS_ADDRB[6]\, 
        C => \U200B_ELINKS/GP_PG_SM[10]_net_1\, Y => 
        HIEFFPLA_NET_0_120221);
    
    HIEFFPLA_INST_0_112168 : AO13
      port map(A => HIEFFPLA_NET_0_115818, B => 
        \U200A_TFC/LOC_STOP_ADDR[4]\, C => \TFC_ADDRB[4]\, Y => 
        HIEFFPLA_NET_0_120294);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_6[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_115982, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_16, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_6[3]\);
    
    AFLSDF_INV_64 : INV
      port map(A => \U_ELK4_CH/U_DDR_ELK1/ELK_IN_DDR_F\, Y => 
        \AFLSDF_INV_64\);
    
    \U50_PATTERNS/U4C_REGCROSS/SAMP_TWO[6]\ : DFN1C0
      port map(D => \U50_PATTERNS/U4C_REGCROSS/SAMP_ONE[6]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_22_0, Q => 
        \U50_PATTERNS/U4C_REGCROSS/SAMP_TWO[6]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_0[6]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116818, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_3, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_0[6]\);
    
    HIEFFPLA_INST_0_53814 : AO1C
      port map(A => HIEFFPLA_NET_0_117329, B => 
        HIEFFPLA_NET_0_117116, C => HIEFFPLA_NET_0_117180, Y => 
        HIEFFPLA_NET_0_117348);
    
    \U50_PATTERNS/ELINK_BLKA[1]/U1\ : DFN1P0
      port map(D => HIEFFPLA_NET_0_119924, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_19, Q => 
        \U50_PATTERNS/ELINK_BLKA[1]\);
    
    \P_OP_MODE6_EE_pad/U0/U0\ : IOPAD_TRI_U
      port map(D => \P_OP_MODE6_EE_pad/U0/NET1\, E => 
        \P_OP_MODE6_EE_pad/U0/NET2\, PAD => P_OP_MODE6_EE);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_15[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116520, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_15, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_15[0]\);
    
    \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[2]\ : DFN1C0
      port map(D => \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\);
    
    HIEFFPLA_INST_0_44329 : XOR2
      port map(A => \TFC_STRT_ADDR[0]\, B => 
        \U50_PATTERNS/U4A_REGCROSS/SAMP_TWO[0]_net_1\, Y => 
        HIEFFPLA_NET_0_119140);
    
    HIEFFPLA_INST_0_38330 : MX2
      port map(A => \U50_PATTERNS/ELINKS_STOP_ADDR_T[3]\, B => 
        \U50_PATTERNS/RD_USB_ADBUS[3]\, S => 
        HIEFFPLA_NET_0_119413, Y => HIEFFPLA_NET_0_120116);
    
    HIEFFPLA_INST_0_46937 : MX2
      port map(A => HIEFFPLA_NET_0_118575, B => 
        HIEFFPLA_NET_0_118589, S => \BIT_OS_SEL_4[1]\, Y => 
        HIEFFPLA_NET_0_118582);
    
    \U200B_ELINKS/GP_PG_SM[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120217, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_29, Q => 
        \U200B_ELINKS/GP_PG_SM[0]_net_1\);
    
    HIEFFPLA_INST_0_51805 : AND3A
      port map(A => HIEFFPLA_NET_0_117682, B => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[5]\, C => 
        HIEFFPLA_NET_0_117686, Y => HIEFFPLA_NET_0_117690);
    
    \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[14]\ : DFN1C0
      port map(D => 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]_net_1\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[14]_net_1\);
    
    HIEFFPLA_INST_0_53907 : AND3A
      port map(A => HIEFFPLA_NET_0_117237, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[0]_net_1\, C
         => \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_1[3]_net_1\, 
        Y => HIEFFPLA_NET_0_117335);
    
    \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[3]\ : DFN1C0
      port map(D => \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\);
    
    HIEFFPLA_INST_0_56433 : AND3
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[7]_net_1\, B => 
        HIEFFPLA_NET_0_117427, C => HIEFFPLA_NET_0_117423, Y => 
        HIEFFPLA_NET_0_116868);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_0[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116821, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_3, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_0[3]\);
    
    \U_ELK6_CH/ELK_IN_R\ : DFN1C0
      port map(D => \U_ELK6_CH/ELK_IN_DDR_R\, CLK => CCC_160M_ADJ, 
        CLR => DEV_RST_B_c, Q => \U_ELK6_CH/ELK_IN_R_net_1\);
    
    HIEFFPLA_INST_0_50634 : MX2
      port map(A => HIEFFPLA_NET_0_117903, B => 
        HIEFFPLA_NET_0_117901, S => \BIT_OS_SEL_4[1]\, Y => 
        HIEFFPLA_NET_0_117913);
    
    HIEFFPLA_INST_0_47833 : MX2
      port map(A => 
        \U_ELK15_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]_net_1\, B => 
        \U_ELK15_CH/ELK_TX_DAT[2]\, S => 
        \U_ELK15_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118426);
    
    HIEFFPLA_INST_0_42322 : NAND3A
      port map(A => \U50_PATTERNS/RD_USB_ADBUS[7]\, B => 
        HIEFFPLA_NET_0_119378, C => HIEFFPLA_NET_0_119586, Y => 
        HIEFFPLA_NET_0_119572);
    
    HIEFFPLA_INST_0_60971 : MX2
      port map(A => HIEFFPLA_NET_0_117190, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_18[0]\, S => 
        HIEFFPLA_NET_0_117134, Y => HIEFFPLA_NET_0_116190);
    
    \U_ELK12_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL\ : DFN1C0
      port map(D => 
        \U_ELK12_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL_net_1\);
    
    HIEFFPLA_INST_0_56461 : AOI1D
      port map(A => HIEFFPLA_NET_0_117432, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_SEL[3]_net_1\, C
         => \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[4]_net_1\, Y
         => HIEFFPLA_NET_0_116860);
    
    HIEFFPLA_INST_0_54221 : MX2
      port map(A => HIEFFPLA_NET_0_116172, B => 
        HIEFFPLA_NET_0_116059, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_1[3]_net_1\, Y
         => HIEFFPLA_NET_0_117293);
    
    HIEFFPLA_INST_0_49178 : MX2
      port map(A => HIEFFPLA_NET_0_118179, B => 
        HIEFFPLA_NET_0_118175, S => \BIT_OS_SEL_0[1]\, Y => 
        HIEFFPLA_NET_0_118177);
    
    \U_ELK7_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]\ : DFN1C0
      port map(D => \U_ELK7_CH/U_SLAVE_1ELK/Q[7]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]_net_1\);
    
    \U50_PATTERNS/ELINK_RWA[13]/U1\ : DFN1P0
      port map(D => HIEFFPLA_NET_0_119707, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_11, Q => 
        \U50_PATTERNS/ELINK_RWA[13]\);
    
    HIEFFPLA_INST_0_54758 : NAND3A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[3]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[0]_net_1\, C => 
        HIEFFPLA_NET_0_117235, Y => HIEFFPLA_NET_0_117207);
    
    HIEFFPLA_INST_0_52722 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_25[2]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_26[2]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_3[0]\, Y => 
        HIEFFPLA_NET_0_117522);
    
    HIEFFPLA_INST_0_54652 : MX2
      port map(A => HIEFFPLA_NET_0_116185, B => 
        HIEFFPLA_NET_0_116074, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[3]_net_1\, Y => 
        HIEFFPLA_NET_0_117227);
    
    \U_EXEC_MASTER/DEL_CNT[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117788, CLK => CLK_40M_GL, CLR
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i\, Q => 
        \U_EXEC_MASTER/DEL_CNT[7]\);
    
    \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[12]\ : DFN1C0
      port map(D => \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\, 
        CLK => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\);
    
    \U0A_40M_REFCLK/\\\\BIBUF_LVDS[0]\\\\/U0/U0\ : IOPADP_BI
      port map(N2PIN => 
        \U0A_40M_REFCLK/\\\\BIBUF_LVDS[0]\\\\/U0/U2_N2P\, D => 
        \U0A_40M_REFCLK/\\\\BIBUF_LVDS[0]\\\\/U0/NET1\, E => 
        \U0A_40M_REFCLK/\\\\BIBUF_LVDS[0]\\\\/U0/NET2\, PAD => 
        BIDIR_CLK40M_P, Y => 
        \U0A_40M_REFCLK/\\\\BIBUF_LVDS[0]\\\\/U0/NET4\);
    
    HIEFFPLA_INST_0_46875 : NAND2B
      port map(A => \OP_MODE_c[1]\, B => \PATT_ELK_DAT_11[3]\, Y
         => HIEFFPLA_NET_0_118595);
    
    HIEFFPLA_INST_0_52672 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_17[3]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_18[3]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_3[0]\, Y => 
        HIEFFPLA_NET_0_117529);
    
    \U_ELK16_CH/U_ELK1_CMD_TX/START_RISE\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118374, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_0, Q => 
        \U_ELK16_CH/U_ELK1_CMD_TX/START_RISE_net_1\);
    
    \U50_PATTERNS/ELINK_ADDRA_5[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119972, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_3, Q => 
        \U50_PATTERNS/ELINK_ADDRA_5[3]\);
    
    HIEFFPLA_INST_0_42432 : AND2
      port map(A => HIEFFPLA_NET_0_119473, B => 
        \U50_PATTERNS/RD_XFER_TYPE[6]_net_1\, Y => 
        HIEFFPLA_NET_0_119535);
    
    HIEFFPLA_INST_0_41305 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_4[7]\, B => 
        HIEFFPLA_NET_0_119560, S => HIEFFPLA_NET_0_119284, Y => 
        HIEFFPLA_NET_0_119752);
    
    HIEFFPLA_INST_0_40684 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_15[2]\, B => 
        HIEFFPLA_NET_0_119575, S => HIEFFPLA_NET_0_119297, Y => 
        HIEFFPLA_NET_0_119821);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_17[4]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116201, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_7, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_17[4]\);
    
    HIEFFPLA_INST_0_49879 : MX2
      port map(A => HIEFFPLA_NET_0_118046, B => 
        HIEFFPLA_NET_0_118044, S => \BIT_OS_SEL_6[1]\, Y => 
        HIEFFPLA_NET_0_118049);
    
    HIEFFPLA_INST_0_48917 : MX2
      port map(A => HIEFFPLA_NET_0_118226, B => 
        HIEFFPLA_NET_0_118218, S => \BIT_OS_SEL_0[1]\, Y => 
        HIEFFPLA_NET_0_118224);
    
    HIEFFPLA_INST_0_51200 : MX2
      port map(A => HIEFFPLA_NET_0_117815, B => 
        HIEFFPLA_NET_0_117811, S => \BIT_OS_SEL_3[1]\, Y => 
        HIEFFPLA_NET_0_117813);
    
    \U_ELK17_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U0\ : IOPADP_BI
      port map(N2PIN => 
        \U_ELK17_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2_N2P\, D => 
        \U_ELK17_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, E => 
        \U_ELK17_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET2\, PAD => 
        ELK17_DAT_P, Y => 
        \U_ELK17_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\);
    
    HIEFFPLA_INST_0_46100 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_15[6]\, C => 
        \U50_PATTERNS/SM_BANK_SEL[4]\, Y => HIEFFPLA_NET_0_118766);
    
    HIEFFPLA_INST_0_43157 : NAND3B
      port map(A => \U50_PATTERNS/REG_STATE_0[1]_net_1\, B => 
        HIEFFPLA_NET_0_119366, C => 
        \U50_PATTERNS/REG_STATE_0[4]_net_1\, Y => 
        HIEFFPLA_NET_0_119359);
    
    \U_ELK6_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]\ : DFN1C0
      port map(D => \U_ELK6_CH/U_SLAVE_1ELK/Q[10]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]_net_1\);
    
    \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[11]\ : DFN1C0
      port map(D => 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]_net_1\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[11]_net_1\);
    
    HIEFFPLA_INST_0_45230 : NAND3C
      port map(A => HIEFFPLA_NET_0_118738, B => 
        HIEFFPLA_NET_0_118748, C => HIEFFPLA_NET_0_118757, Y => 
        HIEFFPLA_NET_0_118961);
    
    \U_ELK18_CH/U_ELK1_SERDAT_SOURCE/SERDAT[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118283, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_13, Q => 
        \U_ELK18_CH/ELK_TX_DAT[0]\);
    
    HIEFFPLA_INST_0_41125 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_2[3]\, B => 
        HIEFFPLA_NET_0_119574, S => HIEFFPLA_NET_0_119278, Y => 
        HIEFFPLA_NET_0_119772);
    
    \U50_PATTERNS/U102_PATT_ELINK_BLK/DPRT_512X9_SRAM_R0C0\ : 
        RAM4K9
      generic map(MEMORYFILE => "DPRT_512X9_SRAM_R0C0.mem")

      port map(ADDRA11 => AFLSDF_GND, ADDRA10 => AFLSDF_GND, 
        ADDRA9 => AFLSDF_GND, ADDRA8 => \GND\, ADDRA7 => 
        \U50_PATTERNS/ELINK_ADDRA_2[7]\, ADDRA6 => 
        \U50_PATTERNS/ELINK_ADDRA_2[6]\, ADDRA5 => 
        \U50_PATTERNS/ELINK_ADDRA_2[5]\, ADDRA4 => 
        \U50_PATTERNS/ELINK_ADDRA_2[4]\, ADDRA3 => 
        \U50_PATTERNS/ELINK_ADDRA_2[3]\, ADDRA2 => 
        \U50_PATTERNS/ELINK_ADDRA_2[2]\, ADDRA1 => 
        \U50_PATTERNS/ELINK_ADDRA_2[1]\, ADDRA0 => 
        \U50_PATTERNS/ELINK_ADDRA_2[0]\, ADDRB11 => AFLSDF_GND, 
        ADDRB10 => AFLSDF_GND, ADDRB9 => AFLSDF_GND, ADDRB8 => 
        \GND\, ADDRB7 => \ELKS_ADDRB[7]\, ADDRB6 => 
        \ELKS_ADDRB[6]\, ADDRB5 => \ELKS_ADDRB[5]\, ADDRB4 => 
        \ELKS_ADDRB[4]\, ADDRB3 => \ELKS_ADDRB[3]\, ADDRB2 => 
        \ELKS_ADDRB[2]\, ADDRB1 => \ELKS_ADDRB[1]\, ADDRB0 => 
        \ELKS_ADDRB[0]\, DINA8 => \GND\, DINA7 => 
        \U50_PATTERNS/ELINK_DINA_2[7]\, DINA6 => 
        \U50_PATTERNS/ELINK_DINA_2[6]\, DINA5 => 
        \U50_PATTERNS/ELINK_DINA_2[5]\, DINA4 => 
        \U50_PATTERNS/ELINK_DINA_2[4]\, DINA3 => 
        \U50_PATTERNS/ELINK_DINA_2[3]\, DINA2 => 
        \U50_PATTERNS/ELINK_DINA_2[2]\, DINA1 => 
        \U50_PATTERNS/ELINK_DINA_2[1]\, DINA0 => 
        \U50_PATTERNS/ELINK_DINA_2[0]\, DINB8 => \GND\, DINB7 => 
        \ELK_RX_SER_WORD_2[7]\, DINB6 => \ELK_RX_SER_WORD_2[6]\, 
        DINB5 => \ELK_RX_SER_WORD_2[5]\, DINB4 => 
        \ELK_RX_SER_WORD_2[4]\, DINB3 => \ELK_RX_SER_WORD_2[3]\, 
        DINB2 => \ELK_RX_SER_WORD_2[2]\, DINB1 => 
        \ELK_RX_SER_WORD_2[1]\, DINB0 => \ELK_RX_SER_WORD_2[0]\, 
        WIDTHA0 => \VCC\, WIDTHA1 => \VCC\, WIDTHB0 => \VCC\, 
        WIDTHB1 => \VCC\, PIPEA => \VCC\, PIPEB => \VCC\, WMODEA
         => \GND\, WMODEB => \GND\, BLKA => 
        \U50_PATTERNS/ELINK_BLKA[2]\, BLKB => ELKS_RAM_BLKB_EN, 
        WENA => \U50_PATTERNS/ELINK_RWA[2]\, WENB => ELKS_RWB, 
        CLKA => CLK60MHZ, CLKB => CLK_40M_GL, RESET => 
        P_USB_MASTER_EN_c_0, DOUTA8 => OPEN, DOUTA7 => 
        \U50_PATTERNS/ELINK_DOUTA_2[7]\, DOUTA6 => 
        \U50_PATTERNS/ELINK_DOUTA_2[6]\, DOUTA5 => 
        \U50_PATTERNS/ELINK_DOUTA_2[5]\, DOUTA4 => 
        \U50_PATTERNS/ELINK_DOUTA_2[4]\, DOUTA3 => 
        \U50_PATTERNS/ELINK_DOUTA_2[3]\, DOUTA2 => 
        \U50_PATTERNS/ELINK_DOUTA_2[2]\, DOUTA1 => 
        \U50_PATTERNS/ELINK_DOUTA_2[1]\, DOUTA0 => 
        \U50_PATTERNS/ELINK_DOUTA_2[0]\, DOUTB8 => OPEN, DOUTB7
         => \PATT_ELK_DAT_2[7]\, DOUTB6 => \PATT_ELK_DAT_2[6]\, 
        DOUTB5 => \PATT_ELK_DAT_2[5]\, DOUTB4 => 
        \PATT_ELK_DAT_2[4]\, DOUTB3 => \PATT_ELK_DAT_2[3]\, 
        DOUTB2 => \PATT_ELK_DAT_2[2]\, DOUTB1 => 
        \PATT_ELK_DAT_2[1]\, DOUTB0 => \PATT_ELK_DAT_2[0]\);
    
    \U50_PATTERNS/ELINK_ADDRA_15[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120045, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_6, Q => 
        \U50_PATTERNS/ELINK_ADDRA_15[2]\);
    
    \U50_PATTERNS/ELINK_ADDRA_17[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120024, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_11, Q => 
        \U50_PATTERNS/ELINK_ADDRA_17[7]\);
    
    \U_ELK8_CH/U_SLAVE_1ELK/Q[11]\ : DFN1C0
      port map(D => \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/Q[11]_net_1\);
    
    \U50_PATTERNS/ELINK_DINA_5[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119746, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_14, Q => 
        \U50_PATTERNS/ELINK_DINA_5[5]\);
    
    HIEFFPLA_INST_0_58719 : AND3
      port map(A => HIEFFPLA_NET_0_116620, B => 
        HIEFFPLA_NET_0_117204, C => HIEFFPLA_NET_0_116649, Y => 
        HIEFFPLA_NET_0_116483);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_12[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116253, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_21, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_12[2]\);
    
    HIEFFPLA_INST_0_60953 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_17[4]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_18[4]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_4[0]\, Y => 
        HIEFFPLA_NET_0_116193);
    
    \U50_PATTERNS/ELINK_ADDRA_10[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120084, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_22, Q => 
        \U50_PATTERNS/ELINK_ADDRA_10[3]\);
    
    \U50_PATTERNS/ELINKS_STRT_ADDR_T[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120098, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_21, Q => 
        \U50_PATTERNS/ELINKS_STRT_ADDR_T[5]\);
    
    HIEFFPLA_INST_0_50913 : MX2
      port map(A => \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[2]_net_1\, B
         => \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\, S => 
        \BIT_OS_SEL_3[2]\, Y => HIEFFPLA_NET_0_117864);
    
    HIEFFPLA_INST_0_47875 : NAND2B
      port map(A => \OP_MODE_c_6[1]\, B => \PATT_ELK_DAT_15[7]\, 
        Y => HIEFFPLA_NET_0_118411);
    
    HIEFFPLA_INST_0_49194 : MX2
      port map(A => \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\, B
         => \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\, S => 
        \BIT_OS_SEL[2]\, Y => HIEFFPLA_NET_0_118175);
    
    HIEFFPLA_INST_0_55312 : AND2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[6]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[3]_net_1\, Y => 
        HIEFFPLA_NET_0_117063);
    
    \U_EXEC_MASTER/MPOR_B_34\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117787, CLK => CLK_40M_GL, CLR
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_0\, Q => 
        P_MASTER_POR_B_c_34);
    
    \U_ELK18_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118285, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_0, Q => 
        \U_ELK18_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]_net_1\);
    
    HIEFFPLA_INST_0_46044 : AND3
      port map(A => \U50_PATTERNS/TFC_DOUTA[2]\, B => 
        HIEFFPLA_NET_0_118997, C => HIEFFPLA_NET_0_119365, Y => 
        HIEFFPLA_NET_0_118779);
    
    \U50_PATTERNS/ELINK_ADDRA_14[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120055, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_5, Q => 
        \U50_PATTERNS/ELINK_ADDRA_14[0]\);
    
    \U50_PATTERNS/ELINK_ADDRA_13[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120060, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_3, Q => 
        \U50_PATTERNS/ELINK_ADDRA_13[3]\);
    
    HIEFFPLA_INST_0_54079 : MX2
      port map(A => HIEFFPLA_NET_0_117351, B => 
        HIEFFPLA_NET_0_117223, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[1]_net_1\, Y
         => HIEFFPLA_NET_0_117311);
    
    HIEFFPLA_INST_0_38993 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_15[7]\, B => 
        HIEFFPLA_NET_0_119516, S => HIEFFPLA_NET_0_119297, Y => 
        HIEFFPLA_NET_0_120040);
    
    \U61_TS_WR_BUF/\\\\TRIBUFF_F_24U[0]\\\\/U0/U0\ : IOPAD_TRI_U
      port map(D => 
        \U61_TS_WR_BUF/\\\\TRIBUFF_F_24U[0]\\\\/U0/NET1\, E => 
        \U61_TS_WR_BUF/\\\\TRIBUFF_F_24U[0]\\\\/U0/NET2\, PAD => 
        USB_WR_B);
    
    HIEFFPLA_INST_0_51491 : MX2
      port map(A => HIEFFPLA_NET_0_117758, B => 
        \U_EXEC_MASTER/PRESCALE[3]\, S => HIEFFPLA_NET_0_117787, 
        Y => HIEFFPLA_NET_0_117765);
    
    HIEFFPLA_INST_0_37483 : MX2
      port map(A => \U200A_TFC/LOC_STRT_ADDR[5]\, B => 
        \TFC_STRT_ADDR[5]\, S => \U200A_TFC/GP_PG_SM_0[10]_net_1\, 
        Y => HIEFFPLA_NET_0_120277);
    
    \U50_PATTERNS/ELINK_DINA_11[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119851, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_11, Q => 
        \U50_PATTERNS/ELINK_DINA_11[4]\);
    
    HIEFFPLA_INST_0_51841 : XA1
      port map(A => \U_MASTER_DES/U13A_ADJ_160M/BITCNT[2]\, B => 
        HIEFFPLA_NET_0_117684, C => HIEFFPLA_NET_0_117631, Y => 
        HIEFFPLA_NET_0_117679);
    
    \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[9]\ : DFN1C0
      port map(D => \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\);
    
    HIEFFPLA_INST_0_56814 : AND2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_0[0]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_0[1]\, Y => 
        HIEFFPLA_NET_0_116791);
    
    \U_ELK7_CH/U_SLAVE_1ELK/Q[13]\ : DFN1C0
      port map(D => \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[13]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/Q[13]_net_1\);
    
    HIEFFPLA_INST_0_111288 : AOI1D
      port map(A => HIEFFPLA_NET_0_116740, B => 
        HIEFFPLA_NET_0_116345, C => HIEFFPLA_NET_0_117337, Y => 
        HIEFFPLA_NET_0_115842);
    
    \U_ELK14_CH/U_ELK1_CMD_TX/SER_OUT_FI\ : DFN1C0
      port map(D => 
        \U_ELK14_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_10, Q
         => \U_ELK14_CH/U_ELK1_CMD_TX/SER_OUT_FI_net_1\);
    
    HIEFFPLA_INST_0_37234 : AO1
      port map(A => HIEFFPLA_NET_0_120327, B => 
        HIEFFPLA_NET_0_120308, C => HIEFFPLA_NET_0_120300, Y => 
        HIEFFPLA_NET_0_120318);
    
    HIEFFPLA_INST_0_49065 : MX2
      port map(A => \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[0]_net_1\, 
        B => \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\, S => 
        \BIT_OS_SEL[2]\, Y => HIEFFPLA_NET_0_118204);
    
    HIEFFPLA_INST_0_38669 : MX2
      port map(A => HIEFFPLA_NET_0_119520, B => 
        \U50_PATTERNS/ELINK_ADDRA_11[3]\, S => 
        HIEFFPLA_NET_0_119280, Y => HIEFFPLA_NET_0_120076);
    
    HIEFFPLA_INST_0_62155 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_30[1]\, B => 
        HIEFFPLA_NET_0_117167, S => HIEFFPLA_NET_0_117330, Y => 
        HIEFFPLA_NET_0_116029);
    
    \U_ELK2_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]\ : DFN1C0
      port map(D => \U_ELK2_CH/U_SLAVE_1ELK/Q[6]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[13]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_115930, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_21, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[13]\);
    
    \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[9]\ : DFN1C0
      port map(D => \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\);
    
    \U200B_ELINKS/ADDR_POINTER[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120251, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_32, Q => \ELKS_ADDRB[3]\);
    
    HIEFFPLA_INST_0_113072 : AO18
      port map(A => HIEFFPLA_NET_0_115811, B => 
        \U200A_TFC/LOC_STOP_ADDR[3]\, C => \TFC_ADDRB[3]\, Y => 
        HIEFFPLA_NET_0_115818);
    
    HIEFFPLA_INST_0_54862 : NAND2A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_0[8]_net_1\, B => 
        HIEFFPLA_NET_0_115871, Y => HIEFFPLA_NET_0_117187);
    
    HIEFFPLA_INST_0_56082 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/MAX_CNT[2]\, 
        B => HIEFFPLA_NET_0_116937, S => HIEFFPLA_NET_0_117084, Y
         => HIEFFPLA_NET_0_116952);
    
    HIEFFPLA_INST_0_53779 : MX2
      port map(A => HIEFFPLA_NET_0_117230, B => 
        HIEFFPLA_NET_0_117374, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[2]_net_1\, Y
         => HIEFFPLA_NET_0_117353);
    
    HIEFFPLA_INST_0_48262 : MX2
      port map(A => HIEFFPLA_NET_0_118350, B => 
        HIEFFPLA_NET_0_118361, S => \BIT_OS_SEL_3[0]\, Y => 
        \U_ELK16_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[3]\);
    
    \U_ELK14_CH/U_SLAVE_1ELK/Q[5]\ : DFN1C0
      port map(D => \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/Q[5]_net_1\);
    
    \U50_PATTERNS/U4D_REGCROSS/LOCAL_REG_VAL[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119085, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_3, Q => \ELKS_STOP_ADDR[6]\);
    
    \U50_PATTERNS/ELINK_ADDRA_11[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120074, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_2, Q => 
        \U50_PATTERNS/ELINK_ADDRA_11[5]\);
    
    \U50_PATTERNS/ELINKS_STRT_ADDR[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120104, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_18, Q => 
        \U50_PATTERNS/ELINKS_STRT_ADDR[7]\);
    
    HIEFFPLA_INST_0_47122 : NAND2B
      port map(A => \OP_MODE_c_2[1]\, B => \PATT_ELK_DAT_12[1]\, 
        Y => HIEFFPLA_NET_0_118552);
    
    HIEFFPLA_INST_0_49612 : NAND2B
      port map(A => \OP_MODE_c_5[1]\, B => \PATT_ELK_DAT_3[1]\, Y
         => HIEFFPLA_NET_0_118102);
    
    \U200B_ELINKS/GP_PG_SM[5]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120211, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_29, Q => 
        \U200B_ELINKS/GP_PG_SM[5]_net_1\);
    
    HIEFFPLA_INST_0_63239 : NAND2B
      port map(A => \OP_MODE_c_0[1]\, B => \PATT_TFC_DAT[2]\, Y
         => \U_TFC_SERDAT_SOURCE/N_SERDAT[2]\);
    
    HIEFFPLA_INST_0_58833 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_1[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_17[1]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[4]_net_1\, Y
         => HIEFFPLA_NET_0_116470);
    
    HIEFFPLA_INST_0_40639 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_14[5]\, B => 
        HIEFFPLA_NET_0_119567, S => HIEFFPLA_NET_0_119249, Y => 
        HIEFFPLA_NET_0_119826);
    
    \U50_PATTERNS/ELINK_ADDRA_17[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120028, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_10, Q => 
        \U50_PATTERNS/ELINK_ADDRA_17[3]\);
    
    HIEFFPLA_INST_0_54333 : MX2
      port map(A => HIEFFPLA_NET_0_116445, B => 
        HIEFFPLA_NET_0_116352, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_2[3]_net_1\, Y
         => HIEFFPLA_NET_0_117279);
    
    HIEFFPLA_INST_0_37826 : AOI1B
      port map(A => \OP_MODE[4]\, B => 
        \U200B_ELINKS/GP_PG_SM[6]_net_1\, C => 
        HIEFFPLA_NET_0_120191, Y => HIEFFPLA_NET_0_120197);
    
    \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[77]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117704, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_33, Q => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[77]_net_1\);
    
    HIEFFPLA_INST_0_50867 : MX2
      port map(A => HIEFFPLA_NET_0_117866, B => 
        HIEFFPLA_NET_0_117863, S => \BIT_OS_SEL_3[1]\, Y => 
        HIEFFPLA_NET_0_117870);
    
    HIEFFPLA_INST_0_46878 : AND2A
      port map(A => \OP_MODE_c[1]\, B => \PATT_ELK_DAT_11[6]\, Y
         => HIEFFPLA_NET_0_118592);
    
    \U_ELK16_CH/U_ELK1_SERDAT_SOURCE/SERDAT[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118372, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_9, Q => 
        \U_ELK16_CH/ELK_TX_DAT[1]\);
    
    \U200B_ELINKS/GP_PG_SM[7]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120207, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_29, Q => 
        \U200B_ELINKS/GP_PG_SM[7]_net_1\);
    
    \U_ELK13_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]\ : DFN1C0
      port map(D => \U_ELK13_CH/U_SLAVE_1ELK/Q[10]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]_net_1\);
    
    \EXT_INT_REF_SEL_pad/U0/U0\ : IOPAD_IN_U
      port map(PAD => EXT_INT_REF_SEL, Y => 
        \EXT_INT_REF_SEL_pad/U0/NET1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_13[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116542, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_12, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_13[0]\);
    
    \U50_PATTERNS/ELINK_ADDRA_9[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119943, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_10, Q => 
        \U50_PATTERNS/ELINK_ADDRA_9[0]\);
    
    HIEFFPLA_INST_0_38750 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_12[4]\, B => 
        HIEFFPLA_NET_0_119519, S => HIEFFPLA_NET_0_119295, Y => 
        HIEFFPLA_NET_0_120067);
    
    HIEFFPLA_INST_0_52050 : AND2A
      port map(A => \U_MASTER_DES/U13A_ADJ_160M/BITCNT[0]\, B => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[44]_net_1\, Y => 
        HIEFFPLA_NET_0_117646);
    
    HIEFFPLA_INST_0_44754 : MX2
      port map(A => \OP_MODE_c_6[1]\, B => 
        \U50_PATTERNS/U4E_REGCROSS/SAMP_TWO[1]_net_1\, S => 
        HIEFFPLA_NET_0_119072, Y => HIEFFPLA_NET_0_119056);
    
    HIEFFPLA_INST_0_49887 : MX2
      port map(A => \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[1]_net_1\, B
         => \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\, S => 
        \BIT_OS_SEL_6[2]\, Y => HIEFFPLA_NET_0_118048);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_1[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116788, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_4, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_1[0]\);
    
    \U_ELK8_CH/ELK_IN_F\ : DFN1C0
      port map(D => \U_ELK8_CH/ELK_IN_DDR_F\, CLK => CCC_160M_ADJ, 
        CLR => DEV_RST_B_c, Q => \U_ELK8_CH/ELK_IN_F_net_1\);
    
    \U50_PATTERNS/ELINK_DINA_1[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119777, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_7, Q => 
        \U50_PATTERNS/ELINK_DINA_1[6]\);
    
    HIEFFPLA_INST_0_62257 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_31[4]\, B => 
        HIEFFPLA_NET_0_117166, S => HIEFFPLA_NET_0_117319, Y => 
        HIEFFPLA_NET_0_116016);
    
    HIEFFPLA_INST_0_56596 : AND3
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[8]_net_1\, B => 
        HIEFFPLA_NET_0_117424, C => HIEFFPLA_NET_0_117427, Y => 
        HIEFFPLA_NET_0_116831);
    
    HIEFFPLA_INST_0_53724 : NAND2B
      port map(A => HIEFFPLA_NET_0_117371, B => 
        HIEFFPLA_NET_0_117406, Y => HIEFFPLA_NET_0_117364);
    
    HIEFFPLA_INST_0_49614 : NAND2B
      port map(A => \OP_MODE_c_5[1]\, B => \PATT_ELK_DAT_3[3]\, Y
         => HIEFFPLA_NET_0_118100);
    
    HIEFFPLA_INST_0_44456 : MX2
      port map(A => \ELKS_STRT_ADDR[1]\, B => 
        \U50_PATTERNS/U4C_REGCROSS/SAMP_TWO[1]_net_1\, S => 
        HIEFFPLA_NET_0_119114, Y => HIEFFPLA_NET_0_119111);
    
    HIEFFPLA_INST_0_58727 : MX2B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_18[3]\, B => 
        HIEFFPLA_NET_0_116774, S => HIEFFPLA_NET_0_117204, Y => 
        HIEFFPLA_NET_0_116482);
    
    HIEFFPLA_INST_0_60534 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_12[2]\, B => 
        HIEFFPLA_NET_0_117131, S => HIEFFPLA_NET_0_117133, Y => 
        HIEFFPLA_NET_0_116253);
    
    HIEFFPLA_INST_0_45668 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_15[3]\, C => 
        \U50_PATTERNS/SM_BANK_SEL[4]\, Y => HIEFFPLA_NET_0_118868);
    
    HIEFFPLA_INST_0_41476 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_7[2]\, B => 
        HIEFFPLA_NET_0_119575, S => HIEFFPLA_NET_0_119289, Y => 
        HIEFFPLA_NET_0_119733);
    
    HIEFFPLA_INST_0_59871 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_31[3]\, B => 
        HIEFFPLA_NET_0_116815, S => HIEFFPLA_NET_0_117097, Y => 
        HIEFFPLA_NET_0_116340);
    
    HIEFFPLA_INST_0_47788 : MX2
      port map(A => HIEFFPLA_NET_0_118446, B => 
        HIEFFPLA_NET_0_118442, S => \BIT_OS_SEL_4[0]\, Y => 
        \U_ELK14_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[6]\);
    
    HIEFFPLA_INST_0_45171 : NAND3C
      port map(A => HIEFFPLA_NET_0_118963, B => 
        HIEFFPLA_NET_0_118759, C => HIEFFPLA_NET_0_118972, Y => 
        HIEFFPLA_NET_0_118973);
    
    \U_ELK2_CH/U_SLAVE_1ELK/Q[12]\ : DFN1C0
      port map(D => \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/Q[12]_net_1\);
    
    \U200B_ELINKS/RX_SER_WORD_2DEL[2]\ : DFN1C0
      port map(D => \U200B_ELINKS/RX_SER_WORD_1DEL[2]_net_1\, CLK
         => CLK_40M_GL, CLR => P_MASTER_POR_B_c_25, Q => 
        \U200B_ELINKS/RX_SER_WORD_2DEL[2]_net_1\);
    
    HIEFFPLA_INST_0_48776 : MX2
      port map(A => HIEFFPLA_NET_0_118267, B => 
        HIEFFPLA_NET_0_118261, S => \BIT_OS_SEL_2[0]\, Y => 
        \U_ELK18_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[5]\);
    
    HIEFFPLA_INST_0_44545 : XOR2
      port map(A => \ELKS_STRT_ADDR[7]\, B => 
        \U50_PATTERNS/U4C_REGCROSS/SAMP_TWO[7]_net_1\, Y => 
        HIEFFPLA_NET_0_119095);
    
    HIEFFPLA_INST_0_42476 : MX2
      port map(A => \U50_PATTERNS/REG_ADDR[4]\, B => 
        HIEFFPLA_NET_0_119505, S => HIEFFPLA_NET_0_119007, Y => 
        HIEFFPLA_NET_0_119529);
    
    \U_EXEC_MASTER/MPOR_B_27\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117787, CLK => CLK_40M_GL, CLR
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_0\, Q => 
        P_MASTER_POR_B_c_27);
    
    HIEFFPLA_INST_0_52109 : MX2A
      port map(A => HIEFFPLA_NET_0_117665, B => 
        HIEFFPLA_NET_0_117664, S => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[4]\, Y => 
        HIEFFPLA_NET_0_117634);
    
    \U_ELK7_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]\ : DFN1C0
      port map(D => \U_ELK7_CH/U_SLAVE_1ELK/Q[8]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]_net_1\);
    
    HIEFFPLA_INST_0_53652 : OR3B
      port map(A => HIEFFPLA_NET_0_117085, B => 
        HIEFFPLA_NET_0_116686, C => HIEFFPLA_NET_0_117325, Y => 
        HIEFFPLA_NET_0_117377);
    
    HIEFFPLA_INST_0_54063 : MX2
      port map(A => HIEFFPLA_NET_0_116452, B => 
        HIEFFPLA_NET_0_116373, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[3]_net_1\, Y
         => HIEFFPLA_NET_0_117313);
    
    HIEFFPLA_INST_0_111898 : XO1
      port map(A => \U50_PATTERNS/U4E_REGCROSS/LOCAL_REG_VAL[7]\, 
        B => \U50_PATTERNS/U4E_REGCROSS/SAMP_TWO[7]_net_1\, C => 
        HIEFFPLA_NET_0_119049, Y => HIEFFPLA_NET_0_115825);
    
    \U_ELK1_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]\ : DFN1C0
      port map(D => \U_ELK1_CH/U_SLAVE_1ELK/Q[4]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]_net_1\);
    
    HIEFFPLA_INST_0_60384 : MX2
      port map(A => HIEFFPLA_NET_0_117131, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_10[2]\, S => 
        HIEFFPLA_NET_0_117154, Y => HIEFFPLA_NET_0_116273);
    
    HIEFFPLA_INST_0_46792 : MX2
      port map(A => HIEFFPLA_NET_0_118630, B => 
        HIEFFPLA_NET_0_118627, S => \BIT_OS_SEL_0[0]\, Y => 
        \U_ELK10_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[6]\);
    
    HIEFFPLA_INST_0_47485 : MX2
      port map(A => \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[1]_net_1\, 
        B => \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\, S => 
        \BIT_OS_SEL_2[2]\, Y => HIEFFPLA_NET_0_118485);
    
    HIEFFPLA_INST_0_62794 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/TUNE_CLKPHASE[3]\, B => 
        HIEFFPLA_NET_0_115953, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[1]_net_1\, Y => 
        HIEFFPLA_NET_0_115946);
    
    HIEFFPLA_INST_0_51066 : AND2
      port map(A => \U_ELK9_CH/ELK_TX_DAT[0]\, B => 
        \U_ELK9_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_117842);
    
    \U_EXEC_MASTER/CCC_1_LOCK_STAT_0D\ : DFN1C0
      port map(D => CCC_MAIN_LOCK, CLK => CLK_40M_GL, CLR => 
        \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i\, Q => 
        \U_EXEC_MASTER/CCC_1_LOCK_STAT_0D_net_1\);
    
    HIEFFPLA_INST_0_55957 : MX2
      port map(A => HIEFFPLA_NET_0_116983, B => 
        HIEFFPLA_NET_0_117031, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[4]\, Y => 
        HIEFFPLA_NET_0_116968);
    
    HIEFFPLA_INST_0_37663 : AND3B
      port map(A => HIEFFPLA_NET_0_120148, B => 
        \U200B_ELINKS/GP_PG_SM[10]_net_1\, C => 
        HIEFFPLA_NET_0_120220, Y => HIEFFPLA_NET_0_120237);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_21[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116144, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_3, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_21[1]\);
    
    \U_ELK4_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U1\ : IOBI_ID_OD_EB
      port map(DR => \U_ELK4_CH/ELK_OUT_R_i_0\, DF => 
        \U_ELK4_CH/ELK_OUT_F_i_0\, CLR => \GND\, E => 
        \AFLSDF_INV_40\, ICLK => CCC_160M_ADJ, OCLK => 
        CCC_160M_FXD, YIN => 
        \U_ELK4_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\, DOUT => 
        \U_ELK4_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, EOUT => 
        \U_ELK4_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET2\, YR => 
        \U_ELK4_CH/U_DDR_ELK1/ELK_IN_DDR_R\, YF => 
        \U_ELK4_CH/U_DDR_ELK1/ELK_IN_DDR_F\);
    
    HIEFFPLA_INST_0_46556 : AND2
      port map(A => \ELK0_TX_DAT[1]\, B => 
        \U_ELK0_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118665);
    
    HIEFFPLA_INST_0_43693 : NAND2B
      port map(A => \U50_PATTERNS/SM_BANK_SEL[21]\, B => 
        \U50_PATTERNS/SM_BANK_SEL[9]\, Y => HIEFFPLA_NET_0_119239);
    
    \U_EXEC_MASTER/USB_MASTER_EN/TEST_SM[2]\ : DFN1P0
      port map(D => HIEFFPLA_NET_0_117751, CLK => CLK_40M_GL, PRE
         => P_MASTER_POR_B_c_24, Q => 
        \U_EXEC_MASTER/USB_MASTER_EN/TEST_SM_i_0[2]\);
    
    \U_ELK1_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U1\ : IOBI_ID_OD_EB
      port map(DR => \U_ELK1_CH/ELK_OUT_R_i_0\, DF => 
        \U_ELK1_CH/ELK_OUT_F_i_0\, CLR => \GND\, E => 
        \AFLSDF_INV_34\, ICLK => CCC_160M_ADJ, OCLK => 
        CCC_160M_FXD, YIN => 
        \U_ELK1_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\, DOUT => 
        \U_ELK1_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, EOUT => 
        \U_ELK1_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET2\, YR => 
        \U_ELK1_CH/U_DDR_ELK1/ELK_IN_DDR_R\, YF => 
        \U_ELK1_CH/U_DDR_ELK1/ELK_IN_DDR_F\);
    
    HIEFFPLA_INST_0_46909 : MX2
      port map(A => HIEFFPLA_NET_0_118577, B => 
        HIEFFPLA_NET_0_118590, S => \BIT_OS_SEL_4[1]\, Y => 
        HIEFFPLA_NET_0_118586);
    
    HIEFFPLA_INST_0_48391 : MX2
      port map(A => \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[2]_net_1\, 
        B => \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\, S => 
        \BIT_OS_SEL_0[2]\, Y => HIEFFPLA_NET_0_118318);
    
    HIEFFPLA_INST_0_48543 : MX2
      port map(A => HIEFFPLA_NET_0_118305, B => 
        HIEFFPLA_NET_0_118295, S => \BIT_OS_SEL_3[0]\, Y => 
        \U_ELK17_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[7]\);
    
    HIEFFPLA_INST_0_46364 : AO1A
      port map(A => HIEFFPLA_NET_0_118865, B => 
        \U50_PATTERNS/SM_BANK_SEL[15]\, C => 
        HIEFFPLA_NET_0_118706, Y => HIEFFPLA_NET_0_118707);
    
    HIEFFPLA_INST_0_53324 : AND3A
      port map(A => \BIT_OS_SEL_1[1]\, B => HIEFFPLA_NET_0_117423, 
        C => \BIT_OS_SEL_1[0]\, Y => HIEFFPLA_NET_0_117429);
    
    HIEFFPLA_INST_0_61760 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_9[4]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_25[4]\, S
         => \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_4[4]_net_1\, 
        Y => HIEFFPLA_NET_0_116081);
    
    \U_TFC_CMD_TX/START_RISE\ : DFN1C0
      port map(D => \U_TFC_CMD_TX/N_START_RISE\, CLK => 
        CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_TFC_CMD_TX/START_RISE_net_1\);
    
    HIEFFPLA_INST_0_57303 : XA1C
      port map(A => HIEFFPLA_NET_0_116711, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_3[4]\, C => 
        HIEFFPLA_NET_0_117179, Y => HIEFFPLA_NET_0_116703);
    
    HIEFFPLA_INST_0_46449 : AND3C
      port map(A => HIEFFPLA_NET_0_118671, B => 
        HIEFFPLA_NET_0_118675, C => HIEFFPLA_NET_0_118680, Y => 
        HIEFFPLA_NET_0_118688);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_26[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116406, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_21, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_26[0]\);
    
    \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_2S_8\ : DFN1C0
      port map(D => 
        \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_1S_net_1\, CLK
         => CLK60MHZ, CLR => P_MASTER_POR_B_c_0_0, Q => 
        P_USB_MASTER_EN_c_8);
    
    HIEFFPLA_INST_0_54630 : MX2
      port map(A => HIEFFPLA_NET_0_116181, B => 
        HIEFFPLA_NET_0_116075, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[3]_net_1\, Y => 
        HIEFFPLA_NET_0_117230);
    
    \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117040, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_16_0, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[0]\);
    
    \U_EXEC_MASTER/MPOR_SALT_B_16\ : DFI1P0
      port map(D => HIEFFPLA_NET_0_117781, CLK => CLK_40M_GL, PRE
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_2\, QN => 
        MASTER_SALT_POR_B_i_0_i_16);
    
    HIEFFPLA_INST_0_55085 : AO1
      port map(A => HIEFFPLA_NET_0_115919, B => 
        HIEFFPLA_NET_0_117108, C => HIEFFPLA_NET_0_117081, Y => 
        HIEFFPLA_NET_0_117124);
    
    HIEFFPLA_INST_0_46258 : AO1
      port map(A => HIEFFPLA_NET_0_119476, B => 
        \U50_PATTERNS/CHKSUM[3]\, C => HIEFFPLA_NET_0_118902, Y
         => HIEFFPLA_NET_0_118730);
    
    \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[6]\ : DFN1C0
      port map(D => 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\);
    
    \U50_PATTERNS/ELINK_DINA_9[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119716, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_20, Q => 
        \U50_PATTERNS/ELINK_DINA_9[3]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_5[8]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116653, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_11, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_5[8]\);
    
    \U_EXEC_MASTER/MPOR_B_21\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117787, CLK => CLK_40M_GL, CLR
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_1\, Q => 
        P_MASTER_POR_B_c_21);
    
    \U_ELK8_CH/U_ELK1_CMD_TX/SER_OUT_RI\ : DFN1C0
      port map(D => 
        \U_ELK8_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_3, Q => 
        \U_ELK8_CH/U_ELK1_CMD_TX/SER_OUT_RI_net_1\);
    
    \U_ELK1_CH/U_ELK1_CMD_TX/START_RISE\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118194, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_4, Q => 
        \U_ELK1_CH/U_ELK1_CMD_TX/START_RISE_net_1\);
    
    HIEFFPLA_INST_0_58820 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_1[3]\, B => 
        HIEFFPLA_NET_0_116468, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_1[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116472);
    
    HIEFFPLA_INST_0_41973 : AND3C
      port map(A => HIEFFPLA_NET_0_119238, B => 
        HIEFFPLA_NET_0_119270, C => 
        \U50_PATTERNS/SM_BANK_SEL[12]\, Y => 
        HIEFFPLA_NET_0_119641);
    
    HIEFFPLA_INST_0_48666 : MX2
      port map(A => HIEFFPLA_NET_0_118270, B => 
        HIEFFPLA_NET_0_118266, S => \BIT_OS_SEL_0[1]\, Y => 
        HIEFFPLA_NET_0_118269);
    
    AFLSDF_INV_28 : INV
      port map(A => DCB_SALT_SEL_c, Y => \AFLSDF_INV_28\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_14[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116235, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_2, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_14[0]\);
    
    HIEFFPLA_INST_0_42570 : NAND3A
      port map(A => HIEFFPLA_NET_0_119521, B => 
        \U50_PATTERNS/REG_ADDR[6]\, C => 
        \U50_PATTERNS/REG_ADDR[5]\, Y => HIEFFPLA_NET_0_119509);
    
    \U50_PATTERNS/WR_XFER_TYPE[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118688, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c, Q => 
        \U50_PATTERNS/WR_XFER_TYPE[1]_net_1\);
    
    \U50_PATTERNS/ELINK_ADDRA_13[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120058, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_3, Q => 
        \U50_PATTERNS/ELINK_ADDRA_13[5]\);
    
    \U_ELK7_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117926, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_11, Q => 
        \U_ELK7_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]_net_1\);
    
    HIEFFPLA_INST_0_42359 : AO1A
      port map(A => HIEFFPLA_NET_0_119581, B => 
        HIEFFPLA_NET_0_119564, C => HIEFFPLA_NET_0_119579, Y => 
        HIEFFPLA_NET_0_119557);
    
    \U50_PATTERNS/ELINK_ADDRA_8[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119950, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_8, Q => 
        \U50_PATTERNS/ELINK_ADDRA_8[1]\);
    
    HIEFFPLA_INST_0_59132 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_24[3]\, B => 
        HIEFFPLA_NET_0_116427, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_2[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116431);
    
    HIEFFPLA_INST_0_52156 : NAND2A
      port map(A => 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM[1]_net_1\, B => 
        HIEFFPLA_NET_0_117626, Y => HIEFFPLA_NET_0_117621);
    
    \U_ELK2_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U0\ : IOPADP_BI
      port map(N2PIN => 
        \U_ELK2_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2_N2P\, D => 
        \U_ELK2_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, E => 
        \U_ELK2_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET2\, PAD => 
        ELK2_DAT_P, Y => 
        \U_ELK2_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\);
    
    HIEFFPLA_INST_0_41758 : MX2
      port map(A => HIEFFPLA_NET_0_119678, B => 
        \U50_PATTERNS/ELINK_RWA[2]\, S => 
        \U50_PATTERNS/SM_BANK_SEL_0[20]\, Y => 
        HIEFFPLA_NET_0_119699);
    
    \U50_PATTERNS/ELINK_ADDRA_6[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119967, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_4, Q => 
        \U50_PATTERNS/ELINK_ADDRA_6[0]\);
    
    HIEFFPLA_INST_0_51823 : AND3
      port map(A => \U_MASTER_DES/U13A_ADJ_160M/BITCNT[1]\, B => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[3]\, C => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[4]\, Y => 
        HIEFFPLA_NET_0_117686);
    
    HIEFFPLA_INST_0_48088 : MX2
      port map(A => 
        \U_ELK16_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]_net_1\, B => 
        \U_ELK16_CH/ELK_TX_DAT[4]\, S => 
        \U_ELK16_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118380);
    
    \U_ELK12_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]\ : DFN1C0
      port map(D => \U_ELK12_CH/U_SLAVE_1ELK/Q[10]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]_net_1\);
    
    HIEFFPLA_INST_0_59889 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_3[1]\, B => 
        HIEFFPLA_NET_0_116677, S => HIEFFPLA_NET_0_117091, Y => 
        HIEFFPLA_NET_0_116338);
    
    HIEFFPLA_INST_0_47009 : MX2
      port map(A => HIEFFPLA_NET_0_118582, B => 
        HIEFFPLA_NET_0_118579, S => \BIT_OS_SEL[0]\, Y => 
        \U_ELK11_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[2]\);
    
    HIEFFPLA_INST_0_63105 : XA1C
      port map(A => HIEFFPLA_NET_0_115907, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[7]\, C => 
        HIEFFPLA_NET_0_117078, Y => HIEFFPLA_NET_0_115887);
    
    HIEFFPLA_INST_0_42093 : MX2
      port map(A => \U50_PATTERNS/OP_MODE[0]\, B => 
        \U50_PATTERNS/OP_MODE_T[0]\, S => HIEFFPLA_NET_0_119472, 
        Y => HIEFFPLA_NET_0_119617);
    
    HIEFFPLA_INST_0_62595 : MX2
      port map(A => HIEFFPLA_NET_0_117114, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_8[1]\, S => 
        HIEFFPLA_NET_0_117153, Y => HIEFFPLA_NET_0_115969);
    
    HIEFFPLA_INST_0_53860 : AND3A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[0]_net_1\, B
         => HIEFFPLA_NET_0_117235, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[3]_net_1\, Y
         => HIEFFPLA_NET_0_117341);
    
    HIEFFPLA_INST_0_37173 : AND3C
      port map(A => \U200A_TFC/GP_PG_SM[4]_net_1\, B => 
        \U200A_TFC/GP_PG_SM[5]_net_1\, C => HIEFFPLA_NET_0_120328, 
        Y => HIEFFPLA_NET_0_120334);
    
    HIEFFPLA_INST_0_60861 : AND2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[4]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_16[3]\, Y => 
        HIEFFPLA_NET_0_116207);
    
    \U_MASTER_DES/U13C_MASTER_DESER/BEST_CLKPHASE[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117450, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_10, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_CLKPHASE[2]\);
    
    \U_ELK4_CH/U_ELK1_CMD_TX/SER_OUT_FDEL\ : DFN1P0
      port map(D => \U_ELK4_CH/U_ELK1_CMD_TX/SER_OUT_FI_i\, CLK
         => CCC_160M_FXD, PRE => MASTER_SALT_POR_B_i_0_i_16, Q
         => \U_ELK4_CH/ELK_OUT_F_i_0\);
    
    HIEFFPLA_INST_0_57672 : XA1C
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_5[6]\, B => 
        HIEFFPLA_NET_0_116645, C => HIEFFPLA_NET_0_117179, Y => 
        HIEFFPLA_NET_0_116638);
    
    HIEFFPLA_INST_0_46732 : MX2
      port map(A => \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[2]_net_1\, 
        B => \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\, S => 
        \BIT_OS_SEL_5[2]\, Y => HIEFFPLA_NET_0_118621);
    
    HIEFFPLA_INST_0_40414 : MX2
      port map(A => HIEFFPLA_NET_0_119570, B => 
        \U50_PATTERNS/ELINK_DINA_11[4]\, S => 
        HIEFFPLA_NET_0_119280, Y => HIEFFPLA_NET_0_119851);
    
    HIEFFPLA_INST_0_111666 : MX2
      port map(A => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[37]_net_1\, B => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[39]_net_1\, S => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[1]\, Y => 
        HIEFFPLA_NET_0_115833);
    
    \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[71]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117708, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_33, Q => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[71]_net_1\);
    
    \U_ELK5_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118019, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_6, Q => 
        \U_ELK5_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]_net_1\);
    
    \U_ELK15_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]\ : DFN1C0
      port map(D => \U_ELK15_CH/U_SLAVE_1ELK/Q[10]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]_net_1\);
    
    \U_ELK13_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL\ : DFN1C0
      port map(D => \U_ELK13_CH/ELK_IN_R_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/RECD_SER_WORD[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_116904, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_29, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/RECD_SER_WORD[0]_net_1\);
    
    HIEFFPLA_INST_0_50760 : MX2
      port map(A => HIEFFPLA_NET_0_117906, B => 
        HIEFFPLA_NET_0_117905, S => \BIT_OS_SEL_5[0]\, Y => 
        \U_ELK7_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[4]\);
    
    HIEFFPLA_INST_0_58516 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_16[1]\, B => 
        HIEFFPLA_NET_0_116507, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_1[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116511);
    
    HIEFFPLA_INST_0_53664 : MX2
      port map(A => HIEFFPLA_NET_0_117400, B => 
        HIEFFPLA_NET_0_117232, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[1]_net_1\, Y
         => HIEFFPLA_NET_0_117375);
    
    HIEFFPLA_INST_0_53206 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_CLKPHASE[0]\, B => 
        HIEFFPLA_NET_0_117447, S => HIEFFPLA_NET_0_117111, Y => 
        HIEFFPLA_NET_0_117452);
    
    \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[3]\ : DFN1C0
      port map(D => 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[3]_net_1\);
    
    HIEFFPLA_INST_0_41062 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_1[4]\, B => 
        HIEFFPLA_NET_0_119570, S => HIEFFPLA_NET_0_119243, Y => 
        HIEFFPLA_NET_0_119779);
    
    HIEFFPLA_INST_0_44174 : MX2
      port map(A => \U50_PATTERNS/TFC_STRT_ADDR_T[0]\, B => 
        \U50_PATTERNS/RD_USB_ADBUS[0]\, S => 
        HIEFFPLA_NET_0_119491, Y => HIEFFPLA_NET_0_119164);
    
    HIEFFPLA_INST_0_42577 : XA1B
      port map(A => \U50_PATTERNS/REG_ADDR[1]\, B => 
        \U50_PATTERNS/REG_ADDR[0]\, C => HIEFFPLA_NET_0_119452, Y
         => HIEFFPLA_NET_0_119508);
    
    HIEFFPLA_INST_0_44235 : AND2
      port map(A => \U50_PATTERNS/U4A_REGCROSS/DELCNT[0]_net_1\, 
        B => \U50_PATTERNS/U4A_REGCROSS/DELCNT[1]_net_1\, Y => 
        HIEFFPLA_NET_0_119156);
    
    HIEFFPLA_INST_0_55167 : AO1E
      port map(A => HIEFFPLA_NET_0_117349, B => 
        HIEFFPLA_NET_0_117410, C => HIEFFPLA_NET_0_117085, Y => 
        HIEFFPLA_NET_0_117107);
    
    \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[0]\ : DFN1C0
      port map(D => 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[0]_net_1\);
    
    HIEFFPLA_INST_0_50609 : NAND2B
      port map(A => \OP_MODE_c_4[1]\, B => \PATT_ELK_DAT_7[2]\, Y
         => HIEFFPLA_NET_0_117921);
    
    HIEFFPLA_INST_0_50363 : AND2A
      port map(A => \OP_MODE_c_0[1]\, B => \PATT_ELK_DAT_6[5]\, Y
         => HIEFFPLA_NET_0_117963);
    
    HIEFFPLA_INST_0_61688 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_25[3]\, B => 
        HIEFFPLA_NET_0_117186, S => HIEFFPLA_NET_0_117117, Y => 
        HIEFFPLA_NET_0_116092);
    
    \U_EXEC_MASTER/MPOR_B_34_0\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117787, CLK => CLK_40M_GL, CLR
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_0\, Q => 
        P_MASTER_POR_B_c_34_0);
    
    HIEFFPLA_INST_0_54869 : NAND2B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[0]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_0[8]_net_1\, Y => 
        HIEFFPLA_NET_0_117185);
    
    HIEFFPLA_INST_0_56744 : AO1
      port map(A => HIEFFPLA_NET_0_116813, B => 
        HIEFFPLA_NET_0_117354, C => HIEFFPLA_NET_0_117371, Y => 
        HIEFFPLA_NET_0_116810);
    
    \U50_PATTERNS/ELINK_BLKA[10]/U1\ : DFN1P0
      port map(D => HIEFFPLA_NET_0_119934, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_20, Q => 
        \U50_PATTERNS/ELINK_BLKA[10]\);
    
    HIEFFPLA_INST_0_61442 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_22[4]\, B => 
        HIEFFPLA_NET_0_117166, S => HIEFFPLA_NET_0_117080, Y => 
        HIEFFPLA_NET_0_116126);
    
    \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_0[8]\ : DFN1P0
      port map(D => HIEFFPLA_NET_0_117188, CLK => CLK_40M_GL, PRE
         => P_MASTER_POR_B_c_27_1, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_0[8]_net_1\);
    
    \P_OP_MODE2_TE_pad/U0/U1\ : IOTRI_OB_EB
      port map(D => \OP_MODE_c[2]\, E => \VCC\, DOUT => 
        \P_OP_MODE2_TE_pad/U0/NET1\, EOUT => 
        \P_OP_MODE2_TE_pad/U0/NET2\);
    
    HIEFFPLA_INST_0_40252 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_0[2]\, B => 
        HIEFFPLA_NET_0_119575, S => HIEFFPLA_NET_0_119272, Y => 
        HIEFFPLA_NET_0_119869);
    
    \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[11]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_WRD_40M_FIXED[11]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_32_0, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[11]_net_1\);
    
    HIEFFPLA_INST_0_42935 : NOR2A
      port map(A => \U50_PATTERNS/REG_STATE[4]_net_1\, B => 
        HIEFFPLA_NET_0_119419, Y => HIEFFPLA_NET_0_119420);
    
    HIEFFPLA_INST_0_42760 : AO1
      port map(A => \U50_PATTERNS/REG_STATE_0[4]_net_1\, B => 
        HIEFFPLA_NET_0_119446, C => HIEFFPLA_NET_0_119599, Y => 
        HIEFFPLA_NET_0_119467);
    
    \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_1S_0\ : DFN1C0
      port map(D => 
        \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_S_net_1\, CLK => 
        CLK60MHZ, CLR => P_MASTER_POR_B_c_22_0, Q => 
        \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_1S_0_net_1\);
    
    \U_ELK5_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]\ : DFN1C0
      port map(D => \U_ELK5_CH/U_SLAVE_1ELK/Q[12]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]_net_1\);
    
    \U_ELK18_CH/U_SLAVE_1ELK/Q[8]\ : DFN1C0
      port map(D => \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/Q[8]_net_1\);
    
    HIEFFPLA_INST_0_51407 : NAND3
      port map(A => \U_EXEC_MASTER/CCC_1_LOCK_STAT_1D_net_1\, B
         => \U_EXEC_MASTER/DEL_CNT[6]\, C => 
        \U_EXEC_MASTER/DEL_CNT[4]\, Y => HIEFFPLA_NET_0_117784);
    
    HIEFFPLA_INST_0_51668 : AOI1A
      port map(A => \U_GEN_REF_CLK/GEN_40M_REFCNT[1]_net_1\, B
         => \U_GEN_REF_CLK/GEN_40M_REFCNT[2]_net_1\, C => 
        \U_GEN_REF_CLK/GEN_40M_REFCNT[0]_net_1\, Y => 
        HIEFFPLA_NET_0_117730);
    
    \U_ELK3_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]\ : DFN1C0
      port map(D => \U_ELK3_CH/U_SLAVE_1ELK/Q[14]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]_net_1\);
    
    HIEFFPLA_INST_0_51258 : MX2
      port map(A => HIEFFPLA_NET_0_117814, B => 
        HIEFFPLA_NET_0_117813, S => \BIT_OS_SEL_4[0]\, Y => 
        \U_ELK9_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[4]\);
    
    HIEFFPLA_INST_0_38534 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_0[4]\, B => 
        HIEFFPLA_NET_0_119519, S => HIEFFPLA_NET_0_119272, Y => 
        HIEFFPLA_NET_0_120091);
    
    HIEFFPLA_INST_0_38045 : AND3B
      port map(A => \U200B_ELINKS/LOC_STRT_ADDR[4]\, B => 
        HIEFFPLA_NET_0_120190, C => HIEFFPLA_NET_0_120234, Y => 
        HIEFFPLA_NET_0_120166);
    
    \U50_PATTERNS/SM_BANK_SEL[13]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119318, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_1_0, Q => 
        \U50_PATTERNS/SM_BANK_SEL[13]\);
    
    HIEFFPLA_INST_0_50029 : MX2
      port map(A => HIEFFPLA_NET_0_118036, B => 
        HIEFFPLA_NET_0_118050, S => \BIT_OS_SEL_0[0]\, Y => 
        \U_ELK4_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[6]\);
    
    \U_ELK15_CH/U_SLAVE_1ELK/Q[9]\ : DFN1C0
      port map(D => \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/Q[9]_net_1\);
    
    HIEFFPLA_INST_0_42861 : AND3
      port map(A => \U50_PATTERNS/REG_STATE[3]_net_1\, B => 
        HIEFFPLA_NET_0_119430, C => HIEFFPLA_NET_0_119380, Y => 
        HIEFFPLA_NET_0_119445);
    
    HIEFFPLA_INST_0_38018 : MX2
      port map(A => \U200B_ELINKS/LOC_STRT_ADDR[6]\, B => 
        \ELKS_STRT_ADDR[6]\, S => 
        \U200B_ELINKS/GP_PG_SM[10]_net_1\, Y => 
        HIEFFPLA_NET_0_120173);
    
    \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[3]\ : DFN1C0
      port map(D => \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\);
    
    HIEFFPLA_INST_0_60028 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_5[2]\, B => 
        HIEFFPLA_NET_0_116316, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_0[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116320);
    
    HIEFFPLA_INST_0_51338 : MX2
      port map(A => HIEFFPLA_NET_0_117777, B => 
        \U_EXEC_MASTER/DEL_CNT[1]\, S => HIEFFPLA_NET_0_117796, Y
         => HIEFFPLA_NET_0_117794);
    
    \U50_PATTERNS/REG_STATE[5]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119008, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_22_0, Q => 
        \U50_PATTERNS/REG_STATE[5]_net_1\);
    
    HIEFFPLA_INST_0_42228 : AND3B
      port map(A => HIEFFPLA_NET_0_119581, B => 
        HIEFFPLA_NET_0_119598, C => HIEFFPLA_NET_0_119564, Y => 
        HIEFFPLA_NET_0_119599);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_21[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116456, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_14, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_21[0]\);
    
    \U_ELK17_CH/U_SLAVE_1ELK/RECD_SER_WORD[1]\ : DFN1C0
      port map(D => \U_ELK17_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[1]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_17[1]\);
    
    \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[7]\ : DFN1C0
      port map(D => 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\);
    
    HIEFFPLA_INST_0_42417 : AO1A
      port map(A => HIEFFPLA_NET_0_119019, B => 
        \U50_PATTERNS/RD_USB_ADBUS[7]\, C => 
        HIEFFPLA_NET_0_119534, Y => HIEFFPLA_NET_0_119542);
    
    HIEFFPLA_INST_0_60843 : MX2
      port map(A => HIEFFPLA_NET_0_117186, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_16[3]\, S => 
        HIEFFPLA_NET_0_117142, Y => HIEFFPLA_NET_0_116212);
    
    HIEFFPLA_INST_0_55286 : AND3
      port map(A => HIEFFPLA_NET_0_117118, B => 
        HIEFFPLA_NET_0_117361, C => HIEFFPLA_NET_0_117414, Y => 
        HIEFFPLA_NET_0_117070);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_1[4]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116166, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_8, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_1[4]\);
    
    \U200B_ELINKS/LOC_STOP_ADDR[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120187, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_7, Q => 
        \U200B_ELINKS/LOC_STOP_ADDR[0]\);
    
    \U_ELK10_CH/U_SLAVE_1ELK/Q[4]\ : DFN1C0
      port map(D => \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/Q[4]_net_1\);
    
    HIEFFPLA_INST_0_44871 : AND3A
      port map(A => \U50_PATTERNS/REG_STATE_0[2]_net_1\, B => 
        HIEFFPLA_NET_0_119030, C => 
        \U50_PATTERNS/REG_STATE_0[1]_net_1\, Y => 
        HIEFFPLA_NET_0_119031);
    
    HIEFFPLA_INST_0_48870 : AND2A
      port map(A => \OP_MODE_c_6[1]\, B => \PATT_ELK_DAT_19[6]\, 
        Y => HIEFFPLA_NET_0_118232);
    
    HIEFFPLA_INST_0_44781 : XO1
      port map(A => \U50_PATTERNS/U4E_REGCROSS/SAMP_TWO[2]_net_1\, 
        B => \OP_MODE_c[2]\, C => HIEFFPLA_NET_0_119048, Y => 
        HIEFFPLA_NET_0_119051);
    
    \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[3]\ : DFN1C0
      port map(D => \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\);
    
    \U_ELK18_CH/U_SLAVE_1ELK/Q[4]\ : DFN1C0
      port map(D => \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/Q[4]_net_1\);
    
    HIEFFPLA_INST_0_62346 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_4[0]\, 
        B => HIEFFPLA_NET_0_117096, S => HIEFFPLA_NET_0_117148, Y
         => HIEFFPLA_NET_0_116000);
    
    HIEFFPLA_INST_0_43550 : AOI1D
      port map(A => HIEFFPLA_NET_0_119371, B => 
        HIEFFPLA_NET_0_119369, C => HIEFFPLA_NET_0_119296, Y => 
        HIEFFPLA_NET_0_119298);
    
    HIEFFPLA_INST_0_49740 : MX2
      port map(A => HIEFFPLA_NET_0_118084, B => 
        HIEFFPLA_NET_0_118081, S => \BIT_OS_SEL_1[0]\, Y => 
        \U_ELK3_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[1]\);
    
    \U50_PATTERNS/ELINK_ADDRA_2[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119994, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_21, Q => 
        \U50_PATTERNS/ELINK_ADDRA_2[5]\);
    
    \U50_PATTERNS/U4C_REGCROSS/LOCAL_REG_VAL[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119109, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_21, Q => \ELKS_STRT_ADDR[3]\);
    
    HIEFFPLA_INST_0_47839 : MX2
      port map(A => HIEFFPLA_NET_0_161283, B => 
        HIEFFPLA_NET_0_161282, S => HIEFFPLA_NET_0_161281, Y => 
        HIEFFPLA_NET_0_118425);
    
    HIEFFPLA_INST_0_44288 : MX2
      port map(A => \TFC_STRT_ADDR[6]\, B => 
        \U50_PATTERNS/U4A_REGCROSS/SAMP_TWO[6]_net_1\, S => 
        HIEFFPLA_NET_0_119156, Y => HIEFFPLA_NET_0_119148);
    
    \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[9]\ : DFN1C0
      port map(D => 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\);
    
    HIEFFPLA_INST_0_57790 : NAND2A
      port map(A => HIEFFPLA_NET_0_116617, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_6[4]\, Y => 
        HIEFFPLA_NET_0_116622);
    
    HIEFFPLA_INST_0_40230 : NAND3C
      port map(A => HIEFFPLA_NET_0_119389, B => 
        HIEFFPLA_NET_0_119464, C => \U50_PATTERNS/SM_BANK_SEL[8]\, 
        Y => HIEFFPLA_NET_0_119872);
    
    \U_ELK8_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117882, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_15, Q => 
        \U_ELK8_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]_net_1\);
    
    \U50_PATTERNS/ELINK_DINA_14[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119827, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_16, Q => 
        \U50_PATTERNS/ELINK_DINA_14[4]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_SEL_0[2]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_BIT_OS_VAL[2]\, CLK
         => CLK_40M_GL, CLR => P_MASTER_POR_B_c_27_1, Q => 
        \BIT_OS_SEL_0[2]\);
    
    \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[4]\ : DFN1C0
      port map(D => 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\);
    
    HIEFFPLA_INST_0_48107 : MX2
      port map(A => 
        \U_ELK16_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]_net_1\, B => 
        \U_ELK16_CH/ELK_TX_DAT[5]\, S => 
        \U_ELK16_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118376);
    
    HIEFFPLA_INST_0_44182 : MX2
      port map(A => \U50_PATTERNS/TFC_STRT_ADDR_T[1]\, B => 
        \U50_PATTERNS/RD_USB_ADBUS[1]\, S => 
        HIEFFPLA_NET_0_119491, Y => HIEFFPLA_NET_0_119163);
    
    HIEFFPLA_INST_0_38867 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_14[1]\, B => 
        HIEFFPLA_NET_0_119523, S => HIEFFPLA_NET_0_119249, Y => 
        HIEFFPLA_NET_0_120054);
    
    HIEFFPLA_INST_0_54488 : MX2
      port map(A => HIEFFPLA_NET_0_117221, B => 
        HIEFFPLA_NET_0_117384, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[1]_net_1\, Y => 
        HIEFFPLA_NET_0_117259);
    
    \U50_PATTERNS/U4B_REGCROSS/SAMP_TWO[3]\ : DFN1C0
      port map(D => \U50_PATTERNS/U4B_REGCROSS/SAMP_ONE[3]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_29, Q => 
        \U50_PATTERNS/U4B_REGCROSS/SAMP_TWO[3]_net_1\);
    
    HIEFFPLA_INST_0_53510 : MX2
      port map(A => HIEFFPLA_NET_0_117347, B => 
        HIEFFPLA_NET_0_117307, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[2]_net_1\, Y
         => HIEFFPLA_NET_0_117398);
    
    \U_ELK11_CH/U_SLAVE_1ELK/Q[7]\ : DFN1C0
      port map(D => \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/Q[7]_net_1\);
    
    \U_ELK10_CH/U_ELK1_SERDAT_SOURCE/SERDAT[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118640, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_17, Q => 
        \U_ELK10_CH/ELK_TX_DAT[3]\);
    
    HIEFFPLA_INST_0_46373 : AO1A
      port map(A => HIEFFPLA_NET_0_118861, B => 
        \U50_PATTERNS/SM_BANK_SEL[15]\, C => 
        HIEFFPLA_NET_0_118854, Y => HIEFFPLA_NET_0_118704);
    
    \U_ELK7_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]\ : DFN1C0
      port map(D => \U_ELK7_CH/U_SLAVE_1ELK/Q[10]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]_net_1\);
    
    HIEFFPLA_INST_0_48808 : MX2
      port map(A => HIEFFPLA_NET_0_118263, B => 
        HIEFFPLA_NET_0_118248, S => \BIT_OS_SEL_2[1]\, Y => 
        HIEFFPLA_NET_0_118250);
    
    \U_ELK9_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117838, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_0, Q => 
        \U_ELK9_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]_net_1\);
    
    HIEFFPLA_INST_0_48615 : AND2A
      port map(A => \OP_MODE_c_1[1]\, B => \PATT_ELK_DAT_18[0]\, 
        Y => HIEFFPLA_NET_0_118283);
    
    HIEFFPLA_INST_0_43763 : AND3B
      port map(A => HIEFFPLA_NET_0_119208, B => 
        HIEFFPLA_NET_0_119559, C => HIEFFPLA_NET_0_119564, Y => 
        HIEFFPLA_NET_0_119220);
    
    HIEFFPLA_INST_0_41907 : AOI1C
      port map(A => \U50_PATTERNS/ELINK_RWA[9]\, B => 
        HIEFFPLA_NET_0_119637, C => HIEFFPLA_NET_0_119666, Y => 
        HIEFFPLA_NET_0_119667);
    
    HIEFFPLA_INST_0_41847 : AOI1C
      port map(A => \U50_PATTERNS/ELINK_RWA[16]\, B => 
        HIEFFPLA_NET_0_119653, C => HIEFFPLA_NET_0_119683, Y => 
        HIEFFPLA_NET_0_119684);
    
    HIEFFPLA_INST_0_62726 : XNOR2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_CLKPHASE[4]\, B => 
        HIEFFPLA_NET_0_115954, Y => HIEFFPLA_NET_0_115952);
    
    HIEFFPLA_INST_0_51723 : NAND2B
      port map(A => 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM_0[4]_net_1\, B => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[78]_net_1\, Y => 
        HIEFFPLA_NET_0_117703);
    
    \U_ELK0_SERDAT_SOURCE/SERDAT[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118657, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_10, Q => \ELK0_TX_DAT[3]\);
    
    HIEFFPLA_INST_0_59930 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_3[3]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_19[3]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_5[4]_net_1\, Y
         => HIEFFPLA_NET_0_116332);
    
    \U_ELK11_CH/U_SLAVE_1ELK/Q[0]\ : DFN1C0
      port map(D => \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/Q[0]_net_1\);
    
    HIEFFPLA_INST_0_58641 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_18[1]\, B => 
        HIEFFPLA_NET_0_116490, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_2[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116494);
    
    HIEFFPLA_INST_0_46386 : AO1
      port map(A => HIEFFPLA_NET_0_119290, B => 
        \U50_PATTERNS/ELINK_DOUTA_17[2]\, C => 
        HIEFFPLA_NET_0_118843, Y => HIEFFPLA_NET_0_118701);
    
    \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[0]\ : DFN1C0
      port map(D => 
        \U_ELK7_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\);
    
    \U_ELK17_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]\ : DFN1C0
      port map(D => \U_ELK17_CH/U_SLAVE_1ELK/Q[3]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]_net_1\);
    
    HIEFFPLA_INST_0_51750 : MX2
      port map(A => \U_MASTER_DES/U13A_ADJ_160M/BITCNT[2]\, B => 
        HIEFFPLA_NET_0_117679, S => HIEFFPLA_NET_0_117630, Y => 
        HIEFFPLA_NET_0_117696);
    
    HIEFFPLA_INST_0_38768 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_12[6]\, B => 
        HIEFFPLA_NET_0_119517, S => HIEFFPLA_NET_0_119295, Y => 
        HIEFFPLA_NET_0_120065);
    
    HIEFFPLA_INST_0_43573 : NAND2B
      port map(A => \U50_PATTERNS/SM_BANK_SEL[21]\, B => 
        \U50_PATTERNS/SM_BANK_SEL[15]\, Y => 
        HIEFFPLA_NET_0_119284);
    
    HIEFFPLA_INST_0_62801 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/TUNE_CLKPHASE[4]\, B => 
        HIEFFPLA_NET_0_115952, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[1]_net_1\, Y => 
        HIEFFPLA_NET_0_115945);
    
    HIEFFPLA_INST_0_49861 : NAND2B
      port map(A => \OP_MODE_c_1[1]\, B => \PATT_ELK_DAT_4[1]\, Y
         => HIEFFPLA_NET_0_118057);
    
    HIEFFPLA_INST_0_45159 : NAND3C
      port map(A => HIEFFPLA_NET_0_118965, B => 
        HIEFFPLA_NET_0_118761, C => HIEFFPLA_NET_0_118975, Y => 
        HIEFFPLA_NET_0_118976);
    
    \U_MASTER_DES/U13A_ADJ_160M/BITCNT[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117698, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_14, Q => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[0]\);
    
    \U_ELK9_CH/U_SLAVE_1ELK/Q[5]\ : DFN1C0
      port map(D => \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/Q[5]_net_1\);
    
    \U_ELK6_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]\ : DFN1C0
      port map(D => \U_ELK6_CH/U_SLAVE_1ELK/Q[13]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]_net_1\);
    
    \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[13]\ : DFN1C0
      port map(D => \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\, 
        CLK => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[13]_net_1\);
    
    HIEFFPLA_INST_0_45911 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/SM_BANK_SEL[8]\, C => 
        \U50_PATTERNS/ELINK_DOUTA_11[7]\, Y => 
        HIEFFPLA_NET_0_118813);
    
    HIEFFPLA_INST_0_42485 : MX2
      port map(A => \U50_PATTERNS/REG_ADDR[5]\, B => 
        HIEFFPLA_NET_0_119504, S => HIEFFPLA_NET_0_119007, Y => 
        HIEFFPLA_NET_0_119528);
    
    HIEFFPLA_INST_0_40173 : AOI1C
      port map(A => \U50_PATTERNS/ELINK_BLKA[9]\, B => 
        HIEFFPLA_NET_0_119637, C => HIEFFPLA_NET_0_119879, Y => 
        HIEFFPLA_NET_0_119880);
    
    \U_ELK3_CH/U_SLAVE_1ELK/Q[10]\ : DFN1C0
      port map(D => \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/Q[10]_net_1\);
    
    \U_ELK11_CH/U_SLAVE_1ELK/Q[9]\ : DFN1C0
      port map(D => \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/Q[9]_net_1\);
    
    HIEFFPLA_INST_0_46973 : MX2
      port map(A => \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[1]_net_1\, 
        B => \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\, S => 
        \BIT_OS_SEL_4[2]\, Y => HIEFFPLA_NET_0_118577);
    
    HIEFFPLA_INST_0_40981 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_19[3]\, B => 
        HIEFFPLA_NET_0_119574, S => HIEFFPLA_NET_0_119293, Y => 
        HIEFFPLA_NET_0_119788);
    
    \U_ELK14_CH/U_SLAVE_1ELK/Q[13]\ : DFN1C0
      port map(D => \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[13]_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/Q[13]_net_1\);
    
    HIEFFPLA_INST_0_51709 : NAND2B
      port map(A => 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM[4]_net_1\, B => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[2]_net_1\, Y => 
        HIEFFPLA_NET_0_117717);
    
    HIEFFPLA_INST_0_46519 : AOI1C
      port map(A => HIEFFPLA_NET_0_119596, B => 
        HIEFFPLA_NET_0_119571, C => 
        \U50_PATTERNS/WR_XFER_TYPE[3]_net_1\, Y => 
        HIEFFPLA_NET_0_118673);
    
    HIEFFPLA_INST_0_51306 : MX2
      port map(A => \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[0]_net_1\, B
         => \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\, S => 
        \BIT_OS_SEL_2[2]\, Y => HIEFFPLA_NET_0_117799);
    
    \U_ELK16_CH/U_SLAVE_1ELK/RECD_SER_WORD[5]\ : DFN1C0
      port map(D => \U_ELK16_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[5]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_16[5]\);
    
    HIEFFPLA_INST_0_56691 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_0[6]\, B => 
        HIEFFPLA_NET_0_116794, S => HIEFFPLA_NET_0_117602, Y => 
        HIEFFPLA_NET_0_116818);
    
    HIEFFPLA_INST_0_50230 : MX2
      port map(A => HIEFFPLA_NET_0_117981, B => 
        HIEFFPLA_NET_0_117991, S => \BIT_OS_SEL_0[0]\, Y => 
        \U_ELK5_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[0]\);
    
    HIEFFPLA_INST_0_49613 : NAND2B
      port map(A => \OP_MODE_c_5[1]\, B => \PATT_ELK_DAT_3[2]\, Y
         => HIEFFPLA_NET_0_118101);
    
    HIEFFPLA_INST_0_37925 : MX2B
      port map(A => \U200B_ELINKS/N_232_li\, B => DCB_SALT_SEL_c, 
        S => \U200B_ELINKS/GP_PG_SM_0[10]_net_1\, Y => 
        HIEFFPLA_NET_0_120189);
    
    HIEFFPLA_INST_0_112131 : AO13
      port map(A => HIEFFPLA_NET_0_115820, B => 
        \U200B_ELINKS/LOC_STOP_ADDR[7]\, C => \ELKS_ADDRB[7]\, Y
         => HIEFFPLA_NET_0_120190);
    
    \U_DDR_TFC/BIBUF_LVDS_0/U0/U0\ : IOPADP_BI
      port map(N2PIN => \U_DDR_TFC/BIBUF_LVDS_0/U0/U2_N2P\, D => 
        \U_DDR_TFC/BIBUF_LVDS_0/U0/NET1\, E => 
        \U_DDR_TFC/BIBUF_LVDS_0/U0/NET2\, PAD => TFC_DAT_0P, Y
         => \U_DDR_TFC/BIBUF_LVDS_0/U0/NET4\);
    
    HIEFFPLA_INST_0_47373 : NAND2B
      port map(A => \OP_MODE_c[1]\, B => \PATT_ELK_DAT_13[3]\, Y
         => HIEFFPLA_NET_0_118505);
    
    HIEFFPLA_INST_0_43557 : AND3B
      port map(A => \U50_PATTERNS/SM_BANK_SEL_0[21]\, B => 
        \U50_PATTERNS/USB_TXE_B\, C => 
        \U50_PATTERNS/REG_STATE_0[5]_net_1\, Y => 
        HIEFFPLA_NET_0_119296);
    
    \U_MASTER_DES/U13C_MASTER_DESER/RECD_SER_WORD[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_116903, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_29, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/RECD_SER_WORD[1]_net_1\);
    
    \U_ELK11_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL\ : DFN1C0
      port map(D => 
        \U_ELK11_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL_net_1\);
    
    HIEFFPLA_INST_0_49507 : MX2
      port map(A => HIEFFPLA_NET_0_118134, B => 
        HIEFFPLA_NET_0_118130, S => \BIT_OS_SEL_1[0]\, Y => 
        \U_ELK2_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[3]\);
    
    HIEFFPLA_INST_0_38660 : MX2
      port map(A => HIEFFPLA_NET_0_119522, B => 
        \U50_PATTERNS/ELINK_ADDRA_11[2]\, S => 
        HIEFFPLA_NET_0_119280, Y => HIEFFPLA_NET_0_120077);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_6[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_115984, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_16, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_6[1]\);
    
    HIEFFPLA_INST_0_57846 : XA1C
      port map(A => HIEFFPLA_NET_0_116618, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_6[7]\, C => 
        HIEFFPLA_NET_0_117179, Y => HIEFFPLA_NET_0_116608);
    
    \U_ELK1_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118200, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_7, Q => 
        \U_ELK1_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]_net_1\);
    
    HIEFFPLA_INST_0_54830 : MX2
      port map(A => HIEFFPLA_NET_0_117281, B => 
        HIEFFPLA_NET_0_117273, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[2]_net_1\, Y => 
        HIEFFPLA_NET_0_117194);
    
    HIEFFPLA_INST_0_50045 : MX2
      port map(A => HIEFFPLA_NET_0_118024, B => 
        HIEFFPLA_NET_0_118047, S => \BIT_OS_SEL_6[1]\, Y => 
        HIEFFPLA_NET_0_118026);
    
    \U_ELK19_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118240, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_4, Q => 
        \U_ELK19_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]_net_1\);
    
    \U50_PATTERNS/ELINK_ADDRA_6[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119960, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_4, Q => 
        \U50_PATTERNS/ELINK_ADDRA_6[7]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_1[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116472, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_17_0, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_1[3]\);
    
    HIEFFPLA_INST_0_47858 : MX2
      port map(A => 
        \U_ELK15_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]_net_1\, B => 
        \U_ELK15_CH/ELK_TX_DAT[5]\, S => 
        \U_ELK15_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118421);
    
    \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_SEL_2[0]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_BIT_OS_VAL[0]\, CLK
         => CLK_40M_GL, CLR => P_MASTER_POR_B_c_27_0, Q => 
        \BIT_OS_SEL_2[0]\);
    
    HIEFFPLA_INST_0_53242 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_CLKPHASE[4]\, B => 
        HIEFFPLA_NET_0_117443, S => HIEFFPLA_NET_0_117111, Y => 
        HIEFFPLA_NET_0_117448);
    
    HIEFFPLA_INST_0_62307 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_3[4]\, 
        B => HIEFFPLA_NET_0_117100, S => HIEFFPLA_NET_0_117178, Y
         => HIEFFPLA_NET_0_116006);
    
    HIEFFPLA_INST_0_44828 : AND3
      port map(A => HIEFFPLA_NET_0_119442, B => 
        \U50_PATTERNS/REG_STATE[1]_net_1\, C => 
        HIEFFPLA_NET_0_119015, Y => HIEFFPLA_NET_0_119040);
    
    \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[8]\ : DFN1C0
      port map(D => 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\);
    
    \U_ELK17_CH/U_SLAVE_1ELK/RECD_SER_WORD[5]\ : DFN1C0
      port map(D => \U_ELK17_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[5]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_17[5]\);
    
    HIEFFPLA_INST_0_42256 : AOI1A
      port map(A => HIEFFPLA_NET_0_119601, B => 
        HIEFFPLA_NET_0_119587, C => HIEFFPLA_NET_0_119019, Y => 
        HIEFFPLA_NET_0_119588);
    
    HIEFFPLA_INST_0_55186 : AOI1D
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[6]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[8]_net_1\, C => 
        HIEFFPLA_NET_0_116708, Y => HIEFFPLA_NET_0_117101);
    
    HIEFFPLA_INST_0_61754 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_9[3]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_25[3]\, S
         => \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_3[4]_net_1\, 
        Y => HIEFFPLA_NET_0_116082);
    
    \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[14]\ : DFN1C0
      port map(D => \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\, 
        CLK => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[14]_net_1\);
    
    HIEFFPLA_INST_0_52890 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_27[2]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_28[2]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_1[0]\, Y => 
        HIEFFPLA_NET_0_117494);
    
    HIEFFPLA_INST_0_46424 : NAND2B
      port map(A => \U50_PATTERNS/WR_XFER_TYPE[0]_net_1\, B => 
        HIEFFPLA_NET_0_118692, Y => HIEFFPLA_NET_0_118693);
    
    \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[50]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117722, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_19, Q => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[50]\);
    
    HIEFFPLA_INST_0_47973 : MX2
      port map(A => HIEFFPLA_NET_0_118401, B => 
        HIEFFPLA_NET_0_118397, S => \BIT_OS_SEL_2[1]\, Y => 
        HIEFFPLA_NET_0_118396);
    
    HIEFFPLA_INST_0_37047 : AO1A
      port map(A => HIEFFPLA_NET_0_120339, B => 
        HIEFFPLA_NET_0_120325, C => HIEFFPLA_NET_0_120344, Y => 
        HIEFFPLA_NET_0_120359);
    
    \U_ELK11_CH/U_SLAVE_1ELK/Q[10]\ : DFN1C0
      port map(D => \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/Q[10]_net_1\);
    
    HIEFFPLA_INST_0_43524 : MX2
      port map(A => \U50_PATTERNS/SM_BANK_SEL[9]\, B => 
        HIEFFPLA_NET_0_119209, S => HIEFFPLA_NET_0_118691, Y => 
        HIEFFPLA_NET_0_119301);
    
    \U_ELK1_CH/U_SLAVE_1ELK/Q[6]\ : DFN1C0
      port map(D => \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/Q[6]_net_1\);
    
    HIEFFPLA_INST_0_55256 : XA1B
      port map(A => HIEFFPLA_NET_0_117225, B => 
        HIEFFPLA_NET_0_115866, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[8]_net_1\, Y => 
        HIEFFPLA_NET_0_117075);
    
    \U_ELK4_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]\ : DFN1C0
      port map(D => \U_ELK4_CH/U_SLAVE_1ELK/Q[2]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]_net_1\);
    
    \U50_PATTERNS/ELINK_ADDRA_18[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120018, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_12, Q => 
        \U50_PATTERNS/ELINK_ADDRA_18[5]\);
    
    \U0B_TX40M_REFCLK/_OUTBUF_LVDS[0]_/U0/U1\ : IOTRI_OB_EB
      port map(D => CLK_40M_BUF_RECD, E => \VCC\, DOUT => 
        \U0B_TX40M_REFCLK/\\\\OUTBUF_LVDS[0]\\\\/U0/NET1\, EOUT
         => \U0B_TX40M_REFCLK/\\\\OUTBUF_LVDS[0]\\\\/U0/NET2\);
    
    HIEFFPLA_INST_0_40504 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_12[6]\, B => 
        HIEFFPLA_NET_0_119566, S => HIEFFPLA_NET_0_119295, Y => 
        HIEFFPLA_NET_0_119841);
    
    \U_ELK7_CH/U_SLAVE_1ELK/Q[0]\ : DFN1C0
      port map(D => \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/Q[0]_net_1\);
    
    HIEFFPLA_INST_0_55050 : AO1C
      port map(A => HIEFFPLA_NET_0_117210, B => 
        HIEFFPLA_NET_0_117082, C => HIEFFPLA_NET_0_117180, Y => 
        HIEFFPLA_NET_0_117133);
    
    \U_ELK5_CH/U_SLAVE_1ELK/Q[7]\ : DFN1C0
      port map(D => \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/Q[7]_net_1\);
    
    HIEFFPLA_INST_0_62773 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/TUNE_CLKPHASE[0]\, B => 
        HIEFFPLA_NET_0_115959, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[1]_net_1\, Y => 
        HIEFFPLA_NET_0_115949);
    
    \U_ELK18_CH/U_SLAVE_1ELK/RECD_SER_WORD[3]\ : DFN1C0
      port map(D => \U_ELK18_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[3]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_18[3]\);
    
    \U_ELK16_CH/U_ELK1_SERDAT_SOURCE/SERDAT[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118373, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_9, Q => 
        \U_ELK16_CH/ELK_TX_DAT[0]\);
    
    \U200A_TFC/GP_PG_SM[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120322, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_28, Q => 
        \U200A_TFC/GP_PG_SM[0]_net_1\);
    
    HIEFFPLA_INST_0_52694 : MX2
      port map(A => HIEFFPLA_NET_0_117478, B => 
        HIEFFPLA_NET_0_117474, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[4]\, Y => 
        HIEFFPLA_NET_0_117526);
    
    HIEFFPLA_INST_0_47539 : MX2
      port map(A => HIEFFPLA_NET_0_118492, B => 
        HIEFFPLA_NET_0_118487, S => \BIT_OS_SEL_4[0]\, Y => 
        \U_ELK13_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[6]\);
    
    HIEFFPLA_INST_0_38912 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_14[6]\, B => 
        HIEFFPLA_NET_0_119517, S => HIEFFPLA_NET_0_119249, Y => 
        HIEFFPLA_NET_0_120049);
    
    \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[0]\ : DFN1C0
      port map(D => 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[0]_net_1\);
    
    HIEFFPLA_INST_0_55336 : AO1
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[4]_net_1\, B => 
        HIEFFPLA_NET_0_117027, C => HIEFFPLA_NET_0_117269, Y => 
        HIEFFPLA_NET_0_117057);
    
    HIEFFPLA_INST_0_46577 : NAND2B
      port map(A => \OP_MODE_c_4[1]\, B => \PATT_ELK_DAT_0[1]\, Y
         => HIEFFPLA_NET_0_118659);
    
    HIEFFPLA_INST_0_48152 : MX2
      port map(A => HIEFFPLA_NET_0_118362, B => 
        HIEFFPLA_NET_0_118358, S => \BIT_OS_SEL_1[1]\, Y => 
        HIEFFPLA_NET_0_118361);
    
    \U_REFCLKBUF/_BIBUF_LVDS[0]_/U0/U1\ : IOBI_IB_OB_EB
      port map(D => CLK_40M_GL, E => DCB_SALT_SEL_c, YIN => 
        \U_REFCLKBUF/\\\\BIBUF_LVDS[0]\\\\/U0/NET4\, DOUT => 
        \U_REFCLKBUF/\\\\BIBUF_LVDS[0]\\\\/U0/NET1\, EOUT => 
        \U_REFCLKBUF/\\\\BIBUF_LVDS[0]\\\\/U0/NET2\, Y => 
        EXTCLK_40MHZ_c);
    
    HIEFFPLA_INST_0_58458 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_15[1]\, B => 
        HIEFFPLA_NET_0_116677, S => HIEFFPLA_NET_0_117098, Y => 
        HIEFFPLA_NET_0_116519);
    
    \U50_PATTERNS/ELINK_ADDRA_13[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120063, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_3, Q => 
        \U50_PATTERNS/ELINK_ADDRA_13[0]\);
    
    HIEFFPLA_INST_0_50817 : AND2
      port map(A => \U_ELK8_CH/ELK_TX_DAT[0]\, B => 
        \U_ELK8_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_117887);
    
    HIEFFPLA_INST_0_38723 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_12[1]\, B => 
        HIEFFPLA_NET_0_119523, S => HIEFFPLA_NET_0_119295, Y => 
        HIEFFPLA_NET_0_120070);
    
    HIEFFPLA_INST_0_49939 : MX2
      port map(A => \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\, B
         => \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[11]_net_1\, S => 
        \BIT_OS_SEL_6[2]\, Y => HIEFFPLA_NET_0_118040);
    
    \U_ELK12_CH/U_SLAVE_1ELK/Q[6]\ : DFN1C0
      port map(D => \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/Q[6]_net_1\);
    
    \U50_PATTERNS/SM_BANK_SEL[16]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119315, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_1_0, Q => 
        \U50_PATTERNS/SM_BANK_SEL[16]\);
    
    \U50_PATTERNS/U4A_REGCROSS/LOCAL_REG_VAL[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119153, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_17, Q => \TFC_STRT_ADDR[1]\);
    
    \U_ELK8_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117883, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_15, Q => 
        \U_ELK8_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]_net_1\);
    
    \U_ELK9_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL\ : DFN1C0
      port map(D => \U_ELK9_CH/ELK_IN_R_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL_net_1\);
    
    HIEFFPLA_INST_0_57800 : NAND3B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_6[4]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_6[5]\, C => 
        HIEFFPLA_NET_0_116621, Y => HIEFFPLA_NET_0_116619);
    
    HIEFFPLA_INST_0_42611 : XA1B
      port map(A => \U50_PATTERNS/REG_ADDR[8]\, B => 
        HIEFFPLA_NET_0_119497, C => HIEFFPLA_NET_0_119452, Y => 
        HIEFFPLA_NET_0_119501);
    
    HIEFFPLA_INST_0_41620 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_9[2]\, B => 
        HIEFFPLA_NET_0_119575, S => HIEFFPLA_NET_0_119292, Y => 
        HIEFFPLA_NET_0_119717);
    
    \U_ELK13_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118517, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_1, Q => 
        \U_ELK13_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]_net_1\);
    
    \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[13]\ : DFN1C0
      port map(D => 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]_net_1\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[13]_net_1\);
    
    HIEFFPLA_INST_0_40153 : AOI1C
      port map(A => \U50_PATTERNS/ELINK_BLKA[5]\, B => 
        HIEFFPLA_NET_0_119642, C => HIEFFPLA_NET_0_119887, Y => 
        HIEFFPLA_NET_0_119888);
    
    HIEFFPLA_INST_0_56916 : AND2B
      port map(A => HIEFFPLA_NET_0_116774, B => 
        HIEFFPLA_NET_0_116708, Y => HIEFFPLA_NET_0_116776);
    
    HIEFFPLA_INST_0_46219 : AO1A
      port map(A => HIEFFPLA_NET_0_118919, B => 
        \U50_PATTERNS/SM_BANK_SEL[10]\, C => 
        HIEFFPLA_NET_0_118739, Y => HIEFFPLA_NET_0_118740);
    
    HIEFFPLA_INST_0_52600 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_9[3]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_10[3]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_1[0]\, Y => 
        HIEFFPLA_NET_0_117541);
    
    HIEFFPLA_INST_0_63089 : XA1C
      port map(A => HIEFFPLA_NET_0_115905, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[3]\, C => 
        HIEFFPLA_NET_0_117078, Y => HIEFFPLA_NET_0_115891);
    
    HIEFFPLA_INST_0_60720 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_15[1]\, B => 
        HIEFFPLA_NET_0_117167, S => HIEFFPLA_NET_0_117356, Y => 
        HIEFFPLA_NET_0_116229);
    
    HIEFFPLA_INST_0_46175 : AO1
      port map(A => HIEFFPLA_NET_0_119283, B => 
        \U50_PATTERNS/ELINK_DOUTA_13[4]\, C => 
        HIEFFPLA_NET_0_118926, Y => HIEFFPLA_NET_0_118749);
    
    HIEFFPLA_INST_0_41053 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_1[3]\, B => 
        HIEFFPLA_NET_0_119574, S => HIEFFPLA_NET_0_119243, Y => 
        HIEFFPLA_NET_0_119780);
    
    \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[7]\ : DFN1C0
      port map(D => 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\);
    
    \U_ELK15_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL\ : DFN1C0
      port map(D => 
        \U_ELK15_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL_net_1\);
    
    HIEFFPLA_INST_0_49911 : MX2
      port map(A => \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\, B
         => \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\, S => 
        \BIT_OS_SEL_6[2]\, Y => HIEFFPLA_NET_0_118044);
    
    HIEFFPLA_INST_0_47577 : MX2
      port map(A => \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\, 
        B => \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[14]_net_1\, S => 
        \BIT_OS_SEL_6[2]\, Y => HIEFFPLA_NET_0_118473);
    
    \U_ELK7_CH/U_SLAVE_1ELK/Q[12]\ : DFN1C0
      port map(D => \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/Q[12]_net_1\);
    
    \U200B_ELINKS/LOC_STRT_ADDR[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120178, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_11, Q => 
        \U200B_ELINKS/LOC_STRT_ADDR[1]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_3[4]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116006, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_11, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_3[4]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_1[5]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116783, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_4, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_1[5]\);
    
    HIEFFPLA_INST_0_39740 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_7[2]\, B => 
        HIEFFPLA_NET_0_119522, S => HIEFFPLA_NET_0_119289, Y => 
        HIEFFPLA_NET_0_119957);
    
    HIEFFPLA_INST_0_56507 : AO1
      port map(A => HIEFFPLA_NET_0_117428, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[11]_net_1\, C
         => HIEFFPLA_NET_0_116833, Y => HIEFFPLA_NET_0_116849);
    
    HIEFFPLA_INST_0_61904 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_27[0]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_28[0]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[0]\, Y => 
        HIEFFPLA_NET_0_116062);
    
    \U_MASTER_DES/U13C_MASTER_DESER/BEST_CLKPHASE[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117452, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_10, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_CLKPHASE[0]\);
    
    \U_ELK2_CH/U_SLAVE_1ELK/Q[5]\ : DFN1C0
      port map(D => \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/Q[5]_net_1\);
    
    \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[7]\ : DFN1C0
      port map(D => 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\);
    
    HIEFFPLA_INST_0_55141 : XA1B
      port map(A => HIEFFPLA_NET_0_117222, B => 
        HIEFFPLA_NET_0_117338, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[8]_net_1\, Y => 
        HIEFFPLA_NET_0_117114);
    
    \U_ELK1_CH/U_ELK1_SERDAT_SOURCE/SERDAT[5]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118188, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_11, Q => 
        \U_ELK1_CH/ELK_TX_DAT[5]\);
    
    HIEFFPLA_INST_0_48844 : AND2
      port map(A => \U_ELK19_CH/ELK_TX_DAT[1]\, B => 
        \U_ELK19_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118243);
    
    HIEFFPLA_INST_0_42837 : AND3C
      port map(A => \U50_PATTERNS/REG_STATE[5]_net_1\, B => 
        \U50_PATTERNS/REG_STATE[2]_net_1\, C => 
        HIEFFPLA_NET_0_119380, Y => HIEFFPLA_NET_0_119453);
    
    HIEFFPLA_INST_0_59758 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_14[2]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_30[2]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_3[4]_net_1\, Y
         => HIEFFPLA_NET_0_116352);
    
    HIEFFPLA_INST_0_43488 : MX2
      port map(A => \U50_PATTERNS/SM_BANK_SEL[5]\, B => 
        HIEFFPLA_NET_0_119213, S => HIEFFPLA_NET_0_118691, Y => 
        HIEFFPLA_NET_0_119305);
    
    HIEFFPLA_INST_0_49342 : AND2
      port map(A => \U_ELK2_CH/ELK_TX_DAT[1]\, B => 
        \U_ELK2_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118153);
    
    \U50_PATTERNS/ELINK_DINA_1[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119778, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_7, Q => 
        \U50_PATTERNS/ELINK_DINA_1[5]\);
    
    HIEFFPLA_INST_0_58142 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_10[3]\, B => 
        HIEFFPLA_NET_0_116815, S => HIEFFPLA_NET_0_117165, Y => 
        HIEFFPLA_NET_0_116559);
    
    \U_ELK19_CH/U_SLAVE_1ELK/RECD_SER_WORD[2]\ : DFN1C0
      port map(D => \U_ELK19_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[2]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_19[2]\);
    
    \U50_PATTERNS/ELINKS_STRT_ADDR_T[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120099, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_21, Q => 
        \U50_PATTERNS/ELINKS_STRT_ADDR_T[4]\);
    
    HIEFFPLA_INST_0_50246 : MX2
      port map(A => HIEFFPLA_NET_0_118005, B => 
        HIEFFPLA_NET_0_118002, S => \BIT_OS_SEL_0[0]\, Y => 
        \U_ELK5_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[2]\);
    
    \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_2S_13\ : DFN1C0
      port map(D => 
        \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_1S_0_net_1\, CLK
         => CLK60MHZ, CLR => \U_EXEC_MASTER/P_MASTER_POR_B_c_0\, 
        Q => P_USB_MASTER_EN_c_13);
    
    \U_ELK5_CH/U_ELK1_SERDAT_SOURCE/SERDAT[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118011, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_17, Q => 
        \U_ELK5_CH/ELK_TX_DAT[2]\);
    
    \U_TFC_CMD_TX/SER_CMD_WORD_R[3]\ : DFN1C0
      port map(D => \U_TFC_CMD_TX/N_SER_CMD_WORD_R[3]\, CLK => 
        CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_TFC_CMD_TX/SER_CMD_WORD_R[3]_net_1\);
    
    HIEFFPLA_INST_0_40720 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_15[6]\, B => 
        HIEFFPLA_NET_0_119566, S => HIEFFPLA_NET_0_119297, Y => 
        HIEFFPLA_NET_0_119817);
    
    \U50_PATTERNS/U4D_REGCROSS/SAMP_TWO[3]\ : DFN1C0
      port map(D => \U50_PATTERNS/U4D_REGCROSS/SAMP_ONE[3]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_30, Q => 
        \U50_PATTERNS/U4D_REGCROSS/SAMP_TWO[3]_net_1\);
    
    HIEFFPLA_INST_0_55251 : AO1B
      port map(A => HIEFFPLA_NET_0_117129, B => 
        HIEFFPLA_NET_0_117416, C => HIEFFPLA_NET_0_117086, Y => 
        HIEFFPLA_NET_0_117076);
    
    \U_ELK10_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U0\ : IOPADP_BI
      port map(N2PIN => 
        \U_ELK10_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2_N2P\, D => 
        \U_ELK10_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, E => 
        \U_ELK10_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET2\, PAD => 
        ELK10_DAT_P, Y => 
        \U_ELK10_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\);
    
    \U_ELK11_CH/U_ELK1_SERDAT_SOURCE/SERDAT[4]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118594, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_0, Q => 
        \U_ELK11_CH/ELK_TX_DAT[4]\);
    
    \U_ELK9_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]\ : DFN1C0
      port map(D => \U_ELK9_CH/U_SLAVE_1ELK/Q[3]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]_net_1\);
    
    HIEFFPLA_INST_0_49362 : AND2A
      port map(A => \OP_MODE_c_1[1]\, B => \PATT_ELK_DAT_2[0]\, Y
         => HIEFFPLA_NET_0_118148);
    
    \U_ELK2_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118156, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_12, Q => 
        \U_ELK2_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]_net_1\);
    
    \U_ELK11_CH/U_ELK1_CMD_TX/SER_OUT_FDEL\ : DFN1C0
      port map(D => \U_ELK11_CH/U_ELK1_CMD_TX/SER_OUT_FI_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_0, Q
         => \U_ELK11_CH/ELK_OUT_F\);
    
    HIEFFPLA_INST_0_59235 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_25[3]\, B => 
        HIEFFPLA_NET_0_116413, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_2[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116417);
    
    HIEFFPLA_INST_0_57340 : AXOI4
      port map(A => HIEFFPLA_NET_0_117085, B => 
        HIEFFPLA_NET_0_117122, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_4[0]\, Y => 
        HIEFFPLA_NET_0_116696);
    
    \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[1]\ : DFN1C0
      port map(D => 
        \U_ELK2_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\);
    
    \U_ELK15_CH/U_ELK1_CMD_TX/SER_OUT_RI\ : DFN1C0
      port map(D => 
        \U_ELK15_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_1, Q => 
        \U_ELK15_CH/U_ELK1_CMD_TX/SER_OUT_RI_net_1\);
    
    HIEFFPLA_INST_0_62640 : MX2
      port map(A => HIEFFPLA_NET_0_117114, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_9[1]\, S => 
        HIEFFPLA_NET_0_117183, Y => HIEFFPLA_NET_0_115964);
    
    HIEFFPLA_INST_0_43817 : MX2
      port map(A => HIEFFPLA_NET_0_119524, B => 
        \U50_PATTERNS/TFC_ADDRA[0]\, S => HIEFFPLA_NET_0_119294, 
        Y => HIEFFPLA_NET_0_119207);
    
    \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[2]\ : DFN1C0
      port map(D => \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\);
    
    HIEFFPLA_INST_0_42205 : MX2
      port map(A => \U50_PATTERNS/OP_MODE_T[6]\, B => 
        \U50_PATTERNS/RD_USB_ADBUS[6]\, S => 
        HIEFFPLA_NET_0_119440, Y => HIEFFPLA_NET_0_119603);
    
    HIEFFPLA_INST_0_38000 : MX2
      port map(A => \U200B_ELINKS/LOC_STRT_ADDR[3]\, B => 
        \ELKS_STRT_ADDR[3]\, S => 
        \U200B_ELINKS/GP_PG_SM_0[10]_net_1\, Y => 
        HIEFFPLA_NET_0_120176);
    
    HIEFFPLA_INST_0_50860 : AND2A
      port map(A => \OP_MODE_c_0[1]\, B => \PATT_ELK_DAT_8[4]\, Y
         => HIEFFPLA_NET_0_117874);
    
    HIEFFPLA_INST_0_52263 : AND3B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[1]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[0]_net_1\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[7]_net_1\, Y => 
        HIEFFPLA_NET_0_117598);
    
    HIEFFPLA_INST_0_40022 : MX2
      port map(A => HIEFFPLA_NET_0_119894, B => 
        \U50_PATTERNS/ELINK_BLKA[2]\, S => 
        \U50_PATTERNS/SM_BANK_SEL[20]\, Y => 
        HIEFFPLA_NET_0_119923);
    
    \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[8]\ : DFN1C0
      port map(D => \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\);
    
    \U_ELK10_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118652, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_6, Q => 
        \U_ELK10_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]_net_1\);
    
    HIEFFPLA_INST_0_53340 : MX2
      port map(A => HIEFFPLA_NET_0_117413, B => 
        HIEFFPLA_NET_0_117298, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[2]_net_1\, Y
         => HIEFFPLA_NET_0_117422);
    
    \U50_PATTERNS/U4D_REGCROSS/SAMP_ONE[2]\ : DFN1C0
      port map(D => \U50_PATTERNS/ELINKS_STOP_ADDR[2]\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_25, Q => 
        \U50_PATTERNS/U4D_REGCROSS/SAMP_ONE[2]_net_1\);
    
    HIEFFPLA_INST_0_60917 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_17[0]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_18[0]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_3[0]\, Y => 
        HIEFFPLA_NET_0_116199);
    
    HIEFFPLA_INST_0_60729 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_15[2]\, B => 
        HIEFFPLA_NET_0_117181, S => HIEFFPLA_NET_0_117356, Y => 
        HIEFFPLA_NET_0_116228);
    
    HIEFFPLA_INST_0_38813 : MX2
      port map(A => HIEFFPLA_NET_0_119520, B => 
        \U50_PATTERNS/ELINK_ADDRA_13[3]\, S => 
        HIEFFPLA_NET_0_119285, Y => HIEFFPLA_NET_0_120060);
    
    HIEFFPLA_INST_0_55914 : MX2
      port map(A => HIEFFPLA_NET_0_116152, B => 
        HIEFFPLA_NET_0_116057, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[3]\, Y => 
        HIEFFPLA_NET_0_116974);
    
    HIEFFPLA_INST_0_55858 : MX2
      port map(A => HIEFFPLA_NET_0_117015, B => 
        HIEFFPLA_NET_0_116039, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[2]\, Y => 
        HIEFFPLA_NET_0_116981);
    
    HIEFFPLA_INST_0_42089 : AO1A
      port map(A => HIEFFPLA_NET_0_119622, B => 
        \U50_PATTERNS/TFC_STOP_ADDR[7]\, C => 
        HIEFFPLA_NET_0_118670, Y => HIEFFPLA_NET_0_119618);
    
    \U_ELK4_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U0\ : IOPADP_BI
      port map(N2PIN => 
        \U_ELK4_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2_N2P\, D => 
        \U_ELK4_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, E => 
        \U_ELK4_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET2\, PAD => 
        ELK4_DAT_P, Y => 
        \U_ELK4_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\);
    
    HIEFFPLA_INST_0_62087 : MX2
      port map(A => HIEFFPLA_NET_0_116131, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_29[4]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_2[3]\, Y => 
        HIEFFPLA_NET_0_116037);
    
    HIEFFPLA_INST_0_37245 : AO1A
      port map(A => HIEFFPLA_NET_0_120297, B => 
        HIEFFPLA_NET_0_120293, C => HIEFFPLA_NET_0_120315, Y => 
        HIEFFPLA_NET_0_120316);
    
    HIEFFPLA_INST_0_54141 : MX2
      port map(A => HIEFFPLA_NET_0_116136, B => 
        HIEFFPLA_NET_0_116243, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_1[3]_net_1\, Y
         => HIEFFPLA_NET_0_117303);
    
    HIEFFPLA_INST_0_57797 : AND3C
      port map(A => HIEFFPLA_NET_0_116616, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_6[8]\, C => 
        HIEFFPLA_NET_0_116619, Y => HIEFFPLA_NET_0_116620);
    
    HIEFFPLA_INST_0_54157 : MX2
      port map(A => HIEFFPLA_NET_0_116363, B => 
        HIEFFPLA_NET_0_116557, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_1[3]_net_1\, Y
         => HIEFFPLA_NET_0_117301);
    
    HIEFFPLA_INST_0_43658 : NAND3C
      port map(A => HIEFFPLA_NET_0_119273, B => 
        HIEFFPLA_NET_0_119252, C => HIEFFPLA_NET_0_119281, Y => 
        HIEFFPLA_NET_0_119253);
    
    HIEFFPLA_INST_0_42141 : MX2
      port map(A => \U50_PATTERNS/OP_MODE[6]\, B => 
        \U50_PATTERNS/OP_MODE_T[6]\, S => HIEFFPLA_NET_0_119472, 
        Y => HIEFFPLA_NET_0_119611);
    
    \U_ELK1_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U0\ : IOPADP_BI
      port map(N2PIN => 
        \U_ELK1_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2_N2P\, D => 
        \U_ELK1_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, E => 
        \U_ELK1_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET2\, PAD => 
        ELK1_DAT_P, Y => 
        \U_ELK1_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\);
    
    \U_ELK17_CH/U_SLAVE_1ELK/Q[12]\ : DFN1C0
      port map(D => \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/Q[12]_net_1\);
    
    \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[11]\ : DFN1C0
      port map(D => 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]_net_1\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[11]_net_1\);
    
    HIEFFPLA_INST_0_43470 : MX2
      port map(A => \U50_PATTERNS/SM_BANK_SEL[3]\, B => 
        HIEFFPLA_NET_0_119215, S => HIEFFPLA_NET_0_118691, Y => 
        HIEFFPLA_NET_0_119307);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_9[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116282, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_6, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_9[3]\);
    
    HIEFFPLA_INST_0_39686 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_6[4]\, B => 
        HIEFFPLA_NET_0_119519, S => HIEFFPLA_NET_0_119258, Y => 
        HIEFFPLA_NET_0_119963);
    
    HIEFFPLA_INST_0_63221 : MX2
      port map(A => \U_TFC_CMD_TX/SER_CMD_WORD_R[0]_net_1\, B => 
        \TFC_TX_DAT[3]\, S => \U_TFC_CMD_TX/START_RISE_net_1\, Y
         => \U_TFC_CMD_TX/N_SER_CMD_WORD_R[1]\);
    
    HIEFFPLA_INST_0_62080 : MX2
      port map(A => HIEFFPLA_NET_0_116133, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_29[3]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_2[3]\, Y => 
        HIEFFPLA_NET_0_116038);
    
    \U_ELK9_CH/U_ELK1_CMD_TX/START_RISE\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117834, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_2, Q => 
        \U_ELK9_CH/U_ELK1_CMD_TX/START_RISE_net_1\);
    
    HIEFFPLA_INST_0_57880 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_7[1]\, B => 
        HIEFFPLA_NET_0_116583, S => HIEFFPLA_NET_0_117113, Y => 
        HIEFFPLA_NET_0_116602);
    
    HIEFFPLA_INST_0_49298 : MX2
      port map(A => HIEFFPLA_NET_0_118159, B => 
        HIEFFPLA_NET_0_118181, S => \BIT_OS_SEL_0[1]\, Y => 
        HIEFFPLA_NET_0_118161);
    
    HIEFFPLA_INST_0_47609 : MX2
      port map(A => 
        \U_ELK14_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]_net_1\, B => 
        \U_ELK14_CH/ELK_TX_DAT[5]\, S => 
        \U_ELK14_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118466);
    
    \U50_PATTERNS/ELINK_ADDRA_12[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120071, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_2_0, Q => 
        \U50_PATTERNS/ELINK_ADDRA_12[0]\);
    
    HIEFFPLA_INST_0_42253 : AND2
      port map(A => \U50_PATTERNS/RD_USB_ADBUS[6]\, B => 
        \U50_PATTERNS/RD_USB_ADBUS[4]\, Y => 
        HIEFFPLA_NET_0_119589);
    
    \U_ELK7_CH/U_SLAVE_1ELK/Q[5]\ : DFN1C0
      port map(D => \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/Q[5]_net_1\);
    
    HIEFFPLA_INST_0_51108 : NAND2B
      port map(A => \OP_MODE_c_3[1]\, B => \PATT_ELK_DAT_9[3]\, Y
         => HIEFFPLA_NET_0_117830);
    
    HIEFFPLA_INST_0_37208 : AND3B
      port map(A => \U200A_TFC/GP_PG_SM[9]_net_1\, B => 
        \U200A_TFC/GP_PG_SM[1]_net_1\, C => HIEFFPLA_NET_0_120333, 
        Y => HIEFFPLA_NET_0_120324);
    
    \U_ELK7_CH/U_SLAVE_1ELK/Q[6]\ : DFN1C0
      port map(D => \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/Q[6]_net_1\);
    
    \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[12]\ : DFN1C0
      port map(D => \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\);
    
    \U_ELK17_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]\ : DFN1C0
      port map(D => \U_ELK17_CH/U_SLAVE_1ELK/Q[12]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]_net_1\);
    
    \U50_PATTERNS/ELINK_DINA_0[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119864, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_5, Q => 
        \U50_PATTERNS/ELINK_DINA_0[7]\);
    
    HIEFFPLA_INST_0_59498 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_28[0]\, B => 
        HIEFFPLA_NET_0_116680, S => HIEFFPLA_NET_0_117094, Y => 
        HIEFFPLA_NET_0_116386);
    
    AFLSDF_INV_68 : INV
      port map(A => \U_ELK4_CH/U_DDR_ELK1/ELK_IN_DDR_R\, Y => 
        \AFLSDF_INV_68\);
    
    \U_ELK18_CH/U_ELK1_SERDAT_SOURCE/SERDAT[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118280, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_13, Q => 
        \U_ELK18_CH/ELK_TX_DAT[3]\);
    
    HIEFFPLA_INST_0_39551 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_4[5]\, B => 
        HIEFFPLA_NET_0_119518, S => HIEFFPLA_NET_0_119284, Y => 
        HIEFFPLA_NET_0_119978);
    
    HIEFFPLA_INST_0_47413 : MX2
      port map(A => HIEFFPLA_NET_0_118496, B => 
        HIEFFPLA_NET_0_118491, S => \BIT_OS_SEL_3[1]\, Y => 
        HIEFFPLA_NET_0_118495);
    
    HIEFFPLA_INST_0_42157 : MX2
      port map(A => \U50_PATTERNS/OP_MODE_T[0]\, B => 
        \U50_PATTERNS/RD_USB_ADBUS[0]\, S => 
        HIEFFPLA_NET_0_119440, Y => HIEFFPLA_NET_0_119609);
    
    \U_ELK16_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118381, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_14, Q => 
        \U_ELK16_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]_net_1\);
    
    HIEFFPLA_INST_0_44724 : MX2
      port map(A => \OP_MODE_c_1[1]\, B => 
        \U50_PATTERNS/U4E_REGCROSS/SAMP_TWO[1]_net_1\, S => 
        HIEFFPLA_NET_0_119072, Y => HIEFFPLA_NET_0_119061);
    
    HIEFFPLA_INST_0_43126 : NAND2A
      port map(A => \U50_PATTERNS/REG_STATE[0]_net_1\, B => 
        \U50_PATTERNS/REG_STATE[3]_net_1\, Y => 
        HIEFFPLA_NET_0_119366);
    
    HIEFFPLA_INST_0_41702 : MX2
      port map(A => HIEFFPLA_NET_0_119687, B => 
        \U50_PATTERNS/ELINK_RWA[13]\, S => 
        \U50_PATTERNS/SM_BANK_SEL_0[20]\, Y => 
        HIEFFPLA_NET_0_119707);
    
    HIEFFPLA_INST_0_46662 : MX2
      port map(A => \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\, 
        B => \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\, S => 
        \BIT_OS_SEL_5[2]\, Y => HIEFFPLA_NET_0_118631);
    
    HIEFFPLA_INST_0_46020 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/SM_BANK_SEL[3]\, C => 
        \U50_PATTERNS/ELINK_DOUTA_16[3]\, Y => 
        HIEFFPLA_NET_0_118785);
    
    HIEFFPLA_INST_0_44702 : MX2
      port map(A => \OP_MODE_c[6]\, B => 
        \U50_PATTERNS/U4E_REGCROSS/SAMP_TWO[6]_net_1\, S => 
        HIEFFPLA_NET_0_119072, Y => HIEFFPLA_NET_0_119064);
    
    \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_SEL_0[1]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_BIT_OS_VAL[1]\, CLK
         => CLK_40M_GL, CLR => P_MASTER_POR_B_c_27_0, Q => 
        \BIT_OS_SEL_0[1]\);
    
    \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[12]\ : DFN1C0
      port map(D => 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]_net_1\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[12]_net_1\);
    
    \U50_PATTERNS/REG_STATE_0[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119461, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_22_0, Q => 
        \U50_PATTERNS/REG_STATE_0[2]_net_1\);
    
    \U50_PATTERNS/ELINK_DINA_4[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119756, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_13, Q => 
        \U50_PATTERNS/ELINK_DINA_4[3]\);
    
    \U50_PATTERNS/ELINK_RWA[18]/U1\ : DFN1P0
      port map(D => HIEFFPLA_NET_0_119702, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_12, Q => 
        \U50_PATTERNS/ELINK_RWA[18]\);
    
    HIEFFPLA_INST_0_62712 : AO13
      port map(A => HIEFFPLA_NET_0_115955, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_CLKPHASE[3]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_SEQCNT[4]\, Y => 
        HIEFFPLA_NET_0_115954);
    
    HIEFFPLA_INST_0_54480 : MX2
      port map(A => HIEFFPLA_NET_0_116333, B => 
        HIEFFPLA_NET_0_116388, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[3]_net_1\, Y => 
        HIEFFPLA_NET_0_117260);
    
    \U_ELK18_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL\ : DFN1C0
      port map(D => 
        \U_ELK18_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL_net_1\);
    
    \U50_PATTERNS/ELINK_ADDRA_15[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120043, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_6, Q => 
        \U50_PATTERNS/ELINK_ADDRA_15[4]\);
    
    HIEFFPLA_INST_0_54389 : MX2
      port map(A => HIEFFPLA_NET_0_116513, B => 
        HIEFFPLA_NET_0_116296, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_2[3]_net_1\, Y
         => HIEFFPLA_NET_0_117272);
    
    HIEFFPLA_INST_0_50114 : AND2A
      port map(A => \OP_MODE_c_4[1]\, B => \PATT_ELK_DAT_5[5]\, Y
         => HIEFFPLA_NET_0_118008);
    
    HIEFFPLA_INST_0_42858 : AND3B
      port map(A => HIEFFPLA_NET_0_119380, B => 
        \U50_PATTERNS/REG_STATE[3]_net_1\, C => 
        HIEFFPLA_NET_0_119429, Y => HIEFFPLA_NET_0_119446);
    
    HIEFFPLA_INST_0_60317 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_9[3]\, B => 
        HIEFFPLA_NET_0_116276, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_0[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116282);
    
    HIEFFPLA_INST_0_42083 : AO1A
      port map(A => HIEFFPLA_NET_0_119622, B => 
        \U50_PATTERNS/TFC_STOP_ADDR[5]\, C => 
        HIEFFPLA_NET_0_118670, Y => HIEFFPLA_NET_0_119619);
    
    HIEFFPLA_INST_0_39938 : MX2
      port map(A => HIEFFPLA_NET_0_119915, B => 
        \U50_PATTERNS/ELINK_BLKA[0]\, S => 
        \U50_PATTERNS/SM_BANK_SEL_0[20]\, Y => 
        HIEFFPLA_NET_0_119935);
    
    \U_ELK14_CH/U_ELK1_CMD_TX/SER_OUT_FDEL\ : DFN1C0
      port map(D => \U_ELK14_CH/U_ELK1_CMD_TX/SER_OUT_FI_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_15, Q
         => \U_ELK14_CH/ELK_OUT_F\);
    
    HIEFFPLA_INST_0_58387 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_14[0]\, B => 
        HIEFFPLA_NET_0_116680, S => HIEFFPLA_NET_0_117159, Y => 
        HIEFFPLA_NET_0_116528);
    
    HIEFFPLA_INST_0_48140 : MX2
      port map(A => \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[3]_net_1\, 
        B => \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\, S => 
        \BIT_OS_SEL_1[2]\, Y => HIEFFPLA_NET_0_118363);
    
    HIEFFPLA_INST_0_50074 : MX2
      port map(A => 
        \U_ELK5_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]_net_1\, B => 
        \U_ELK5_CH/ELK_TX_DAT[2]\, S => 
        \U_ELK5_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118021);
    
    HIEFFPLA_INST_0_161272 : DFN1C0
      port map(D => 
        \U_ELK15_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_9, Q => 
        HIEFFPLA_NET_0_161283);
    
    \U_ELK13_CH/U_ELK1_SERDAT_SOURCE/SERDAT[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118506, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_4, Q => 
        \U_ELK13_CH/ELK_TX_DAT[2]\);
    
    HIEFFPLA_INST_0_56013 : MX2
      port map(A => HIEFFPLA_NET_0_117021, B => 
        HIEFFPLA_NET_0_117011, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[2]\, Y => 
        HIEFFPLA_NET_0_116961);
    
    HIEFFPLA_INST_0_54971 : OA1A
      port map(A => HIEFFPLA_NET_0_117242, B => 
        HIEFFPLA_NET_0_117245, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_3[6]_net_1\, Y => 
        HIEFFPLA_NET_0_117152);
    
    HIEFFPLA_INST_0_53260 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_SEQCNT[0]\, B => 
        HIEFFPLA_NET_0_117437, S => HIEFFPLA_NET_0_117062, Y => 
        HIEFFPLA_NET_0_117442);
    
    \U_ELK10_CH/U_ELK1_SERDAT_SOURCE/SERDAT[6]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118637, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_17, Q => 
        \U_ELK10_CH/ELK_TX_DAT[6]\);
    
    \U50_PATTERNS/ELINK_DINA_0[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119871, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_5, Q => 
        \U50_PATTERNS/ELINK_DINA_0[0]\);
    
    HIEFFPLA_INST_0_55536 : MX2
      port map(A => HIEFFPLA_NET_0_116165, B => 
        HIEFFPLA_NET_0_116270, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[3]\, Y => 
        HIEFFPLA_NET_0_117024);
    
    HIEFFPLA_INST_0_41944 : NAND2
      port map(A => HIEFFPLA_NET_0_119389, B => 
        \U50_PATTERNS/SM_BANK_SEL[1]\, Y => HIEFFPLA_NET_0_119651);
    
    \P_USB_RXF_B_pad/U0/U0\ : IOPAD_IN_U
      port map(PAD => P_USB_RXF_B, Y => \P_USB_RXF_B_pad/U0/NET1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/Q[4]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[4]_net_1\, CLK => 
        CCC_160M_FXD, CLR => P_MASTER_POR_B_c_34, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/Q[4]_net_1\);
    
    HIEFFPLA_INST_0_62197 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_14[0]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_30[0]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[4]_net_1\, Y => 
        HIEFFPLA_NET_0_116024);
    
    HIEFFPLA_INST_0_46190 : AO1
      port map(A => HIEFFPLA_NET_0_119254, B => 
        \U50_PATTERNS/ELINK_DOUTA_6[7]\, C => 
        HIEFFPLA_NET_0_118923, Y => HIEFFPLA_NET_0_118746);
    
    HIEFFPLA_INST_0_41503 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_7[5]\, B => 
        HIEFFPLA_NET_0_119567, S => HIEFFPLA_NET_0_119289, Y => 
        HIEFFPLA_NET_0_119730);
    
    HIEFFPLA_INST_0_42317 : AND3A
      port map(A => HIEFFPLA_NET_0_119572, B => 
        HIEFFPLA_NET_0_119430, C => HIEFFPLA_NET_0_119557, Y => 
        HIEFFPLA_NET_0_119573);
    
    \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_SEL_7[2]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_BIT_OS_VAL[2]\, CLK
         => CLK_40M_GL, CLR => P_MASTER_POR_B_c_27_0, Q => 
        \BIT_OS_SEL_7[2]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_115937, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_24_0, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[3]_net_1\);
    
    HIEFFPLA_INST_0_39776 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_7[6]\, B => 
        HIEFFPLA_NET_0_119517, S => HIEFFPLA_NET_0_119289, Y => 
        HIEFFPLA_NET_0_119953);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_11[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116264, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_20, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_11[1]\);
    
    HIEFFPLA_INST_0_53395 : AND2A
      port map(A => HIEFFPLA_NET_0_117390, B => 
        HIEFFPLA_NET_0_117325, Y => HIEFFPLA_NET_0_117415);
    
    HIEFFPLA_INST_0_37525 : NAND3C
      port map(A => \U200A_TFC/RX_SER_WORD_3DEL_i_0[1]\, B => 
        \U200A_TFC/RX_SER_WORD_3DEL[0]_net_1\, C => 
        HIEFFPLA_NET_0_120269, Y => HIEFFPLA_NET_0_120267);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_27[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116067, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_13, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_27[3]\);
    
    HIEFFPLA_INST_0_47953 : MX2
      port map(A => HIEFFPLA_NET_0_118409, B => 
        HIEFFPLA_NET_0_118406, S => \BIT_OS_SEL_2[1]\, Y => 
        HIEFFPLA_NET_0_118399);
    
    HIEFFPLA_INST_0_45478 : AO1
      port map(A => HIEFFPLA_NET_0_119288, B => 
        \U50_PATTERNS/ELINK_DOUTA_16[7]\, C => 
        HIEFFPLA_NET_0_118813, Y => HIEFFPLA_NET_0_118906);
    
    HIEFFPLA_INST_0_41098 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_2[0]\, B => 
        HIEFFPLA_NET_0_119578, S => HIEFFPLA_NET_0_119278, Y => 
        HIEFFPLA_NET_0_119775);
    
    HIEFFPLA_INST_0_45732 : AO1
      port map(A => HIEFFPLA_NET_0_119236, B => 
        \U50_PATTERNS/ELINK_DOUTA_0[5]\, C => 
        HIEFFPLA_NET_0_118784, Y => HIEFFPLA_NET_0_118856);
    
    \U_EXEC_MASTER/USB_MASTER_EN/TEST_SM[4]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117749, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_24, Q => 
        \U_EXEC_MASTER/USB_MASTER_EN/TEST_SM[4]_net_1\);
    
    \U50_PATTERNS/ELINK_DINA_0[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119870, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_5, Q => 
        \U50_PATTERNS/ELINK_DINA_0[1]\);
    
    HIEFFPLA_INST_0_53549 : MX2
      port map(A => HIEFFPLA_NET_0_117401, B => 
        HIEFFPLA_NET_0_117372, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[0]_net_1\, Y
         => HIEFFPLA_NET_0_117390);
    
    HIEFFPLA_INST_0_45328 : AO1
      port map(A => HIEFFPLA_NET_0_119246, B => 
        \U50_PATTERNS/ELINK_DOUTA_3[6]\, C => 
        HIEFFPLA_NET_0_118822, Y => HIEFFPLA_NET_0_118939);
    
    \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[5]\ : DFN1C0
      port map(D => 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\);
    
    HIEFFPLA_INST_0_52195 : AND3A
      port map(A => HIEFFPLA_NET_0_117688, B => 
        HIEFFPLA_NET_0_117612, C => HIEFFPLA_NET_0_117681, Y => 
        HIEFFPLA_NET_0_117613);
    
    HIEFFPLA_INST_0_113942 : AO18
      port map(A => HIEFFPLA_NET_0_115808, B => 
        \U200B_ELINKS/LOC_STOP_ADDR[5]\, C => \ELKS_ADDRB[5]\, Y
         => HIEFFPLA_NET_0_115812);
    
    HIEFFPLA_INST_0_49361 : AND2
      port map(A => CLK_40M_GL, B => 
        \U_ELK2_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0_net_1\, Y => 
        HIEFFPLA_NET_0_118149);
    
    HIEFFPLA_INST_0_43805 : AND3A
      port map(A => \U50_PATTERNS/RD_USB_ADBUS[2]\, B => 
        HIEFFPLA_NET_0_119591, C => 
        \U50_PATTERNS/RD_USB_ADBUS[3]\, Y => 
        HIEFFPLA_NET_0_119210);
    
    HIEFFPLA_INST_0_60010 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_5[0]\, B => 
        HIEFFPLA_NET_0_116680, S => HIEFFPLA_NET_0_117156, Y => 
        HIEFFPLA_NET_0_116322);
    
    HIEFFPLA_INST_0_39578 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_5[0]\, B => 
        HIEFFPLA_NET_0_119524, S => HIEFFPLA_NET_0_119251, Y => 
        HIEFFPLA_NET_0_119975);
    
    \U_ELK7_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]\ : DFN1C0
      port map(D => \U_ELK7_CH/U_SLAVE_1ELK/Q[13]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]_net_1\);
    
    \U_ELK17_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]\ : DFN1C0
      port map(D => \U_ELK17_CH/U_SLAVE_1ELK/Q[6]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]_net_1\);
    
    \U50_PATTERNS/ELINK_BLKA[19]/U1\ : DFN1P0
      port map(D => HIEFFPLA_NET_0_119925, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_20, Q => 
        \U50_PATTERNS/ELINK_BLKA[19]\);
    
    HIEFFPLA_INST_0_52800 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_11[3]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_12[3]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_1[0]\, Y => 
        HIEFFPLA_NET_0_117509);
    
    HIEFFPLA_INST_0_51049 : MX2
      port map(A => HIEFFPLA_NET_0_117856, B => 
        HIEFFPLA_NET_0_117843, S => \BIT_OS_SEL_5[1]\, Y => 
        HIEFFPLA_NET_0_117845);
    
    \U_ELK12_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118562, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_15, Q => 
        \U_ELK12_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]_net_1\);
    
    HIEFFPLA_INST_0_49780 : MX2
      port map(A => HIEFFPLA_NET_0_118093, B => 
        HIEFFPLA_NET_0_118090, S => \BIT_OS_SEL_1[0]\, Y => 
        \U_ELK3_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[6]\);
    
    HIEFFPLA_INST_0_50610 : NAND2B
      port map(A => \OP_MODE_c_4[1]\, B => \PATT_ELK_DAT_7[3]\, Y
         => HIEFFPLA_NET_0_117920);
    
    \U_ELK7_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]\ : DFN1C0
      port map(D => \U_ELK7_CH/U_SLAVE_1ELK/Q[4]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]_net_1\);
    
    \U_ELK4_CH/U_SLAVE_1ELK/Q[6]\ : DFN1C0
      port map(D => \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/Q[6]_net_1\);
    
    HIEFFPLA_INST_0_41566 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_8[4]\, B => 
        HIEFFPLA_NET_0_119570, S => HIEFFPLA_NET_0_119291, Y => 
        HIEFFPLA_NET_0_119723);
    
    HIEFFPLA_INST_0_38314 : MX2
      port map(A => \U50_PATTERNS/ELINKS_STOP_ADDR_T[1]\, B => 
        \U50_PATTERNS/RD_USB_ADBUS[1]\, S => 
        HIEFFPLA_NET_0_119413, Y => HIEFFPLA_NET_0_120118);
    
    \U_MASTER_DES/U13A_ADJ_160M/BITCNT[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117696, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_14, Q => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[2]\);
    
    \U_ELK8_CH/ELK_IN_R\ : DFN1C0
      port map(D => \U_ELK8_CH/ELK_IN_DDR_R\, CLK => CCC_160M_ADJ, 
        CLR => DEV_RST_B_c, Q => \U_ELK8_CH/ELK_IN_R_net_1\);
    
    HIEFFPLA_INST_0_39074 : MX2
      port map(A => HIEFFPLA_NET_0_119524, B => 
        \U50_PATTERNS/ELINK_ADDRA_17[0]\, S => 
        HIEFFPLA_NET_0_119260, Y => HIEFFPLA_NET_0_120031);
    
    \U50_PATTERNS/ELINK_ADDRA_16[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120032, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_9, Q => 
        \U50_PATTERNS/ELINK_ADDRA_16[7]\);
    
    HIEFFPLA_INST_0_39632 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_5[6]\, B => 
        HIEFFPLA_NET_0_119517, S => HIEFFPLA_NET_0_119251, Y => 
        HIEFFPLA_NET_0_119969);
    
    \U50_PATTERNS/U4D_REGCROSS/LOCAL_REG_VAL[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119088, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_3, Q => \ELKS_STOP_ADDR[3]\);
    
    HIEFFPLA_INST_0_52758 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_3[0]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_4[0]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[0]\, Y => 
        HIEFFPLA_NET_0_117516);
    
    HIEFFPLA_INST_0_38624 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_10[6]\, B => 
        HIEFFPLA_NET_0_119517, S => HIEFFPLA_NET_0_119239, Y => 
        HIEFFPLA_NET_0_120081);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_7[7]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116596, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_14, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_7[7]\);
    
    \U_ELK10_CH/ELK_IN_R\ : DFN1C0
      port map(D => \U_ELK10_CH/ELK_IN_DDR_R\, CLK => 
        CCC_160M_ADJ, CLR => DEV_RST_B_c, Q => 
        \U_ELK10_CH/ELK_IN_R_net_1\);
    
    HIEFFPLA_INST_0_44650 : XOR2
      port map(A => \U50_PATTERNS/U4D_REGCROSS/DELCNT[0]_net_1\, 
        B => \U50_PATTERNS/U4D_REGCROSS/DELCNT[1]_net_1\, Y => 
        HIEFFPLA_NET_0_119073);
    
    HIEFFPLA_INST_0_54411 : AND3
      port map(A => HIEFFPLA_NET_0_117063, B => 
        HIEFFPLA_NET_0_117386, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_4[4]_net_1\, Y
         => HIEFFPLA_NET_0_117269);
    
    \U200A_TFC/LOC_STOP_ADDR[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120283, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_1, Q => \U200A_TFC/LOC_STOP_ADDR[7]\);
    
    HIEFFPLA_INST_0_38186 : MX2
      port map(A => \U50_PATTERNS/CHKSUM[4]\, B => 
        HIEFFPLA_NET_0_120131, S => HIEFFPLA_NET_0_119470, Y => 
        HIEFFPLA_NET_0_120139);
    
    \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[3]\ : DFN1C0
      port map(D => \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\);
    
    HIEFFPLA_INST_0_59221 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_25[1]\, B => 
        HIEFFPLA_NET_0_116415, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_2[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116419);
    
    \U_ELK12_CH/ELK_IN_R\ : DFN1C0
      port map(D => \U_ELK12_CH/ELK_IN_DDR_R\, CLK => 
        CCC_160M_ADJ, CLR => DEV_RST_B_c, Q => 
        \U_ELK12_CH/ELK_IN_R_net_1\);
    
    HIEFFPLA_INST_0_39767 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_7[5]\, B => 
        HIEFFPLA_NET_0_119518, S => HIEFFPLA_NET_0_119289, Y => 
        HIEFFPLA_NET_0_119954);
    
    HIEFFPLA_INST_0_38290 : MX2
      port map(A => \U50_PATTERNS/ELINKS_STOP_ADDR[6]\, B => 
        \U50_PATTERNS/ELINKS_STOP_ADDR_T[6]\, S => 
        HIEFFPLA_NET_0_119472, Y => HIEFFPLA_NET_0_120121);
    
    \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[2]\ : DFN1C0
      port map(D => \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\);
    
    HIEFFPLA_INST_0_63045 : NAND3
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[0]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[1]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[2]\, Y => 
        HIEFFPLA_NET_0_115905);
    
    HIEFFPLA_INST_0_51712 : NAND2B
      port map(A => 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM[4]_net_1\, B => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[37]_net_1\, Y => 
        HIEFFPLA_NET_0_117714);
    
    \U_ELK11_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]\ : DFN1C0
      port map(D => \U_ELK11_CH/U_SLAVE_1ELK/Q[10]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]_net_1\);
    
    \U_ELK17_CH/U_SLAVE_1ELK/RECD_SER_WORD[3]\ : DFN1C0
      port map(D => \U_ELK17_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[3]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_17[3]\);
    
    \U_ELK17_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]\ : DFN1C0
      port map(D => \U_ELK17_CH/U_SLAVE_1ELK/Q[14]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]_net_1\);
    
    \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[9]\ : DFN1C0
      port map(D => \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\);
    
    \U50_PATTERNS/ELINKS_STRT_ADDR[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120105, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_17, Q => 
        \U50_PATTERNS/ELINKS_STRT_ADDR[6]\);
    
    HIEFFPLA_INST_0_45224 : NAND3C
      port map(A => HIEFFPLA_NET_0_118740, B => 
        HIEFFPLA_NET_0_118749, C => HIEFFPLA_NET_0_118758, Y => 
        HIEFFPLA_NET_0_118962);
    
    HIEFFPLA_INST_0_58957 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_21[2]\, B => 
        HIEFFPLA_NET_0_116687, S => HIEFFPLA_NET_0_117093, Y => 
        HIEFFPLA_NET_0_116454);
    
    HIEFFPLA_INST_0_46130 : AO1
      port map(A => HIEFFPLA_NET_0_119244, B => 
        \U50_PATTERNS/ELINK_DOUTA_2[3]\, C => 
        HIEFFPLA_NET_0_118934, Y => HIEFFPLA_NET_0_118759);
    
    HIEFFPLA_INST_0_43735 : AND3A
      port map(A => \U50_PATTERNS/RD_USB_ADBUS[2]\, B => 
        HIEFFPLA_NET_0_119593, C => 
        \U50_PATTERNS/RD_USB_ADBUS[3]\, Y => 
        HIEFFPLA_NET_0_119227);
    
    HIEFFPLA_INST_0_42992 : AO1A
      port map(A => HIEFFPLA_NET_0_119394, B => 
        HIEFFPLA_NET_0_119448, C => HIEFFPLA_NET_0_119412, Y => 
        HIEFFPLA_NET_0_119407);
    
    \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[13]\ : DFN1C0
      port map(D => \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[13]_net_1\);
    
    \U_ELK12_CH/U_ELK1_SERDAT_SOURCE/SERDAT[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118551, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_2, Q => 
        \U_ELK12_CH/ELK_TX_DAT[2]\);
    
    HIEFFPLA_INST_0_44230 : MX2
      port map(A => \U50_PATTERNS/TFC_STRT_ADDR_T[7]\, B => 
        \U50_PATTERNS/RD_USB_ADBUS[7]\, S => 
        HIEFFPLA_NET_0_119491, Y => HIEFFPLA_NET_0_119157);
    
    HIEFFPLA_INST_0_42986 : NAND3C
      port map(A => HIEFFPLA_NET_0_119416, B => 
        HIEFFPLA_NET_0_119011, C => HIEFFPLA_NET_0_119327, Y => 
        HIEFFPLA_NET_0_119409);
    
    HIEFFPLA_INST_0_62466 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_6[0]\, 
        B => HIEFFPLA_NET_0_117096, S => HIEFFPLA_NET_0_117132, Y
         => HIEFFPLA_NET_0_115985);
    
    HIEFFPLA_INST_0_59079 : MX2
      port map(A => HIEFFPLA_NET_0_116677, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_23[1]\, S => 
        HIEFFPLA_NET_0_117214, Y => HIEFFPLA_NET_0_116437);
    
    HIEFFPLA_INST_0_59688 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_2[3]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_18[3]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_1[4]_net_1\, Y
         => HIEFFPLA_NET_0_116361);
    
    \U_ELK9_CH/U_SLAVE_1ELK/Q[4]\ : DFN1C0
      port map(D => \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/Q[4]_net_1\);
    
    HIEFFPLA_INST_0_51392 : MX2
      port map(A => HIEFFPLA_NET_0_117770, B => 
        \U_EXEC_MASTER/DEL_CNT[7]\, S => HIEFFPLA_NET_0_117796, Y
         => HIEFFPLA_NET_0_117788);
    
    HIEFFPLA_INST_0_48078 : AND2
      port map(A => \U_ELK16_CH/ELK_TX_DAT[0]\, B => 
        \U_ELK16_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118382);
    
    \U_ELK6_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL\ : DFN1C0
      port map(D => 
        \U_ELK6_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL_net_1\);
    
    HIEFFPLA_INST_0_57221 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_3[5]\, B => 
        HIEFFPLA_NET_0_116702, S => HIEFFPLA_NET_0_117120, Y => 
        HIEFFPLA_NET_0_116720);
    
    HIEFFPLA_INST_0_48949 : MX2
      port map(A => \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[1]_net_1\, 
        B => \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\, S => 
        \BIT_OS_SEL[2]\, Y => HIEFFPLA_NET_0_118220);
    
    \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[9]\ : DFN1C0
      port map(D => \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\);
    
    HIEFFPLA_INST_0_61766 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_26[0]\, B => 
        HIEFFPLA_NET_0_117096, S => HIEFFPLA_NET_0_117138, Y => 
        HIEFFPLA_NET_0_116080);
    
    \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[12]\ : DFN1C0
      port map(D => \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\, 
        CLK => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\);
    
    \U_ELK15_CH/U_SLAVE_1ELK/RECD_SER_WORD[4]\ : DFN1C0
      port map(D => \U_ELK15_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[4]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_15[4]\);
    
    HIEFFPLA_INST_0_43808 : AND2A
      port map(A => HIEFFPLA_NET_0_119208, B => 
        HIEFFPLA_NET_0_119568, Y => HIEFFPLA_NET_0_119209);
    
    \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[3]\ : DFN1C0
      port map(D => \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\);
    
    HIEFFPLA_INST_0_54085 : AND3
      port map(A => HIEFFPLA_NET_0_116649, B => 
        HIEFFPLA_NET_0_117334, C => HIEFFPLA_NET_0_117325, Y => 
        HIEFFPLA_NET_0_117310);
    
    HIEFFPLA_INST_0_55315 : AO1A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[4]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_0[8]_net_1\, C => 
        HIEFFPLA_NET_0_117068, Y => HIEFFPLA_NET_0_117062);
    
    \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_2[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117009, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_17_0, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_2[3]\);
    
    \U50_PATTERNS/SM_BANK_SEL[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119307, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_7, Q => 
        \U50_PATTERNS/SM_BANK_SEL[3]\);
    
    HIEFFPLA_INST_0_50385 : MX2
      port map(A => HIEFFPLA_NET_0_117948, B => 
        HIEFFPLA_NET_0_117946, S => \BIT_OS_SEL_5[1]\, Y => 
        HIEFFPLA_NET_0_117958);
    
    HIEFFPLA_INST_0_44062 : MX2
      port map(A => \U50_PATTERNS/TFC_STOP_ADDR_T[2]\, B => 
        \U50_PATTERNS/RD_USB_ADBUS[2]\, S => 
        HIEFFPLA_NET_0_119492, Y => HIEFFPLA_NET_0_119178);
    
    HIEFFPLA_INST_0_44576 : MX2
      port map(A => \ELKS_STOP_ADDR[3]\, B => 
        \U50_PATTERNS/U4D_REGCROSS/SAMP_TWO[3]_net_1\, S => 
        HIEFFPLA_NET_0_119093, Y => HIEFFPLA_NET_0_119088);
    
    \U_ELK14_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]\ : DFN1C0
      port map(D => \U_ELK14_CH/U_SLAVE_1ELK/Q[2]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]_net_1\);
    
    \U50_PATTERNS/ELINK_DINA_9[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119713, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_20, Q => 
        \U50_PATTERNS/ELINK_DINA_9[6]\);
    
    HIEFFPLA_INST_0_44771 : XO1
      port map(A => \OP_MODE_c_6[1]\, B => 
        \U50_PATTERNS/U4E_REGCROSS/SAMP_TWO[1]_net_1\, C => 
        HIEFFPLA_NET_0_119051, Y => HIEFFPLA_NET_0_119053);
    
    HIEFFPLA_INST_0_58866 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_20[1]\, B => 
        HIEFFPLA_NET_0_116459, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_1[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116466);
    
    HIEFFPLA_INST_0_51521 : NAND2
      port map(A => \U_EXEC_MASTER/PRESCALE[2]\, B => 
        \U_EXEC_MASTER/PRESCALE[1]\, Y => HIEFFPLA_NET_0_117755);
    
    HIEFFPLA_INST_0_46316 : NAND3C
      port map(A => HIEFFPLA_NET_0_119619, B => 
        HIEFFPLA_NET_0_119624, C => HIEFFPLA_NET_0_118884, Y => 
        HIEFFPLA_NET_0_118718);
    
    HIEFFPLA_INST_0_40261 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_0[3]\, B => 
        HIEFFPLA_NET_0_119574, S => HIEFFPLA_NET_0_119272, Y => 
        HIEFFPLA_NET_0_119868);
    
    \U200A_TFC/LOC_STRT_ADDR[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120275, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_5, Q => \U200A_TFC/LOC_STRT_ADDR[7]\);
    
    \U50_PATTERNS/ELINK_ADDRA_12[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120065, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_2_0, Q => 
        \U50_PATTERNS/ELINK_ADDRA_12[6]\);
    
    \U50_PATTERNS/ELINKS_STRT_ADDR[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120108, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_17, Q => 
        \U50_PATTERNS/ELINKS_STRT_ADDR[3]\);
    
    HIEFFPLA_INST_0_44335 : XO1
      port map(A => \U50_PATTERNS/U4A_REGCROSS/SAMP_TWO[6]_net_1\, 
        B => \TFC_STRT_ADDR[6]\, C => HIEFFPLA_NET_0_119137, Y
         => HIEFFPLA_NET_0_119138);
    
    HIEFFPLA_INST_0_54668 : MX2
      port map(A => HIEFFPLA_NET_0_117375, B => 
        HIEFFPLA_NET_0_117259, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[0]_net_1\, Y => 
        HIEFFPLA_NET_0_117225);
    
    HIEFFPLA_INST_0_41950 : NAND2B
      port map(A => \U50_PATTERNS/ELINK_RWA[1]\, B => 
        HIEFFPLA_NET_0_119648, Y => HIEFFPLA_NET_0_119649);
    
    HIEFFPLA_INST_0_42412 : AO1A
      port map(A => HIEFFPLA_NET_0_119019, B => 
        \U50_PATTERNS/RD_USB_ADBUS[6]\, C => 
        HIEFFPLA_NET_0_119535, Y => HIEFFPLA_NET_0_119543);
    
    HIEFFPLA_INST_0_48674 : MX2
      port map(A => \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\, 
        B => \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\, S => 
        \BIT_OS_SEL_0[2]\, Y => HIEFFPLA_NET_0_118268);
    
    HIEFFPLA_INST_0_46292 : NAND3C
      port map(A => HIEFFPLA_NET_0_119621, B => 
        HIEFFPLA_NET_0_119626, C => HIEFFPLA_NET_0_118888, Y => 
        HIEFFPLA_NET_0_118724);
    
    \U50_PATTERNS/U4E_REGCROSS/SAMP_TWO[0]\ : DFN1C0
      port map(D => \U50_PATTERNS/U4E_REGCROSS/SAMP_ONE[0]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_23, Q => 
        \U50_PATTERNS/U4E_REGCROSS/SAMP_TWO[0]_net_1\);
    
    \U50_PATTERNS/ELINK_ADDRA_2[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119997, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_21, Q => 
        \U50_PATTERNS/ELINK_ADDRA_2[2]\);
    
    HIEFFPLA_INST_0_51085 : AND2
      port map(A => \U_ELK9_CH/ELK_TX_DAT[1]\, B => 
        \U_ELK9_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_117838);
    
    HIEFFPLA_INST_0_38223 : AND2A
      port map(A => HIEFFPLA_NET_0_119452, B => 
        \U50_PATTERNS/RD_USB_ADBUS[0]\, Y => 
        HIEFFPLA_NET_0_120135);
    
    \U50_PATTERNS/ELINK_DINA_8[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119727, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_18, Q => 
        \U50_PATTERNS/ELINK_DINA_8[0]\);
    
    \U_ELK13_CH/U_SLAVE_1ELK/Q[8]\ : DFN1C0
      port map(D => \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/Q[8]_net_1\);
    
    HIEFFPLA_INST_0_57839 : AND3B
      port map(A => HIEFFPLA_NET_0_117179, B => 
        HIEFFPLA_NET_0_116605, C => HIEFFPLA_NET_0_116618, Y => 
        HIEFFPLA_NET_0_116609);
    
    HIEFFPLA_INST_0_43880 : MX2
      port map(A => HIEFFPLA_NET_0_119516, B => 
        \U50_PATTERNS/TFC_ADDRA[7]\, S => HIEFFPLA_NET_0_119294, 
        Y => HIEFFPLA_NET_0_119200);
    
    \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[4]\ : DFN1C0
      port map(D => 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\);
    
    HIEFFPLA_INST_0_51724 : NAND2B
      port map(A => 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM_0[4]_net_1\, B => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[79]_net_1\, Y => 
        HIEFFPLA_NET_0_117702);
    
    HIEFFPLA_INST_0_42900 : AND2B
      port map(A => \U50_PATTERNS/REG_STATE[5]_net_1\, B => 
        \U50_PATTERNS/REG_STATE[2]_net_1\, Y => 
        HIEFFPLA_NET_0_119429);
    
    HIEFFPLA_INST_0_42754 : AOI1C
      port map(A => HIEFFPLA_NET_0_119488, B => 
        HIEFFPLA_NET_0_119495, C => HIEFFPLA_NET_0_119513, Y => 
        HIEFFPLA_NET_0_119468);
    
    HIEFFPLA_INST_0_50109 : AND2A
      port map(A => \OP_MODE_c_4[1]\, B => \PATT_ELK_DAT_5[0]\, Y
         => HIEFFPLA_NET_0_118013);
    
    \U50_PATTERNS/ELINK_ADDRA_6[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119963, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_4, Q => 
        \U50_PATTERNS/ELINK_ADDRA_6[4]\);
    
    \U_ELK15_CH/U_ELK1_SERDAT_SOURCE/SERDAT[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118416, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_8, Q => 
        \U_ELK15_CH/ELK_TX_DAT[2]\);
    
    HIEFFPLA_INST_0_38250 : MX2
      port map(A => \U50_PATTERNS/ELINKS_STOP_ADDR[1]\, B => 
        \U50_PATTERNS/ELINKS_STOP_ADDR_T[1]\, S => 
        HIEFFPLA_NET_0_119472, Y => HIEFFPLA_NET_0_120126);
    
    \U_ELK2_CH/U_ELK1_CMD_TX/START_RISE\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118149, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_13, Q => 
        \U_ELK2_CH/U_ELK1_CMD_TX/START_RISE_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_SEL_5[0]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_BIT_OS_VAL[0]\, CLK
         => CLK_40M_GL, CLR => P_MASTER_POR_B_c_27_0, Q => 
        \BIT_OS_SEL_5[0]\);
    
    \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[0]\ : DFN1C0
      port map(D => 
        \U_ELK9_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\);
    
    HIEFFPLA_INST_0_57805 : NAND2A
      port map(A => HIEFFPLA_NET_0_116621, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_6[0]\, Y => 
        HIEFFPLA_NET_0_116617);
    
    HIEFFPLA_INST_0_52518 : MX2
      port map(A => HIEFFPLA_NET_0_117497, B => 
        HIEFFPLA_NET_0_117493, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_1[3]\, Y => 
        HIEFFPLA_NET_0_117553);
    
    \U50_PATTERNS/ELINK_ADDRA_16[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120038, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_8, Q => 
        \U50_PATTERNS/ELINK_ADDRA_16[1]\);
    
    HIEFFPLA_INST_0_57369 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_4[3]\, B => 
        HIEFFPLA_NET_0_116668, S => HIEFFPLA_NET_0_117122, Y => 
        HIEFFPLA_NET_0_116693);
    
    HIEFFPLA_INST_0_61394 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_5[3]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_21[3]\, S
         => \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_1[4]_net_1\, 
        Y => HIEFFPLA_NET_0_116132);
    
    \U_ELK19_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]\ : DFN1C0
      port map(D => \U_ELK19_CH/U_SLAVE_1ELK/Q[0]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]_net_1\);
    
    HIEFFPLA_INST_0_43650 : NAND3C
      port map(A => HIEFFPLA_NET_0_119274, B => 
        HIEFFPLA_NET_0_119281, C => HIEFFPLA_NET_0_119252, Y => 
        HIEFFPLA_NET_0_119255);
    
    HIEFFPLA_INST_0_55217 : NAND2B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[8]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[7]_net_1\, Y => 
        HIEFFPLA_NET_0_117084);
    
    HIEFFPLA_INST_0_43015 : NAND3C
      port map(A => HIEFFPLA_NET_0_118996, B => 
        HIEFFPLA_NET_0_119384, C => HIEFFPLA_NET_0_119401, Y => 
        HIEFFPLA_NET_0_119402);
    
    \U50_PATTERNS/ELINK_DINA_16[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119814, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_18, Q => 
        \U50_PATTERNS/ELINK_DINA_16[1]\);
    
    \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[5]\ : DFN1C0
      port map(D => 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\);
    
    HIEFFPLA_INST_0_53533 : MX2
      port map(A => HIEFFPLA_NET_0_117402, B => 
        HIEFFPLA_NET_0_117373, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[0]_net_1\, Y
         => HIEFFPLA_NET_0_117392);
    
    \U_ELK1_CH/U_SLAVE_1ELK/Q[5]\ : DFN1C0
      port map(D => \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/Q[5]_net_1\);
    
    \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[6]\ : DFN1C0
      port map(D => 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\);
    
    HIEFFPLA_INST_0_57967 : AO1A
      port map(A => HIEFFPLA_NET_0_116591, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_7[1]\, C => 
        HIEFFPLA_NET_0_116588, Y => HIEFFPLA_NET_0_116589);
    
    HIEFFPLA_INST_0_53708 : MX2
      port map(A => HIEFFPLA_NET_0_117272, B => 
        HIEFFPLA_NET_0_117257, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[2]_net_1\, Y
         => HIEFFPLA_NET_0_117368);
    
    HIEFFPLA_INST_0_37214 : OA1A
      port map(A => HIEFFPLA_NET_0_120328, B => 
        HIEFFPLA_NET_0_120293, C => 
        \U200A_TFC/GP_PG_SM[10]_net_1\, Y => 
        HIEFFPLA_NET_0_120323);
    
    HIEFFPLA_INST_0_42353 : NAND2B
      port map(A => \U50_PATTERNS/RD_USB_ADBUS[3]\, B => 
        \U50_PATTERNS/RD_USB_ADBUS[2]\, Y => 
        HIEFFPLA_NET_0_119559);
    
    HIEFFPLA_INST_0_37607 : AOI1A
      port map(A => \ELKS_STRT_ADDR[7]\, B => 
        HIEFFPLA_NET_0_120219, C => HIEFFPLA_NET_0_120247, Y => 
        HIEFFPLA_NET_0_120248);
    
    HIEFFPLA_INST_0_56251 : AND3B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/RECD_SER_WORD[0]_net_1\, 
        B => 
        \U_MASTER_DES/U13C_MASTER_DESER/RECD_SER_WORD[4]_net_1\, 
        C => 
        \U_MASTER_DES/U13C_MASTER_DESER/RECD_SER_WORD[3]_net_1\, 
        Y => HIEFFPLA_NET_0_116907);
    
    HIEFFPLA_INST_0_44054 : MX2
      port map(A => \U50_PATTERNS/TFC_STOP_ADDR_T[1]\, B => 
        \U50_PATTERNS/RD_USB_ADBUS[1]\, S => 
        HIEFFPLA_NET_0_119492, Y => HIEFFPLA_NET_0_119179);
    
    HIEFFPLA_INST_0_39866 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_9[0]\, B => 
        HIEFFPLA_NET_0_119524, S => HIEFFPLA_NET_0_119292, Y => 
        HIEFFPLA_NET_0_119943);
    
    HIEFFPLA_INST_0_38322 : MX2
      port map(A => \U50_PATTERNS/ELINKS_STOP_ADDR_T[2]\, B => 
        \U50_PATTERNS/RD_USB_ADBUS[2]\, S => 
        HIEFFPLA_NET_0_119413, Y => HIEFFPLA_NET_0_120117);
    
    \U_ELK6_CH/U_ELK1_SERDAT_SOURCE/SERDAT[6]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117962, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_2, Q => 
        \U_ELK6_CH/ELK_TX_DAT[6]\);
    
    HIEFFPLA_INST_0_58677 : AO1C
      port map(A => HIEFFPLA_NET_0_117204, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_18[2]\, C => 
        HIEFFPLA_NET_0_117231, Y => HIEFFPLA_NET_0_116489);
    
    \U50_PATTERNS/ELINK_DINA_6[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119737, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_16, Q => 
        \U50_PATTERNS/ELINK_DINA_6[6]\);
    
    HIEFFPLA_INST_0_51324 : AO1
      port map(A => \U_EXEC_MASTER/CCC_1_LOCK_STAT_1D_net_1\, B
         => HIEFFPLA_NET_0_117797, C => HIEFFPLA_NET_0_117787, Y
         => HIEFFPLA_NET_0_117796);
    
    HIEFFPLA_INST_0_48021 : MX2
      port map(A => HIEFFPLA_NET_0_118407, B => 
        HIEFFPLA_NET_0_118404, S => \BIT_OS_SEL_3[0]\, Y => 
        \U_ELK15_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[4]\);
    
    HIEFFPLA_INST_0_44400 : MX2
      port map(A => \TFC_STOP_ADDR[7]\, B => 
        \U50_PATTERNS/U4B_REGCROSS/SAMP_TWO[7]_net_1\, S => 
        HIEFFPLA_NET_0_119135, Y => HIEFFPLA_NET_0_119126);
    
    HIEFFPLA_INST_0_37601 : AOI1A
      port map(A => \ELKS_STRT_ADDR[5]\, B => 
        HIEFFPLA_NET_0_120219, C => HIEFFPLA_NET_0_120249, Y => 
        HIEFFPLA_NET_0_120250);
    
    AFLSDF_INV_20 : INV
      port map(A => DCB_SALT_SEL_c, Y => \AFLSDF_INV_20\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/MAX_CNT[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_116951, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_16, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/MAX_CNT[3]\);
    
    \U_ELK11_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118602, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_7, Q => 
        \U_ELK11_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]_net_1\);
    
    \U_ELK10_CH/U_SLAVE_1ELK/RECD_SER_WORD[4]\ : DFN1C0
      port map(D => \U_ELK10_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[4]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_10[4]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_1[6]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116782, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_4, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_1[6]\);
    
    HIEFFPLA_INST_0_56202 : XA1C
      port map(A => HIEFFPLA_NET_0_116929, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/MAX_CNT[8]\, C => 
        HIEFFPLA_NET_0_117112, Y => HIEFFPLA_NET_0_116931);
    
    HIEFFPLA_INST_0_41931 : AND3C
      port map(A => HIEFFPLA_NET_0_119271, B => 
        HIEFFPLA_NET_0_119262, C => 
        \U50_PATTERNS/SM_BANK_SEL[10]\, Y => 
        HIEFFPLA_NET_0_119657);
    
    \U50_PATTERNS/TFC_STOP_ADDR[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119187, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_8, Q => 
        \U50_PATTERNS/TFC_STOP_ADDR[1]\);
    
    \U_ELK15_CH/U_SLAVE_1ELK/Q[8]\ : DFN1C0
      port map(D => \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/Q[8]_net_1\);
    
    \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[8]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117700, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_31, Q => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[8]_net_1\);
    
    \U_ELK1_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL\ : DFN1C0
      port map(D => \U_ELK1_CH/ELK_IN_R_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL_net_1\);
    
    \U50_PATTERNS/ELINK_DINA_8[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119722, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_18, Q => 
        \U50_PATTERNS/ELINK_DINA_8[5]\);
    
    HIEFFPLA_INST_0_63018 : AND3A
      port map(A => HIEFFPLA_NET_0_115911, B => 
        HIEFFPLA_NET_0_115899, C => HIEFFPLA_NET_0_115901, Y => 
        HIEFFPLA_NET_0_115913);
    
    HIEFFPLA_INST_0_53467 : AOI1
      port map(A => HIEFFPLA_NET_0_117337, B => 
        HIEFFPLA_NET_0_116593, C => HIEFFPLA_NET_0_117403, Y => 
        HIEFFPLA_NET_0_117404);
    
    HIEFFPLA_INST_0_41251 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_4[1]\, B => 
        HIEFFPLA_NET_0_119576, S => HIEFFPLA_NET_0_119284, Y => 
        HIEFFPLA_NET_0_119758);
    
    \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[0]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_SER_IN_R_1DEL_net_1\, 
        CLK => CCC_160M_ADJ, CLR => P_MASTER_POR_B_c_34_0, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[0]_net_1\);
    
    \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[48]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117724, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_19, Q => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[48]\);
    
    \U_ELK18_CH/U_ELK1_SERDAT_SOURCE/SERDAT[6]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118277, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_13, Q => 
        \U_ELK18_CH/ELK_TX_DAT[6]\);
    
    \U_MASTER_DES/U13A_ADJ_160M/BITCNT[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117691, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_14, Q => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[7]\);
    
    HIEFFPLA_INST_0_58296 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_13[3]\, B => 
        HIEFFPLA_NET_0_116534, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_1[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116539);
    
    HIEFFPLA_INST_0_43020 : AND3B
      port map(A => \U50_PATTERNS/USB_RXF_B\, B => 
        \U50_PATTERNS/REG_STATE[4]_net_1\, C => 
        \U50_PATTERNS/REG_STATE[3]_net_1\, Y => 
        HIEFFPLA_NET_0_119400);
    
    HIEFFPLA_INST_0_111367 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_18[0]\, B => 
        HIEFFPLA_NET_0_116735, S => HIEFFPLA_NET_0_117204, Y => 
        HIEFFPLA_NET_0_116484);
    
    HIEFFPLA_INST_0_61157 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_1[4]\, 
        B => HIEFFPLA_NET_0_117166, S => HIEFFPLA_NET_0_117149, Y
         => HIEFFPLA_NET_0_116166);
    
    \U50_PATTERNS/U4A_REGCROSS/LOCAL_REG_VAL[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119154, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_17, Q => \TFC_STRT_ADDR[0]\);
    
    HIEFFPLA_INST_0_111285 : MX2A
      port map(A => HIEFFPLA_NET_0_115843, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_29[3]\, S => 
        HIEFFPLA_NET_0_117395, Y => HIEFFPLA_NET_0_116368);
    
    \U_ELK3_CH/U_SLAVE_1ELK/Q[1]\ : DFN1C0
      port map(D => \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/Q[1]_net_1\);
    
    HIEFFPLA_INST_0_40693 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_15[3]\, B => 
        HIEFFPLA_NET_0_119574, S => HIEFFPLA_NET_0_119297, Y => 
        HIEFFPLA_NET_0_119820);
    
    \U50_PATTERNS/ELINKS_STOP_ADDR_T[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120119, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_7, Q => 
        \U50_PATTERNS/ELINKS_STOP_ADDR_T[0]\);
    
    \U200B_ELINKS/GP_PG_SM[8]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120206, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_29, Q => 
        \U200B_ELINKS/GP_PG_SM[8]_net_1\);
    
    HIEFFPLA_INST_0_56249 : AND2A
      port map(A => DCB_SALT_SEL_c, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/RECD_SER_WORD[7]_net_1\, 
        Y => \TFC_RX_SER_WORD[7]\);
    
    HIEFFPLA_INST_0_43061 : AND3B
      port map(A => HIEFFPLA_NET_0_119451, B => 
        HIEFFPLA_NET_0_119422, C => HIEFFPLA_NET_0_119021, Y => 
        HIEFFPLA_NET_0_119389);
    
    \U_ELK10_CH/U_SLAVE_1ELK/Q[1]\ : DFN1C0
      port map(D => \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/Q[1]_net_1\);
    
    HIEFFPLA_INST_0_58041 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_0[0]\, B => 
        HIEFFPLA_NET_0_116680, S => HIEFFPLA_NET_0_117088, Y => 
        HIEFFPLA_NET_0_116572);
    
    HIEFFPLA_INST_0_49226 : MX2
      port map(A => HIEFFPLA_NET_0_118175, B => 
        HIEFFPLA_NET_0_118173, S => \BIT_OS_SEL_0[1]\, Y => 
        HIEFFPLA_NET_0_118170);
    
    HIEFFPLA_INST_0_57814 : XA1B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_6[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_6[0]\, C => 
        HIEFFPLA_NET_0_117179, Y => HIEFFPLA_NET_0_116615);
    
    \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[12]\ : DFN1C0
      port map(D => \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\);
    
    \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[10]\ : DFN1C0
      port map(D => 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\);
    
    \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[8]\ : DFN1C0
      port map(D => 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\);
    
    \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[11]\ : DFN1C0
      port map(D => 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[11]_net_1\);
    
    HIEFFPLA_INST_0_61370 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_5[1]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_21[1]\, S
         => \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_1[4]_net_1\, 
        Y => HIEFFPLA_NET_0_116136);
    
    HIEFFPLA_INST_0_43497 : MX2
      port map(A => \U50_PATTERNS/SM_BANK_SEL[6]\, B => 
        HIEFFPLA_NET_0_119212, S => HIEFFPLA_NET_0_118691, Y => 
        HIEFFPLA_NET_0_119304);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_1[8]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116780, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_4, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_1[8]\);
    
    \U50_PATTERNS/U4B_REGCROSS/LOCAL_REG_VAL[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119131, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_19, Q => \TFC_STOP_ADDR[2]\);
    
    HIEFFPLA_INST_0_39209 : MX2
      port map(A => HIEFFPLA_NET_0_119516, B => 
        \U50_PATTERNS/ELINK_ADDRA_18[7]\, S => 
        HIEFFPLA_NET_0_119264, Y => HIEFFPLA_NET_0_120016);
    
    \U_ELK13_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0\ : DFN1C0
      port map(D => CLK_40M_GL, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_6, Q => 
        \U_ELK13_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0_net_1\);
    
    HIEFFPLA_INST_0_42783 : AOI1C
      port map(A => HIEFFPLA_NET_0_119496, B => 
        HIEFFPLA_NET_0_119636, C => 
        \U50_PATTERNS/REG_STATE_0[4]_net_1\, Y => 
        HIEFFPLA_NET_0_119463);
    
    \U_ELK19_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U3\ : IOBI_ID_OD_EB
      port map(DR => \U_ELK19_CH/ELK_OUT_R\, DF => 
        \U_ELK19_CH/ELK_OUT_F\, CLR => \GND\, E => 
        \AFLSDF_INV_33\, ICLK => CCC_160M_ADJ, OCLK => 
        CCC_160M_FXD, YIN => 
        \U_ELK19_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\, DOUT => 
        OPEN, EOUT => 
        \U_ELK19_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET3\, YR => OPEN, 
        YF => OPEN);
    
    \U_ELK13_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL\ : DFN1C0
      port map(D => \U_ELK13_CH/ELK_IN_F_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL_net_1\);
    
    \U50_PATTERNS/SM_BANK_SEL[9]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119301, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_8, Q => 
        \U50_PATTERNS/SM_BANK_SEL[9]\);
    
    HIEFFPLA_INST_0_50614 : NAND2B
      port map(A => \OP_MODE_c_4[1]\, B => \PATT_ELK_DAT_7[7]\, Y
         => HIEFFPLA_NET_0_117916);
    
    HIEFFPLA_INST_0_45858 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_18[2]\, C => 
        \U50_PATTERNS/SM_BANK_SEL[1]\, Y => HIEFFPLA_NET_0_118826);
    
    HIEFFPLA_INST_0_45602 : AO1A
      port map(A => HIEFFPLA_NET_0_119428, B => 
        \U50_PATTERNS/ELINKS_STRT_ADDR[7]\, C => 
        HIEFFPLA_NET_0_118788, Y => HIEFFPLA_NET_0_118882);
    
    HIEFFPLA_INST_0_38948 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_15[2]\, B => 
        HIEFFPLA_NET_0_119522, S => HIEFFPLA_NET_0_119297, Y => 
        HIEFFPLA_NET_0_120045);
    
    \U50_PATTERNS/TFC_DINA[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119190, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_4, Q => \U50_PATTERNS/TFC_DINA[7]\);
    
    \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_2S_4\ : DFN1C0
      port map(D => 
        \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_1S_net_1\, CLK
         => CLK60MHZ, CLR => P_MASTER_POR_B_c_0_0, Q => 
        P_USB_MASTER_EN_c_4);
    
    HIEFFPLA_INST_0_56091 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/MAX_CNT[3]\, 
        B => HIEFFPLA_NET_0_116936, S => HIEFFPLA_NET_0_117084, Y
         => HIEFFPLA_NET_0_116951);
    
    HIEFFPLA_INST_0_40405 : MX2
      port map(A => HIEFFPLA_NET_0_119574, B => 
        \U50_PATTERNS/ELINK_DINA_11[3]\, S => 
        HIEFFPLA_NET_0_119280, Y => HIEFFPLA_NET_0_119852);
    
    \U50_PATTERNS/SM_BANK_SEL[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119308, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_7, Q => 
        \U50_PATTERNS/SM_BANK_SEL[2]\);
    
    HIEFFPLA_INST_0_46225 : AO1A
      port map(A => HIEFFPLA_NET_0_118918, B => 
        \U50_PATTERNS/SM_BANK_SEL[15]\, C => 
        HIEFFPLA_NET_0_118737, Y => HIEFFPLA_NET_0_118738);
    
    HIEFFPLA_INST_0_58360 : MX2A
      port map(A => HIEFFPLA_NET_0_116774, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_13[3]\, S => 
        HIEFFPLA_NET_0_117396, Y => HIEFFPLA_NET_0_116530);
    
    HIEFFPLA_INST_0_42980 : AND3B
      port map(A => \U50_PATTERNS/REG_STATE[3]_net_1\, B => 
        \U50_PATTERNS/USB_RXF_B\, C => 
        \U50_PATTERNS/REG_STATE[2]_net_1\, Y => 
        HIEFFPLA_NET_0_119411);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_31[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116019, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_10, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_31[1]\);
    
    HIEFFPLA_INST_0_60063 : MX2
      port map(A => HIEFFPLA_NET_0_116815, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_5[3]\, S => 
        HIEFFPLA_NET_0_117218, Y => HIEFFPLA_NET_0_116315);
    
    HIEFFPLA_INST_0_48431 : MX2
      port map(A => \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\, 
        B => \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\, S => 
        \BIT_OS_SEL_0[2]\, Y => HIEFFPLA_NET_0_118312);
    
    HIEFFPLA_INST_0_47670 : MX2
      port map(A => \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\, 
        B => \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\, S => 
        \BIT_OS_SEL_2[2]\, Y => HIEFFPLA_NET_0_118449);
    
    HIEFFPLA_INST_0_38597 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_10[3]\, B => 
        HIEFFPLA_NET_0_119520, S => HIEFFPLA_NET_0_119239, Y => 
        HIEFFPLA_NET_0_120084);
    
    \U_ELK18_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118289, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_3, Q => 
        \U_ELK18_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]_net_1\);
    
    HIEFFPLA_INST_0_61604 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_24[2]\, B => 
        HIEFFPLA_NET_0_117181, S => HIEFFPLA_NET_0_117074, Y => 
        HIEFFPLA_NET_0_116103);
    
    HIEFFPLA_INST_0_52105 : AND3C
      port map(A => HIEFFPLA_NET_0_117667, B => 
        HIEFFPLA_NET_0_117666, C => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[4]\, Y => 
        HIEFFPLA_NET_0_117635);
    
    HIEFFPLA_INST_0_58326 : AO1A
      port map(A => HIEFFPLA_NET_0_117396, B => 
        HIEFFPLA_NET_0_116589, C => HIEFFPLA_NET_0_116529, Y => 
        HIEFFPLA_NET_0_116533);
    
    HIEFFPLA_INST_0_44796 : XOR2
      port map(A => \U50_PATTERNS/U4E_REGCROSS/DELCNT[0]_net_1\, 
        B => \U50_PATTERNS/U4E_REGCROSS/DELCNT[1]_net_1\, Y => 
        HIEFFPLA_NET_0_119046);
    
    \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[0]\ : DFN1C0
      port map(D => 
        \U_ELK2_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\);
    
    HIEFFPLA_INST_0_37736 : NAND2B
      port map(A => HIEFFPLA_NET_0_120190, B => 
        HIEFFPLA_NET_0_120226, Y => HIEFFPLA_NET_0_120220);
    
    \U_ELK9_CH/U_SLAVE_1ELK/Q[14]\ : DFN1C0
      port map(D => \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[14]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/Q[14]_net_1\);
    
    \U50_PATTERNS/U104_PATT_ELINK_BLK/DPRT_512X9_SRAM_R0C0\ : 
        RAM4K9
      generic map(MEMORYFILE => "DPRT_512X9_SRAM_R0C0.mem")

      port map(ADDRA11 => AFLSDF_GND, ADDRA10 => AFLSDF_GND, 
        ADDRA9 => AFLSDF_GND, ADDRA8 => \GND\, ADDRA7 => 
        \U50_PATTERNS/ELINK_ADDRA_4[7]\, ADDRA6 => 
        \U50_PATTERNS/ELINK_ADDRA_4[6]\, ADDRA5 => 
        \U50_PATTERNS/ELINK_ADDRA_4[5]\, ADDRA4 => 
        \U50_PATTERNS/ELINK_ADDRA_4[4]\, ADDRA3 => 
        \U50_PATTERNS/ELINK_ADDRA_4[3]\, ADDRA2 => 
        \U50_PATTERNS/ELINK_ADDRA_4[2]\, ADDRA1 => 
        \U50_PATTERNS/ELINK_ADDRA_4[1]\, ADDRA0 => 
        \U50_PATTERNS/ELINK_ADDRA_4[0]\, ADDRB11 => AFLSDF_GND, 
        ADDRB10 => AFLSDF_GND, ADDRB9 => AFLSDF_GND, ADDRB8 => 
        \GND\, ADDRB7 => \ELKS_ADDRB[7]\, ADDRB6 => 
        \ELKS_ADDRB[6]\, ADDRB5 => \ELKS_ADDRB[5]\, ADDRB4 => 
        \ELKS_ADDRB[4]\, ADDRB3 => \ELKS_ADDRB[3]\, ADDRB2 => 
        \ELKS_ADDRB[2]\, ADDRB1 => \ELKS_ADDRB[1]\, ADDRB0 => 
        \ELKS_ADDRB[0]\, DINA8 => \GND\, DINA7 => 
        \U50_PATTERNS/ELINK_DINA_4[7]\, DINA6 => 
        \U50_PATTERNS/ELINK_DINA_4[6]\, DINA5 => 
        \U50_PATTERNS/ELINK_DINA_4[5]\, DINA4 => 
        \U50_PATTERNS/ELINK_DINA_4[4]\, DINA3 => 
        \U50_PATTERNS/ELINK_DINA_4[3]\, DINA2 => 
        \U50_PATTERNS/ELINK_DINA_4[2]\, DINA1 => 
        \U50_PATTERNS/ELINK_DINA_4[1]\, DINA0 => 
        \U50_PATTERNS/ELINK_DINA_4[0]\, DINB8 => \GND\, DINB7 => 
        \ELK_RX_SER_WORD_4[7]\, DINB6 => \ELK_RX_SER_WORD_4[6]\, 
        DINB5 => \ELK_RX_SER_WORD_4[5]\, DINB4 => 
        \ELK_RX_SER_WORD_4[4]\, DINB3 => \ELK_RX_SER_WORD_4[3]\, 
        DINB2 => \ELK_RX_SER_WORD_4[2]\, DINB1 => 
        \ELK_RX_SER_WORD_4[1]\, DINB0 => \ELK_RX_SER_WORD_4[0]\, 
        WIDTHA0 => \VCC\, WIDTHA1 => \VCC\, WIDTHB0 => \VCC\, 
        WIDTHB1 => \VCC\, PIPEA => \VCC\, PIPEB => \VCC\, WMODEA
         => \GND\, WMODEB => \GND\, BLKA => 
        \U50_PATTERNS/ELINK_BLKA[4]\, BLKB => ELKS_RAM_BLKB_EN, 
        WENA => \U50_PATTERNS/ELINK_RWA[4]\, WENB => ELKS_RWB, 
        CLKA => CLK60MHZ, CLKB => CLK_40M_GL, RESET => 
        P_USB_MASTER_EN_c_0, DOUTA8 => OPEN, DOUTA7 => 
        \U50_PATTERNS/ELINK_DOUTA_4[7]\, DOUTA6 => 
        \U50_PATTERNS/ELINK_DOUTA_4[6]\, DOUTA5 => 
        \U50_PATTERNS/ELINK_DOUTA_4[5]\, DOUTA4 => 
        \U50_PATTERNS/ELINK_DOUTA_4[4]\, DOUTA3 => 
        \U50_PATTERNS/ELINK_DOUTA_4[3]\, DOUTA2 => 
        \U50_PATTERNS/ELINK_DOUTA_4[2]\, DOUTA1 => 
        \U50_PATTERNS/ELINK_DOUTA_4[1]\, DOUTA0 => 
        \U50_PATTERNS/ELINK_DOUTA_4[0]\, DOUTB8 => OPEN, DOUTB7
         => \PATT_ELK_DAT_4[7]\, DOUTB6 => \PATT_ELK_DAT_4[6]\, 
        DOUTB5 => \PATT_ELK_DAT_4[5]\, DOUTB4 => 
        \PATT_ELK_DAT_4[4]\, DOUTB3 => \PATT_ELK_DAT_4[3]\, 
        DOUTB2 => \PATT_ELK_DAT_4[2]\, DOUTB1 => 
        \PATT_ELK_DAT_4[1]\, DOUTB0 => \PATT_ELK_DAT_4[0]\);
    
    \U_ELK8_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]\ : DFN1C0
      port map(D => \U_ELK8_CH/U_SLAVE_1ELK/Q[8]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]_net_1\);
    
    HIEFFPLA_INST_0_58939 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_21[0]\, B => 
        HIEFFPLA_NET_0_116680, S => HIEFFPLA_NET_0_117093, Y => 
        HIEFFPLA_NET_0_116456);
    
    \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[9]\ : DFN1C0
      port map(D => 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\);
    
    HIEFFPLA_INST_0_59853 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_31[1]\, B => 
        HIEFFPLA_NET_0_116677, S => HIEFFPLA_NET_0_117097, Y => 
        HIEFFPLA_NET_0_116342);
    
    HIEFFPLA_INST_0_42329 : AND3
      port map(A => HIEFFPLA_NET_0_119429, B => 
        HIEFFPLA_NET_0_119561, C => HIEFFPLA_NET_0_119568, Y => 
        HIEFFPLA_NET_0_119569);
    
    HIEFFPLA_INST_0_56235 : AND2A
      port map(A => DCB_SALT_SEL_c, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/RECD_SER_WORD[0]_net_1\, 
        Y => \TFC_RX_SER_WORD[0]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/PHASE_ADJ[3]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[3]_net_1\, CLK
         => CLK_40M_GL, CLR => P_MASTER_POR_B_c, Q => 
        \U_MASTER_DES/PHASE_ADJ_160_L[3]\);
    
    \U50_PATTERNS/ELINK_ADDRA_14[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120053, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_5, Q => 
        \U50_PATTERNS/ELINK_ADDRA_14[2]\);
    
    \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_2S_20\ : DFN1C0
      port map(D => 
        \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_1S_0_net_1\, CLK
         => CLK60MHZ, CLR => \U_EXEC_MASTER/P_MASTER_POR_B_c_0\, 
        Q => P_USB_MASTER_EN_c_20);
    
    HIEFFPLA_INST_0_50856 : AND2A
      port map(A => \OP_MODE_c_0[1]\, B => \PATT_ELK_DAT_8[0]\, Y
         => HIEFFPLA_NET_0_117878);
    
    HIEFFPLA_INST_0_37317 : AND3A
      port map(A => \U200A_TFC/N_232_li\, B => 
        HIEFFPLA_NET_0_120333, C => \U200A_TFC/GP_PG_SM[9]_net_1\, 
        Y => HIEFFPLA_NET_0_120296);
    
    \U_ELK18_CH/U_SLAVE_1ELK/RECD_SER_WORD[5]\ : DFN1C0
      port map(D => \U_ELK18_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[5]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_18[5]\);
    
    HIEFFPLA_INST_0_52221 : AND2
      port map(A => \U_MASTER_DES/CCC_RX_CLK_LOCK\, B => 
        CCC_MAIN_LOCK, Y => ALL_PLL_LOCK_c);
    
    HIEFFPLA_INST_0_39290 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_1[0]\, B => 
        HIEFFPLA_NET_0_119524, S => HIEFFPLA_NET_0_119243, Y => 
        HIEFFPLA_NET_0_120007);
    
    HIEFFPLA_INST_0_37604 : AO1A
      port map(A => HIEFFPLA_NET_0_120240, B => 
        HIEFFPLA_NET_0_120234, C => HIEFFPLA_NET_0_120237, Y => 
        HIEFFPLA_NET_0_120249);
    
    \U_ELK9_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]\ : DFN1C0
      port map(D => \U_ELK9_CH/U_SLAVE_1ELK/Q[14]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]_net_1\);
    
    HIEFFPLA_INST_0_47290 : MX2
      port map(A => HIEFFPLA_NET_0_118536, B => 
        HIEFFPLA_NET_0_118532, S => \BIT_OS_SEL_5[0]\, Y => 
        \U_ELK12_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[6]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_0[8]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116816, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_3, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_0[8]\);
    
    \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[2]\\\\/U0/U0\ : 
        IOPAD_BI_U
      port map(D => 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[2]\\\\/U0/NET1\, 
        E => 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[2]\\\\/U0/NET2\, 
        Y => 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[2]\\\\/U0/NET3\, 
        PAD => BIDIR_USB_ADBUS(2));
    
    HIEFFPLA_INST_0_37681 : NAND2B
      port map(A => \U200B_ELINKS/GP_PG_SM[4]_net_1\, B => 
        \U200B_ELINKS/GP_PG_SM[5]_net_1\, Y => 
        HIEFFPLA_NET_0_120231);
    
    \U_ELK4_CH/U_SLAVE_1ELK/Q[7]\ : DFN1C0
      port map(D => \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/Q[7]_net_1\);
    
    \U50_PATTERNS/U101_PATT_ELINK_BLK/DPRT_512X9_SRAM_R0C0\ : 
        RAM4K9
      generic map(MEMORYFILE => "DPRT_512X9_SRAM_R0C0.mem")

      port map(ADDRA11 => AFLSDF_GND, ADDRA10 => AFLSDF_GND, 
        ADDRA9 => AFLSDF_GND, ADDRA8 => \GND\, ADDRA7 => 
        \U50_PATTERNS/ELINK_ADDRA_1[7]\, ADDRA6 => 
        \U50_PATTERNS/ELINK_ADDRA_1[6]\, ADDRA5 => 
        \U50_PATTERNS/ELINK_ADDRA_1[5]\, ADDRA4 => 
        \U50_PATTERNS/ELINK_ADDRA_1[4]\, ADDRA3 => 
        \U50_PATTERNS/ELINK_ADDRA_1[3]\, ADDRA2 => 
        \U50_PATTERNS/ELINK_ADDRA_1[2]\, ADDRA1 => 
        \U50_PATTERNS/ELINK_ADDRA_1[1]\, ADDRA0 => 
        \U50_PATTERNS/ELINK_ADDRA_1[0]\, ADDRB11 => AFLSDF_GND, 
        ADDRB10 => AFLSDF_GND, ADDRB9 => AFLSDF_GND, ADDRB8 => 
        \GND\, ADDRB7 => \ELKS_ADDRB[7]\, ADDRB6 => 
        \ELKS_ADDRB_0[6]\, ADDRB5 => \ELKS_ADDRB[5]\, ADDRB4 => 
        \ELKS_ADDRB_0[4]\, ADDRB3 => \ELKS_ADDRB[3]\, ADDRB2 => 
        \ELKS_ADDRB_0[2]\, ADDRB1 => \ELKS_ADDRB[1]\, ADDRB0 => 
        \ELKS_ADDRB[0]\, DINA8 => \GND\, DINA7 => 
        \U50_PATTERNS/ELINK_DINA_1[7]\, DINA6 => 
        \U50_PATTERNS/ELINK_DINA_1[6]\, DINA5 => 
        \U50_PATTERNS/ELINK_DINA_1[5]\, DINA4 => 
        \U50_PATTERNS/ELINK_DINA_1[4]\, DINA3 => 
        \U50_PATTERNS/ELINK_DINA_1[3]\, DINA2 => 
        \U50_PATTERNS/ELINK_DINA_1[2]\, DINA1 => 
        \U50_PATTERNS/ELINK_DINA_1[1]\, DINA0 => 
        \U50_PATTERNS/ELINK_DINA_1[0]\, DINB8 => \GND\, DINB7 => 
        \ELK_RX_SER_WORD_1[7]\, DINB6 => \ELK_RX_SER_WORD_1[6]\, 
        DINB5 => \ELK_RX_SER_WORD_1[5]\, DINB4 => 
        \ELK_RX_SER_WORD_1[4]\, DINB3 => \ELK_RX_SER_WORD_1[3]\, 
        DINB2 => \ELK_RX_SER_WORD_1[2]\, DINB1 => 
        \ELK_RX_SER_WORD_1[1]\, DINB0 => \ELK_RX_SER_WORD_1[0]\, 
        WIDTHA0 => \VCC\, WIDTHA1 => \VCC\, WIDTHB0 => \VCC\, 
        WIDTHB1 => \VCC\, PIPEA => \VCC\, PIPEB => \VCC\, WMODEA
         => \GND\, WMODEB => \GND\, BLKA => 
        \U50_PATTERNS/ELINK_BLKA[1]\, BLKB => ELKS_RAM_BLKB_EN, 
        WENA => \U50_PATTERNS/ELINK_RWA[1]\, WENB => ELKS_RWB, 
        CLKA => CLK60MHZ, CLKB => CLK_40M_GL, RESET => 
        P_USB_MASTER_EN_c_0, DOUTA8 => OPEN, DOUTA7 => 
        \U50_PATTERNS/ELINK_DOUTA_1[7]\, DOUTA6 => 
        \U50_PATTERNS/ELINK_DOUTA_1[6]\, DOUTA5 => 
        \U50_PATTERNS/ELINK_DOUTA_1[5]\, DOUTA4 => 
        \U50_PATTERNS/ELINK_DOUTA_1[4]\, DOUTA3 => 
        \U50_PATTERNS/ELINK_DOUTA_1[3]\, DOUTA2 => 
        \U50_PATTERNS/ELINK_DOUTA_1[2]\, DOUTA1 => 
        \U50_PATTERNS/ELINK_DOUTA_1[1]\, DOUTA0 => 
        \U50_PATTERNS/ELINK_DOUTA_1[0]\, DOUTB8 => OPEN, DOUTB7
         => \PATT_ELK_DAT_1[7]\, DOUTB6 => \PATT_ELK_DAT_1[6]\, 
        DOUTB5 => \PATT_ELK_DAT_1[5]\, DOUTB4 => 
        \PATT_ELK_DAT_1[4]\, DOUTB3 => \PATT_ELK_DAT_1[3]\, 
        DOUTB2 => \PATT_ELK_DAT_1[2]\, DOUTB1 => 
        \PATT_ELK_DAT_1[1]\, DOUTB0 => \PATT_ELK_DAT_1[0]\);
    
    HIEFFPLA_INST_0_50208 : MX2
      port map(A => \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\, B
         => \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[13]_net_1\, S => 
        \BIT_OS_SEL_6[2]\, Y => HIEFFPLA_NET_0_117992);
    
    HIEFFPLA_INST_0_55301 : AO1A
      port map(A => HIEFFPLA_NET_0_117109, B => 
        HIEFFPLA_NET_0_116813, C => HIEFFPLA_NET_0_117066, Y => 
        HIEFFPLA_NET_0_117067);
    
    HIEFFPLA_INST_0_42519 : OA1A
      port map(A => HIEFFPLA_NET_0_119433, B => 
        HIEFFPLA_NET_0_119010, C => \U50_PATTERNS/REG_ADDR[0]\, Y
         => HIEFFPLA_NET_0_119524);
    
    HIEFFPLA_INST_0_49871 : MX2
      port map(A => HIEFFPLA_NET_0_118040, B => 
        HIEFFPLA_NET_0_118037, S => \BIT_OS_SEL_6[1]\, Y => 
        HIEFFPLA_NET_0_118050);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_4[6]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116690, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_9, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_4[6]\);
    
    \U_ELK16_CH/U_ELK1_SERDAT_SOURCE/SERDAT[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118370, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_9, Q => 
        \U_ELK16_CH/ELK_TX_DAT[3]\);
    
    \U50_PATTERNS/ELINK_DINA_7[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119732, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_17, Q => 
        \U50_PATTERNS/ELINK_DINA_7[3]\);
    
    \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[10]\ : DFN1C0
      port map(D => \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\);
    
    HIEFFPLA_INST_0_37830 : AND3B
      port map(A => \U200B_ELINKS/GP_PG_SM[2]_net_1\, B => 
        HIEFFPLA_NET_0_120195, C => 
        \U200B_ELINKS/GP_PG_SM[3]_net_1\, Y => 
        HIEFFPLA_NET_0_120196);
    
    \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_2S\ : DFN1C0
      port map(D => 
        \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_1S_net_1\, CLK
         => CLK60MHZ, CLR => P_MASTER_POR_B_c_22_0, Q => 
        P_USB_MASTER_EN_c);
    
    \U_ELK1_CH/U_SLAVE_1ELK/Q[10]\ : DFN1C0
      port map(D => \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/Q[10]_net_1\);
    
    \U_ELK15_CH/U_SLAVE_1ELK/Q[1]\ : DFN1C0
      port map(D => \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/Q[1]_net_1\);
    
    HIEFFPLA_INST_0_40243 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_0[1]\, B => 
        HIEFFPLA_NET_0_119576, S => HIEFFPLA_NET_0_119272, Y => 
        HIEFFPLA_NET_0_119870);
    
    \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[3]\ : DFN1C0
      port map(D => \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\);
    
    HIEFFPLA_INST_0_56992 : AOI1
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_1[0]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_1[1]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_1[2]\, Y => 
        HIEFFPLA_NET_0_116758);
    
    HIEFFPLA_INST_0_38642 : MX2
      port map(A => HIEFFPLA_NET_0_119524, B => 
        \U50_PATTERNS/ELINK_ADDRA_11[0]\, S => 
        HIEFFPLA_NET_0_119280, Y => HIEFFPLA_NET_0_120079);
    
    \U_ELK4_CH/U_SLAVE_1ELK/Q[14]\ : DFN1C0
      port map(D => \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[14]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/Q[14]_net_1\);
    
    \U_ELK9_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]\ : DFN1C0
      port map(D => \U_ELK9_CH/U_SLAVE_1ELK/Q[8]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]_net_1\);
    
    HIEFFPLA_INST_0_49381 : MX2
      port map(A => \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\, B
         => \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[13]_net_1\, S => 
        \BIT_OS_SEL[2]\, Y => HIEFFPLA_NET_0_118139);
    
    HIEFFPLA_INST_0_58050 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_0[1]\, B => 
        HIEFFPLA_NET_0_116677, S => HIEFFPLA_NET_0_117088, Y => 
        HIEFFPLA_NET_0_116571);
    
    \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[10]\ : DFN1C0
      port map(D => 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\);
    
    \U200A_TFC/GP_PG_SM[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120321, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_28, Q => 
        \U200A_TFC/GP_PG_SM[1]_net_1\);
    
    HIEFFPLA_INST_0_63054 : AND2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[9]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[10]\, Y => 
        HIEFFPLA_NET_0_115902);
    
    HIEFFPLA_INST_0_42902 : NAND3B
      port map(A => HIEFFPLA_NET_0_119438, B => 
        HIEFFPLA_NET_0_119372, C => HIEFFPLA_NET_0_119431, Y => 
        HIEFFPLA_NET_0_119428);
    
    \U_ELK12_CH/U_SLAVE_1ELK/Q[14]\ : DFN1C0
      port map(D => \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[14]_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/Q[14]_net_1\);
    
    HIEFFPLA_INST_0_37279 : AND2A
      port map(A => HIEFFPLA_NET_0_120307, B => \OP_MODE[0]\, Y
         => HIEFFPLA_NET_0_120308);
    
    \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[0]\ : DFN1C0
      port map(D => 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[0]_net_1\);
    
    \U50_PATTERNS/ELINK_RWA[6]/U1\ : DFN1P0
      port map(D => HIEFFPLA_NET_0_119695, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_6, Q => \U50_PATTERNS/ELINK_RWA[6]\);
    
    \U_MASTER_DES/U13A_ADJ_160M/BITCNT[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117695, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_14, Q => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[3]\);
    
    \U_ELK13_CH/U_SLAVE_1ELK/Q[1]\ : DFN1C0
      port map(D => \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/Q[1]_net_1\);
    
    \U50_PATTERNS/ELINK_DINA_14[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119828, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_16, Q => 
        \U50_PATTERNS/ELINK_DINA_14[3]\);
    
    HIEFFPLA_INST_0_51418 : NAND3A
      port map(A => HIEFFPLA_NET_0_117785, B => 
        \U_EXEC_MASTER/DEL_CNT[6]\, C => 
        \U_EXEC_MASTER/DEL_CNT[5]\, Y => HIEFFPLA_NET_0_117779);
    
    HIEFFPLA_INST_0_51186 : MX2
      port map(A => \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\, B
         => \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\, S => 
        \BIT_OS_SEL_2[2]\, Y => HIEFFPLA_NET_0_117815);
    
    HIEFFPLA_INST_0_49825 : MX2
      port map(A => 
        \U_ELK4_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]_net_1\, B => 
        \U_ELK4_CH/ELK_TX_DAT[2]\, S => 
        \U_ELK4_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118066);
    
    \U_ELK11_CH/U_SLAVE_1ELK/RECD_SER_WORD[2]\ : DFN1C0
      port map(D => \U_ELK11_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[2]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_11[2]\);
    
    HIEFFPLA_INST_0_42281 : AO1
      port map(A => \U50_PATTERNS/RD_USB_ADBUS[1]\, B => 
        \U50_PATTERNS/RD_USB_ADBUS[0]\, C => 
        HIEFFPLA_NET_0_119581, Y => HIEFFPLA_NET_0_119583);
    
    HIEFFPLA_INST_0_57290 : AND3B
      port map(A => HIEFFPLA_NET_0_117179, B => 
        HIEFFPLA_NET_0_116698, C => HIEFFPLA_NET_0_116714, Y => 
        HIEFFPLA_NET_0_116706);
    
    HIEFFPLA_INST_0_54888 : AND2A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_0[8]_net_1\, B => 
        HIEFFPLA_NET_0_115867, Y => HIEFFPLA_NET_0_117181);
    
    HIEFFPLA_INST_0_48616 : NAND2B
      port map(A => \OP_MODE_c_1[1]\, B => \PATT_ELK_DAT_18[1]\, 
        Y => HIEFFPLA_NET_0_118282);
    
    HIEFFPLA_INST_0_48310 : MX2
      port map(A => HIEFFPLA_NET_0_118355, B => 
        HIEFFPLA_NET_0_118338, S => \BIT_OS_SEL_3[1]\, Y => 
        HIEFFPLA_NET_0_118340);
    
    HIEFFPLA_INST_0_45775 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/SM_BANK_SEL[6]\, C => 
        \U50_PATTERNS/ELINK_DOUTA_13[7]\, Y => 
        HIEFFPLA_NET_0_118846);
    
    \U_ELK17_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]\ : DFN1C0
      port map(D => \U_ELK17_CH/U_SLAVE_1ELK/Q[9]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]_net_1\);
    
    HIEFFPLA_INST_0_46040 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_14[1]\, C => 
        \U50_PATTERNS/SM_BANK_SEL[5]\, Y => HIEFFPLA_NET_0_118780);
    
    HIEFFPLA_INST_0_53720 : AO1E
      port map(A => HIEFFPLA_NET_0_116678, B => 
        HIEFFPLA_NET_0_116593, C => HIEFFPLA_NET_0_117394, Y => 
        HIEFFPLA_NET_0_117366);
    
    \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[13]\ : DFN1C0
      port map(D => \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\, 
        CLK => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[13]_net_1\);
    
    \U_ELK8_CH/U_SLAVE_1ELK/RECD_SER_WORD[4]\ : DFN1C0
      port map(D => \U_ELK8_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[4]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_8[4]\);
    
    \U50_PATTERNS/ELINK_BLKA[11]/U1\ : DFN1P0
      port map(D => HIEFFPLA_NET_0_119933, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_20, Q => 
        \U50_PATTERNS/ELINK_BLKA[11]\);
    
    HIEFFPLA_INST_0_61328 : MX2
      port map(A => HIEFFPLA_NET_0_117186, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_21[3]\, S => 
        HIEFFPLA_NET_0_117144, Y => HIEFFPLA_NET_0_116142);
    
    HIEFFPLA_INST_0_52510 : MX2
      port map(A => HIEFFPLA_NET_0_117498, B => 
        HIEFFPLA_NET_0_117494, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_1[3]\, Y => 
        HIEFFPLA_NET_0_117554);
    
    \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[13]\ : DFN1C0
      port map(D => \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[13]_net_1\);
    
    \U_ELK4_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL\ : DFN1C0
      port map(D => 
        \U_ELK4_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL_net_1\);
    
    HIEFFPLA_INST_0_111824 : MX2B
      port map(A => 
        \U_EXEC_MASTER/USB_MASTER_EN/CNT_EN_60M2S_net_1\, B => 
        HIEFFPLA_NET_0_115827, S => HIEFFPLA_NET_0_117753, Y => 
        HIEFFPLA_NET_0_117741);
    
    \U_ELK5_CH/U_ELK1_SERDAT_SOURCE/SERDAT[5]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118008, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i, Q => 
        \U_ELK5_CH/ELK_TX_DAT[5]\);
    
    HIEFFPLA_INST_0_56820 : NAND3A
      port map(A => HIEFFPLA_NET_0_116801, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_0[6]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_0[7]\, Y => 
        HIEFFPLA_NET_0_116789);
    
    \U_ELK12_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U3\ : IOBI_ID_OD_EB
      port map(DR => \U_ELK12_CH/ELK_OUT_R\, DF => 
        \U_ELK12_CH/ELK_OUT_F\, CLR => \GND\, E => 
        \AFLSDF_INV_19\, ICLK => CCC_160M_ADJ, OCLK => 
        CCC_160M_FXD, YIN => 
        \U_ELK12_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\, DOUT => 
        OPEN, EOUT => 
        \U_ELK12_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET3\, YR => OPEN, 
        YF => OPEN);
    
    HIEFFPLA_INST_0_62003 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_12[2]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_28[2]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_3[4]_net_1\, Y
         => HIEFFPLA_NET_0_116048);
    
    HIEFFPLA_INST_0_54961 : AND3B
      port map(A => HIEFFPLA_NET_0_117246, B => 
        HIEFFPLA_NET_0_117241, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_3[6]_net_1\, Y => 
        HIEFFPLA_NET_0_117155);
    
    HIEFFPLA_INST_0_51250 : MX2
      port map(A => HIEFFPLA_NET_0_117818, B => 
        HIEFFPLA_NET_0_117814, S => \BIT_OS_SEL_4[0]\, Y => 
        \U_ELK9_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[3]\);
    
    HIEFFPLA_INST_0_63233 : MX2
      port map(A => \U_TFC_CMD_TX/SER_CMD_WORD_R[2]_net_1\, B => 
        \TFC_TX_DAT[7]\, S => \U_TFC_CMD_TX/START_RISE_net_1\, Y
         => \U_TFC_CMD_TX/N_SER_CMD_WORD_R[3]\);
    
    HIEFFPLA_INST_0_42831 : AND3A
      port map(A => \U50_PATTERNS/REG_STATE[1]_net_1\, B => 
        HIEFFPLA_NET_0_119370, C => 
        \U50_PATTERNS/REG_STATE[5]_net_1\, Y => 
        HIEFFPLA_NET_0_119454);
    
    \U200A_TFC/RX_SER_WORD_3DEL[5]\ : DFN1C0
      port map(D => \U200A_TFC/RX_SER_WORD_2DEL[5]_net_1\, CLK
         => CLK_40M_GL, CLR => P_MASTER_POR_B_c_24, Q => 
        \U200A_TFC/RX_SER_WORD_3DEL[5]_net_1\);
    
    HIEFFPLA_INST_0_38939 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_15[1]\, B => 
        HIEFFPLA_NET_0_119523, S => HIEFFPLA_NET_0_119297, Y => 
        HIEFFPLA_NET_0_120046);
    
    \P_CLK_40M_GL_pad/U0/U1\ : IOTRI_OB_EB
      port map(D => CLK_40M_GL, E => \VCC\, DOUT => 
        \P_CLK_40M_GL_pad/U0/NET1\, EOUT => 
        \P_CLK_40M_GL_pad/U0/NET2\);
    
    HIEFFPLA_INST_0_54133 : MX2
      port map(A => HIEFFPLA_NET_0_116171, B => 
        HIEFFPLA_NET_0_116065, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_1[3]_net_1\, Y
         => HIEFFPLA_NET_0_117304);
    
    \U_MASTER_DES/U13C_MASTER_DESER/ARB_WRD_40M_FIXED[1]\ : 
        DFN1C0
      port map(D => \U_MASTER_DES/U13C_MASTER_DESER/Q[1]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_26, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_WRD_40M_FIXED[1]_net_1\);
    
    \U_ELK4_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]\ : DFN1C0
      port map(D => \U_ELK4_CH/U_SLAVE_1ELK/Q[7]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]_net_1\);
    
    HIEFFPLA_INST_0_42872 : AND3A
      port map(A => HIEFFPLA_NET_0_119450, B => 
        \U50_PATTERNS/REG_STATE_0[1]_net_1\, C => 
        HIEFFPLA_NET_0_119411, Y => HIEFFPLA_NET_0_119440);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_15[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116517, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_15, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_15[3]\);
    
    HIEFFPLA_INST_0_45983 : NAND3C
      port map(A => HIEFFPLA_NET_0_118940, B => 
        HIEFFPLA_NET_0_118952, C => HIEFFPLA_NET_0_118697, Y => 
        HIEFFPLA_NET_0_118797);
    
    HIEFFPLA_INST_0_38466 : MX2
      port map(A => \U50_PATTERNS/ELINKS_STRT_ADDR_T[4]\, B => 
        \U50_PATTERNS/RD_USB_ADBUS[4]\, S => 
        HIEFFPLA_NET_0_119493, Y => HIEFFPLA_NET_0_120099);
    
    HIEFFPLA_INST_0_111287 : AND3A
      port map(A => HIEFFPLA_NET_0_115842, B => 
        HIEFFPLA_NET_0_116395, C => HIEFFPLA_NET_0_117404, Y => 
        HIEFFPLA_NET_0_116399);
    
    HIEFFPLA_INST_0_61892 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_11[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_27[1]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_2[4]_net_1\, Y
         => HIEFFPLA_NET_0_116064);
    
    HIEFFPLA_INST_0_42305 : AOI1
      port map(A => HIEFFPLA_NET_0_119583, B => 
        HIEFFPLA_NET_0_119580, C => HIEFFPLA_NET_0_119571, Y => 
        HIEFFPLA_NET_0_119577);
    
    HIEFFPLA_INST_0_42219 : AO1D
      port map(A => \U50_PATTERNS/RD_USB_ADBUS[5]\, B => 
        HIEFFPLA_NET_0_119565, C => 
        \U50_PATTERNS/RD_USB_ADBUS[6]\, Y => 
        HIEFFPLA_NET_0_119601);
    
    HIEFFPLA_INST_0_37572 : AND3
      port map(A => HIEFFPLA_NET_0_120257, B => \TFC_ADDRB[3]\, C
         => \TFC_ADDRB[2]\, Y => HIEFFPLA_NET_0_120258);
    
    \U_ELK15_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118421, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_6, Q => 
        \U_ELK15_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]_net_1\);
    
    \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[13]\ : DFN1C0
      port map(D => 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]_net_1\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[13]_net_1\);
    
    \U50_PATTERNS/ELINK_ADDRA_8[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119951, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_8, Q => 
        \U50_PATTERNS/ELINK_ADDRA_8[0]\);
    
    \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[1]\ : DFN1C0
      port map(D => 
        \U_ELK3_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\);
    
    \U_ELK14_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]\ : DFN1C0
      port map(D => \U_ELK14_CH/U_SLAVE_1ELK/Q[9]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_3[7]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116718, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_7, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_3[7]\);
    
    HIEFFPLA_INST_0_43047 : AND3A
      port map(A => HIEFFPLA_NET_0_119380, B => 
        HIEFFPLA_NET_0_119429, C => HIEFFPLA_NET_0_119393, Y => 
        HIEFFPLA_NET_0_119392);
    
    HIEFFPLA_INST_0_37459 : MX2
      port map(A => \U200A_TFC/LOC_STRT_ADDR[1]\, B => 
        \TFC_STRT_ADDR[1]\, S => \U200A_TFC/GP_PG_SM_0[10]_net_1\, 
        Y => HIEFFPLA_NET_0_120281);
    
    \U50_PATTERNS/ELINK_ADDRA_0[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120093, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_18, Q => 
        \U50_PATTERNS/ELINK_ADDRA_0[2]\);
    
    HIEFFPLA_INST_0_39945 : MX2
      port map(A => HIEFFPLA_NET_0_119913, B => 
        \U50_PATTERNS/ELINK_BLKA[10]\, S => 
        \U50_PATTERNS/SM_BANK_SEL[20]\, Y => 
        HIEFFPLA_NET_0_119934);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_16[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116511, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_16_0, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_16[1]\);
    
    \U_EXEC_MASTER/MPOR_SALT_B_13\ : DFI1P0
      port map(D => HIEFFPLA_NET_0_117781, CLK => CLK_40M_GL, PRE
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_2\, QN => 
        MASTER_SALT_POR_B_i_0_i_13);
    
    \U_ELK7_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL\ : DFN1C0
      port map(D => \U_ELK7_CH/ELK_IN_R_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL_net_1\);
    
    \U_ELK6_CH/U_SLAVE_1ELK/RECD_SER_WORD[0]\ : DFN1C0
      port map(D => \U_ELK6_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[0]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_6[0]\);
    
    HIEFFPLA_INST_0_57635 : NAND3C
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_5[8]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_5[7]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_5[6]\, Y => 
        HIEFFPLA_NET_0_116646);
    
    \U_ELK2_CH/U_SLAVE_1ELK/Q[7]\ : DFN1C0
      port map(D => \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/Q[7]_net_1\);
    
    \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[13]\ : DFN1C0
      port map(D => \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\, 
        CLK => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[13]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_10[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116559, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_6, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_10[3]\);
    
    HIEFFPLA_INST_0_63027 : AND3
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[12]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[8]\, C => 
        HIEFFPLA_NET_0_115909, Y => HIEFFPLA_NET_0_115910);
    
    HIEFFPLA_INST_0_51374 : MX2
      port map(A => HIEFFPLA_NET_0_117773, B => 
        \U_EXEC_MASTER/DEL_CNT[5]\, S => HIEFFPLA_NET_0_117796, Y
         => HIEFFPLA_NET_0_117790);
    
    \U_ELK8_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]\ : DFN1C0
      port map(D => \U_ELK8_CH/U_SLAVE_1ELK/Q[1]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]_net_1\);
    
    \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[13]\ : DFN1C0
      port map(D => 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[13]_net_1\);
    
    \U50_PATTERNS/ELINK_ADDRA_14[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120050, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_5, Q => 
        \U50_PATTERNS/ELINK_ADDRA_14[5]\);
    
    HIEFFPLA_INST_0_62863 : AOI1B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[8]_net_1\, B => 
        \OP_MODE_c[5]\, C => HIEFFPLA_NET_0_115938, Y => 
        HIEFFPLA_NET_0_115935);
    
    HIEFFPLA_INST_0_48113 : MX2
      port map(A => HIEFFPLA_NET_0_161286, B => 
        HIEFFPLA_NET_0_161285, S => HIEFFPLA_NET_0_161284, Y => 
        HIEFFPLA_NET_0_118375);
    
    HIEFFPLA_INST_0_56981 : AND3B
      port map(A => HIEFFPLA_NET_0_116756, B => 
        HIEFFPLA_NET_0_117179, C => HIEFFPLA_NET_0_116778, Y => 
        HIEFFPLA_NET_0_116760);
    
    HIEFFPLA_INST_0_50642 : MX2
      port map(A => \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[1]_net_1\, B
         => \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\, S => 
        \BIT_OS_SEL_4[2]\, Y => HIEFFPLA_NET_0_117912);
    
    \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[7]\ : DFN1C0
      port map(D => 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\);
    
    \U50_PATTERNS/U4B_REGCROSS/SAMP_TWO[0]\ : DFN1C0
      port map(D => \U50_PATTERNS/U4B_REGCROSS/SAMP_ONE[0]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_29, Q => 
        \U50_PATTERNS/U4B_REGCROSS/SAMP_TWO[0]_net_1\);
    
    HIEFFPLA_INST_0_56248 : AND2
      port map(A => DCB_SALT_SEL_c, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/RECD_SER_WORD[7]_net_1\, 
        Y => \ELK_RX_SER_WORD_0[7]\);
    
    \U_ELK8_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]\ : DFN1C0
      port map(D => \U_ELK8_CH/U_SLAVE_1ELK/Q[6]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]_net_1\);
    
    \U200B_ELINKS/RX_SER_WORD_3DEL[4]\ : DFN1C0
      port map(D => \U200B_ELINKS/RX_SER_WORD_2DEL[4]_net_1\, CLK
         => CLK_40M_GL, CLR => P_MASTER_POR_B_c_31_0, Q => 
        \U200B_ELINKS/RX_SER_WORD_3DEL[4]_net_1\);
    
    HIEFFPLA_INST_0_61172 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_1[1]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_2[1]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_1[0]\, Y => 
        HIEFFPLA_NET_0_116164);
    
    HIEFFPLA_INST_0_63020 : NAND3A
      port map(A => HIEFFPLA_NET_0_115916, B => 
        HIEFFPLA_NET_0_115902, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[11]\, Y => 
        HIEFFPLA_NET_0_115912);
    
    HIEFFPLA_INST_0_43632 : NAND2B
      port map(A => HIEFFPLA_NET_0_119270, B => 
        HIEFFPLA_NET_0_119279, Y => HIEFFPLA_NET_0_119261);
    
    HIEFFPLA_INST_0_51900 : MX2
      port map(A => HIEFFPLA_NET_0_117658, B => 
        HIEFFPLA_NET_0_117648, S => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[2]\, Y => 
        HIEFFPLA_NET_0_117669);
    
    HIEFFPLA_INST_0_47001 : MX2
      port map(A => HIEFFPLA_NET_0_118586, B => 
        HIEFFPLA_NET_0_118582, S => \BIT_OS_SEL[0]\, Y => 
        \U_ELK11_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[1]\);
    
    HIEFFPLA_INST_0_37554 : AND3
      port map(A => \TFC_ADDRB[1]\, B => HIEFFPLA_NET_0_120262, C
         => \TFC_ADDRB[2]\, Y => HIEFFPLA_NET_0_120261);
    
    \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[2]\ : DFN1C0
      port map(D => 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[2]_net_1\);
    
    HIEFFPLA_INST_0_47127 : AND2A
      port map(A => \OP_MODE_c_3[1]\, B => \PATT_ELK_DAT_12[6]\, 
        Y => HIEFFPLA_NET_0_118547);
    
    HIEFFPLA_INST_0_49617 : AND2A
      port map(A => \OP_MODE_c_5[1]\, B => \PATT_ELK_DAT_3[6]\, Y
         => HIEFFPLA_NET_0_118097);
    
    HIEFFPLA_INST_0_48592 : MX2
      port map(A => 
        \U_ELK18_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]_net_1\, B => 
        \U_ELK18_CH/ELK_TX_DAT[6]\, S => 
        \U_ELK18_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118289);
    
    \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[4]\ : DFN1C0
      port map(D => \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\);
    
    HIEFFPLA_INST_0_57103 : NAND2B
      port map(A => HIEFFPLA_NET_0_116708, B => 
        HIEFFPLA_NET_0_116740, Y => HIEFFPLA_NET_0_116742);
    
    \U50_PATTERNS/ELINK_DINA_17[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119807, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_19, Q => 
        \U50_PATTERNS/ELINK_DINA_17[0]\);
    
    HIEFFPLA_INST_0_43012 : AND3
      port map(A => HIEFFPLA_NET_0_119430, B => 
        HIEFFPLA_NET_0_119016, C => HIEFFPLA_NET_0_119379, Y => 
        HIEFFPLA_NET_0_119403);
    
    \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[8]\ : DFN1C0
      port map(D => 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\);
    
    \U50_PATTERNS/ELINK_DINA_1[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119781, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_7, Q => 
        \U50_PATTERNS/ELINK_DINA_1[2]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_17[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116202, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_7, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_17[3]\);
    
    \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[11]\ : DFN1C0
      port map(D => \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\);
    
    \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[4]\ : DFN1C0
      port map(D => \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117039, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_17_0, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[2]\);
    
    HIEFFPLA_INST_0_50115 : AND2A
      port map(A => \OP_MODE_c_5[1]\, B => \PATT_ELK_DAT_5[6]\, Y
         => HIEFFPLA_NET_0_118007);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_4[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116694, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_9, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_4[2]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_SEL_2[2]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_BIT_OS_VAL[2]\, CLK
         => CLK_40M_GL, CLR => P_MASTER_POR_B_c_27_1, Q => 
        \BIT_OS_SEL_2[2]\);
    
    HIEFFPLA_INST_0_112148 : OA1C
      port map(A => HIEFFPLA_NET_0_120234, B => 
        HIEFFPLA_NET_0_120190, C => HIEFFPLA_NET_0_115819, Y => 
        HIEFFPLA_NET_0_120219);
    
    \U_ELK6_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]\ : DFN1C0
      port map(D => \U_ELK6_CH/U_SLAVE_1ELK/Q[0]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]_net_1\);
    
    \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[12]\ : DFN1C0
      port map(D => \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\);
    
    HIEFFPLA_INST_0_44908 : AND3
      port map(A => \U50_PATTERNS/REG_STATE_0[1]_net_1\, B => 
        HIEFFPLA_NET_0_119561, C => HIEFFPLA_NET_0_119568, Y => 
        HIEFFPLA_NET_0_119023);
    
    \U200A_TFC/R_RWB/U1\ : DFN1P0
      port map(D => HIEFFPLA_NET_0_120263, CLK => CLK_40M_GL, PRE
         => P_MASTER_POR_B_c_16_0, Q => TFC_RWB);
    
    \U_EXEC_MASTER/MPOR_B_27_1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117787, CLK => CLK_40M_GL, CLR
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_0\, Q => 
        P_MASTER_POR_B_c_27_1);
    
    \U50_PATTERNS/U4E_REGCROSS/SAMP_ONE[4]\ : DFN1C0
      port map(D => \U50_PATTERNS/OP_MODE[4]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c, Q => 
        \U50_PATTERNS/U4E_REGCROSS/SAMP_ONE[4]_net_1\);
    
    HIEFFPLA_INST_0_63012 : NOR3B
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[4]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[2]\, C => 
        HIEFFPLA_NET_0_115914, Y => HIEFFPLA_NET_0_115915);
    
    \U50_PATTERNS/U4D_REGCROSS/DELCNT[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119092, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_26, Q => 
        \U50_PATTERNS/U4D_REGCROSS/DELCNT[0]_net_1\);
    
    HIEFFPLA_INST_0_45016 : AND3A
      port map(A => \U50_PATTERNS/USB_TXE_B\, B => 
        \U50_PATTERNS/REG_STATE_0[1]_net_1\, C => 
        \U50_PATTERNS/REG_STATE_0[5]_net_1\, Y => 
        HIEFFPLA_NET_0_118999);
    
    HIEFFPLA_INST_0_44795 : XOR2
      port map(A => \OP_MODE_c[5]\, B => 
        \U50_PATTERNS/U4E_REGCROSS/SAMP_TWO[5]_net_1\, Y => 
        HIEFFPLA_NET_0_119047);
    
    HIEFFPLA_INST_0_43581 : NAND2B
      port map(A => \U50_PATTERNS/SM_BANK_SEL[7]\, B => 
        \U50_PATTERNS/SM_BANK_SEL[3]\, Y => HIEFFPLA_NET_0_119281);
    
    HIEFFPLA_INST_0_39875 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_9[1]\, B => 
        HIEFFPLA_NET_0_119523, S => HIEFFPLA_NET_0_119292, Y => 
        HIEFFPLA_NET_0_119942);
    
    \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[13]\ : DFN1C0
      port map(D => 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]_net_1\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[13]_net_1\);
    
    \U50_PATTERNS/TFC_STOP_ADDR_T[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119179, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_15, Q => 
        \U50_PATTERNS/TFC_STOP_ADDR_T[1]\);
    
    HIEFFPLA_INST_0_52812 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_7[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_8[1]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_2[0]\, Y => 
        HIEFFPLA_NET_0_117507);
    
    HIEFFPLA_INST_0_46629 : AND2A
      port map(A => \OP_MODE_c_3[1]\, B => \PATT_ELK_DAT_10[6]\, 
        Y => HIEFFPLA_NET_0_118637);
    
    \U_ELK8_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]\ : DFN1C0
      port map(D => \U_ELK8_CH/U_SLAVE_1ELK/Q[0]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]_net_1\);
    
    \U_ELK2_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118153, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_8, Q => 
        \U_ELK2_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]_net_1\);
    
    HIEFFPLA_INST_0_47650 : MX2
      port map(A => \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[3]_net_1\, 
        B => \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\, S => 
        \BIT_OS_SEL_2[2]\, Y => HIEFFPLA_NET_0_118452);
    
    \U200A_TFC/ADDR_POINTER[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120366, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_30, Q => \TFC_ADDRB[1]\);
    
    \P_USB_TXE_B_pad/U0/U1\ : IOIN_IRP
      port map(PRE => \AFLSDF_INV_1\, ICLK => CLK60MHZ, YIN => 
        \P_USB_TXE_B_pad/U0/NET1\, Y => \U50_PATTERNS/USB_TXE_B\);
    
    HIEFFPLA_INST_0_56740 : AND3
      port map(A => HIEFFPLA_NET_0_117414, B => 
        HIEFFPLA_NET_0_117359, C => HIEFFPLA_NET_0_116813, Y => 
        HIEFFPLA_NET_0_116811);
    
    HIEFFPLA_INST_0_55930 : MX2
      port map(A => HIEFFPLA_NET_0_116987, B => 
        HIEFFPLA_NET_0_117003, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[2]\, Y => 
        HIEFFPLA_NET_0_116972);
    
    HIEFFPLA_INST_0_53331 : AND2
      port map(A => \BIT_OS_SEL[1]\, B => \BIT_OS_SEL[0]\, Y => 
        HIEFFPLA_NET_0_117427);
    
    HIEFFPLA_INST_0_47369 : AND2
      port map(A => CLK_40M_GL, B => 
        \U_ELK13_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0_net_1\, Y => 
        HIEFFPLA_NET_0_118509);
    
    HIEFFPLA_INST_0_37283 : AND2A
      port map(A => \OP_MODE[0]\, B => 
        \U200A_TFC/GP_PG_SM[6]_net_1\, Y => HIEFFPLA_NET_0_120306);
    
    \U_ELK6_CH/U_SLAVE_1ELK/Q[3]\ : DFN1C0
      port map(D => \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/Q[3]_net_1\);
    
    \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[10]\ : DFN1C0
      port map(D => 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]_net_1\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\);
    
    \U50_PATTERNS/ELINK_DINA_12[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119840, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_12, Q => 
        \U50_PATTERNS/ELINK_DINA_12[7]\);
    
    HIEFFPLA_INST_0_39973 : MX2
      port map(A => HIEFFPLA_NET_0_119905, B => 
        \U50_PATTERNS/ELINK_BLKA[14]\, S => 
        \U50_PATTERNS/SM_BANK_SEL[20]\, Y => 
        HIEFFPLA_NET_0_119930);
    
    AFLSDF_INV_32 : INV
      port map(A => DCB_SALT_SEL_c, Y => \AFLSDF_INV_32\);
    
    \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[12]\ : DFN1C0
      port map(D => 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]_net_1\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[12]_net_1\);
    
    \U50_PATTERNS/TFC_STRT_ADDR_T[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119159, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_4, Q => 
        \U50_PATTERNS/TFC_STRT_ADDR_T[5]\);
    
    HIEFFPLA_INST_0_53332 : AND2
      port map(A => \BIT_OS_SEL[2]\, B => \BIT_OS_SEL[0]\, Y => 
        HIEFFPLA_NET_0_117426);
    
    HIEFFPLA_INST_0_51721 : NAND2B
      port map(A => 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM_0[4]_net_1\, B => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[76]_net_1\, Y => 
        HIEFFPLA_NET_0_117705);
    
    HIEFFPLA_INST_0_49413 : MX2
      port map(A => HIEFFPLA_NET_0_118136, B => 
        HIEFFPLA_NET_0_118133, S => \BIT_OS_SEL[1]\, Y => 
        HIEFFPLA_NET_0_118134);
    
    \U_ELK19_CH/U_ELK1_CMD_TX/SER_OUT_FDEL\ : DFN1C0
      port map(D => \U_ELK19_CH/U_ELK1_CMD_TX/SER_OUT_FI_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_16, Q
         => \U_ELK19_CH/ELK_OUT_F\);
    
    \U_ELK8_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]\ : DFN1C0
      port map(D => \U_ELK8_CH/U_SLAVE_1ELK/Q[11]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]_net_1\);
    
    HIEFFPLA_INST_0_62230 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_31[1]\, B => 
        HIEFFPLA_NET_0_117167, S => HIEFFPLA_NET_0_117319, Y => 
        HIEFFPLA_NET_0_116019);
    
    AFLSDF_INV_2 : INV
      port map(A => EXT_INT_REF_SEL_c, Y => \AFLSDF_INV_2\);
    
    HIEFFPLA_INST_0_57261 : NAND3
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_3[0]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_3[2]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_3[1]\, Y => 
        HIEFFPLA_NET_0_116714);
    
    \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[1]\ : DFN1C0
      port map(D => 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[1]_net_1\);
    
    HIEFFPLA_INST_0_43225 : AO1D
      port map(A => HIEFFPLA_NET_0_119357, B => 
        HIEFFPLA_NET_0_119366, C => HIEFFPLA_NET_0_119356, Y => 
        HIEFFPLA_NET_0_119343);
    
    \U_ELK14_CH/U_SLAVE_1ELK/RECD_SER_WORD[6]\ : DFN1C0
      port map(D => \U_ELK14_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[6]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_14[6]\);
    
    HIEFFPLA_INST_0_60498 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_11[2]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_12[2]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_4[0]\, Y => 
        HIEFFPLA_NET_0_116258);
    
    HIEFFPLA_INST_0_56571 : AND3
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[9]_net_1\, B => 
        HIEFFPLA_NET_0_117426, C => HIEFFPLA_NET_0_117425, Y => 
        HIEFFPLA_NET_0_116836);
    
    HIEFFPLA_INST_0_115744 : AO18
      port map(A => HIEFFPLA_NET_0_115806, B => 
        \U200B_ELINKS/LOC_STOP_ADDR[1]\, C => \ELKS_ADDRB[1]\, Y
         => HIEFFPLA_NET_0_115809);
    
    \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[13]\ : DFN1C0
      port map(D => 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]_net_1\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[13]_net_1\);
    
    HIEFFPLA_INST_0_46253 : AO1
      port map(A => HIEFFPLA_NET_0_119476, B => 
        \U50_PATTERNS/CHKSUM[2]\, C => HIEFFPLA_NET_0_118903, Y
         => HIEFFPLA_NET_0_118731);
    
    AFLSDF_INV_8 : INV
      port map(A => P_USB_MASTER_EN_c_22, Y => \AFLSDF_INV_8\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_26[4]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116076, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_12, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_26[4]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_7[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116600, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_14, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_7[3]\);
    
    \U_ELK11_CH/U_SLAVE_1ELK/Q[6]\ : DFN1C0
      port map(D => \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/Q[6]_net_1\);
    
    HIEFFPLA_INST_0_50559 : MX2
      port map(A => \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[0]_net_1\, B
         => \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\, S => 
        \BIT_OS_SEL_5[2]\, Y => HIEFFPLA_NET_0_117934);
    
    HIEFFPLA_INST_0_41909 : AND2
      port map(A => HIEFFPLA_NET_0_119389, B => 
        \U50_PATTERNS/SM_BANK_SEL[10]\, Y => 
        HIEFFPLA_NET_0_119666);
    
    HIEFFPLA_INST_0_58745 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_19[0]\, B => 
        HIEFFPLA_NET_0_116680, S => HIEFFPLA_NET_0_117092, Y => 
        HIEFFPLA_NET_0_116481);
    
    HIEFFPLA_INST_0_41341 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_5[3]\, B => 
        HIEFFPLA_NET_0_119574, S => HIEFFPLA_NET_0_119251, Y => 
        HIEFFPLA_NET_0_119748);
    
    HIEFFPLA_INST_0_60693 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_14[3]\, B => 
        HIEFFPLA_NET_0_117186, S => HIEFFPLA_NET_0_117228, Y => 
        HIEFFPLA_NET_0_116232);
    
    \U50_PATTERNS/ELINK_DINA_13[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119832, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_14, Q => 
        \U50_PATTERNS/ELINK_DINA_13[7]\);
    
    \U_ELK11_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]\ : DFN1C0
      port map(D => \U_ELK11_CH/U_SLAVE_1ELK/Q[8]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]_net_1\);
    
    \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[5]\ : DFN1C0
      port map(D => 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\);
    
    HIEFFPLA_INST_0_38176 : MX2
      port map(A => \U50_PATTERNS/CHKSUM[3]\, B => 
        HIEFFPLA_NET_0_120132, S => HIEFFPLA_NET_0_119470, Y => 
        HIEFFPLA_NET_0_120140);
    
    \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[9]\ : DFN1C0
      port map(D => \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\);
    
    \U50_PATTERNS/ELINK_ADDRA_13[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120062, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_3, Q => 
        \U50_PATTERNS/ELINK_ADDRA_13[1]\);
    
    HIEFFPLA_INST_0_51941 : MX2A
      port map(A => HIEFFPLA_NET_0_117654, B => 
        HIEFFPLA_NET_0_117653, S => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[1]\, Y => 
        HIEFFPLA_NET_0_117661);
    
    HIEFFPLA_INST_0_38378 : MX2
      port map(A => \U50_PATTERNS/ELINKS_STRT_ADDR[1]\, B => 
        \U50_PATTERNS/ELINKS_STRT_ADDR_T[1]\, S => 
        HIEFFPLA_NET_0_119472, Y => HIEFFPLA_NET_0_120110);
    
    HIEFFPLA_INST_0_43563 : NAND2B
      port map(A => \U50_PATTERNS/SM_BANK_SEL[21]\, B => 
        \U50_PATTERNS/SM_BANK_SEL[11]\, Y => 
        HIEFFPLA_NET_0_119291);
    
    \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[1]\ : DFN1C0
      port map(D => 
        \U_ELK13_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\);
    
    \U50_PATTERNS/TFC_ADDRA[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119206, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_9, Q => \U50_PATTERNS/TFC_ADDRA[1]\);
    
    HIEFFPLA_INST_0_56774 : NAND2B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_0[8]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_0[7]\, Y => 
        HIEFFPLA_NET_0_116800);
    
    HIEFFPLA_INST_0_46872 : AND2A
      port map(A => \OP_MODE_c[1]\, B => \PATT_ELK_DAT_11[0]\, Y
         => HIEFFPLA_NET_0_118598);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_4[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_115999, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_13, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_4[1]\);
    
    HIEFFPLA_INST_0_46049 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_14[3]\, C => 
        \U50_PATTERNS/SM_BANK_SEL[5]\, Y => HIEFFPLA_NET_0_118778);
    
    \U_ELK1_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]\ : DFN1C0
      port map(D => \U_ELK1_CH/U_SLAVE_1ELK/Q[14]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]_net_1\);
    
    HIEFFPLA_INST_0_57183 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_3[1]\, B => 
        HIEFFPLA_NET_0_116707, S => HIEFFPLA_NET_0_117120, Y => 
        HIEFFPLA_NET_0_116724);
    
    HIEFFPLA_INST_0_48487 : MX2
      port map(A => HIEFFPLA_NET_0_118296, B => 
        HIEFFPLA_NET_0_118310, S => \BIT_OS_SEL_2[0]\, Y => 
        \U_ELK17_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[0]\);
    
    HIEFFPLA_INST_0_51266 : MX2
      port map(A => HIEFFPLA_NET_0_117813, B => 
        HIEFFPLA_NET_0_117823, S => \BIT_OS_SEL_4[0]\, Y => 
        \U_ELK9_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[5]\);
    
    AFLSDF_INV_60 : INV
      port map(A => \U200B_ELINKS/RX_SER_WORD_2DEL[3]_net_1\, Y
         => \AFLSDF_INV_60\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_6[4]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_115981, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_16, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_6[4]\);
    
    AFLSDF_INV_0 : INV
      port map(A => P_USB_MASTER_EN_c, Y => \AFLSDF_INV_0\);
    
    \U50_PATTERNS/ELINK_BLKA[16]/U1\ : DFN1P0
      port map(D => HIEFFPLA_NET_0_119928, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_20, Q => 
        \U50_PATTERNS/ELINK_BLKA[16]\);
    
    HIEFFPLA_INST_0_40171 : AOI1D
      port map(A => HIEFFPLA_NET_0_119389, B => 
        HIEFFPLA_NET_0_119464, C => 
        \U50_PATTERNS/SM_BANK_SEL[11]\, Y => 
        HIEFFPLA_NET_0_119881);
    
    \U_ELK18_CH/U_SLAVE_1ELK/Q[5]\ : DFN1C0
      port map(D => \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/Q[5]_net_1\);
    
    HIEFFPLA_INST_0_53452 : AND3A
      port map(A => HIEFFPLA_NET_0_116620, B => 
        HIEFFPLA_NET_0_117361, C => HIEFFPLA_NET_0_117414, Y => 
        HIEFFPLA_NET_0_117406);
    
    HIEFFPLA_INST_0_43665 : NAND3C
      port map(A => HIEFFPLA_NET_0_119279, B => 
        HIEFFPLA_NET_0_119229, C => HIEFFPLA_NET_0_119256, Y => 
        HIEFFPLA_NET_0_119248);
    
    HIEFFPLA_INST_0_42825 : AND3A
      port map(A => \U50_PATTERNS/REG_STATE[0]_net_1\, B => 
        \U50_PATTERNS/REG_STATE_0[5]_net_1\, C => 
        \U50_PATTERNS/REG_STATE_0[2]_net_1\, Y => 
        HIEFFPLA_NET_0_119455);
    
    \U200A_TFC/GP_PG_SM[8]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120311, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_28, Q => 
        \U200A_TFC/GP_PG_SM[8]_net_1\);
    
    HIEFFPLA_INST_0_43608 : NAND2B
      port map(A => \U50_PATTERNS/SM_BANK_SEL[18]\, B => 
        \U50_PATTERNS/SM_BANK_SEL[17]\, Y => 
        HIEFFPLA_NET_0_119269);
    
    \U_ELK16_CH/U_ELK1_SERDAT_SOURCE/SERDAT[6]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118367, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_9, Q => 
        \U_ELK16_CH/ELK_TX_DAT[6]\);
    
    HIEFFPLA_INST_0_49611 : AND2A
      port map(A => \OP_MODE_c_5[1]\, B => \PATT_ELK_DAT_3[0]\, Y
         => HIEFFPLA_NET_0_118103);
    
    \U_ELK6_CH/U_ELK1_SERDAT_SOURCE/SERDAT[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117968, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_1, Q => 
        \U_ELK6_CH/ELK_TX_DAT[0]\);
    
    \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[1]\ : DFN1C0
      port map(D => 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[1]_net_1\);
    
    HIEFFPLA_INST_0_40540 : MX2
      port map(A => HIEFFPLA_NET_0_119575, B => 
        \U50_PATTERNS/ELINK_DINA_13[2]\, S => 
        HIEFFPLA_NET_0_119285, Y => HIEFFPLA_NET_0_119837);
    
    \U_ELK13_CH/U_ELK1_SERDAT_SOURCE/SERDAT[5]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118503, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_4, Q => 
        \U_ELK13_CH/ELK_TX_DAT[5]\);
    
    \U50_PATTERNS/ELINK_DINA_3[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119760, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_11, Q => 
        \U50_PATTERNS/ELINK_DINA_3[7]\);
    
    \U50_PATTERNS/ELINK_ADDRA_1[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120007, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_20, Q => 
        \U50_PATTERNS/ELINK_ADDRA_1[0]\);
    
    HIEFFPLA_INST_0_59898 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_3[2]\, B => 
        HIEFFPLA_NET_0_116331, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_2[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116337);
    
    HIEFFPLA_INST_0_47872 : AND2A
      port map(A => \OP_MODE_c_6[1]\, B => \PATT_ELK_DAT_15[4]\, 
        Y => HIEFFPLA_NET_0_118414);
    
    HIEFFPLA_INST_0_50329 : MX2
      port map(A => 
        \U_ELK6_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]_net_1\, B => 
        \U_ELK6_CH/ELK_TX_DAT[4]\, S => 
        \U_ELK6_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_117975);
    
    HIEFFPLA_INST_0_43312 : NAND2A
      port map(A => HIEFFPLA_NET_0_119452, B => 
        HIEFFPLA_NET_0_119328, Y => HIEFFPLA_NET_0_119329);
    
    \U_ELK3_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL\ : DFN1C0
      port map(D => 
        \U_ELK3_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL_net_1\);
    
    \U_ELK13_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]\ : DFN1C0
      port map(D => \U_ELK13_CH/U_SLAVE_1ELK/Q[12]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]_net_1\);
    
    HIEFFPLA_INST_0_40315 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_10[1]\, B => 
        HIEFFPLA_NET_0_119576, S => HIEFFPLA_NET_0_119239, Y => 
        HIEFFPLA_NET_0_119862);
    
    HIEFFPLA_INST_0_57916 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_7[5]\, B => 
        HIEFFPLA_NET_0_116579, S => HIEFFPLA_NET_0_117113, Y => 
        HIEFFPLA_NET_0_116598);
    
    \U_ELK12_CH/U_SLAVE_1ELK/Q[5]\ : DFN1C0
      port map(D => \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/Q[5]_net_1\);
    
    \U50_PATTERNS/U4D_REGCROSS/SAMP_ONE[1]\ : DFN1C0
      port map(D => \U50_PATTERNS/ELINKS_STOP_ADDR[1]\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_25, Q => 
        \U50_PATTERNS/U4D_REGCROSS/SAMP_ONE[1]_net_1\);
    
    HIEFFPLA_INST_0_57524 : XA1B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_4[8]\, B => 
        HIEFFPLA_NET_0_116662, C => HIEFFPLA_NET_0_117179, Y => 
        HIEFFPLA_NET_0_116663);
    
    HIEFFPLA_INST_0_45901 : AO1
      port map(A => HIEFFPLA_NET_0_119254, B => 
        \U50_PATTERNS/ELINK_DOUTA_6[4]\, C => 
        HIEFFPLA_NET_0_118763, Y => HIEFFPLA_NET_0_118816);
    
    \U_ELK7_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117927, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_10, Q => 
        \U_ELK7_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]_net_1\);
    
    HIEFFPLA_INST_0_57193 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_3[2]\, B => 
        HIEFFPLA_NET_0_116706, S => HIEFFPLA_NET_0_117120, Y => 
        HIEFFPLA_NET_0_116723);
    
    \U_ELK11_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0\ : DFN1C0
      port map(D => CLK_40M_GL, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_5, Q => 
        \U_ELK11_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0_net_1\);
    
    HIEFFPLA_INST_0_62950 : MX2
      port map(A => HIEFFPLA_NET_0_115889, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[5]\, S => 
        HIEFFPLA_NET_0_117073, Y => HIEFFPLA_NET_0_115925);
    
    \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[13]\ : DFN1C0
      port map(D => \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[13]_net_1\);
    
    HIEFFPLA_INST_0_55307 : AND3B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[0]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[3]_net_1\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[2]_net_1\, Y => 
        HIEFFPLA_NET_0_117065);
    
    \U50_PATTERNS/ELINK_DINA_16[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119815, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_18, Q => 
        \U50_PATTERNS/ELINK_DINA_16[0]\);
    
    HIEFFPLA_INST_0_57483 : AND2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_4[5]\, B => 
        HIEFFPLA_NET_0_116684, Y => HIEFFPLA_NET_0_116672);
    
    \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[3]\ : DFN1C0
      port map(D => 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[3]_net_1\);
    
    HIEFFPLA_INST_0_54205 : MX2
      port map(A => HIEFFPLA_NET_0_116173, B => 
        HIEFFPLA_NET_0_116061, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_1[3]_net_1\, Y
         => HIEFFPLA_NET_0_117295);
    
    HIEFFPLA_INST_0_49724 : MX2
      port map(A => HIEFFPLA_NET_0_118092, B => 
        HIEFFPLA_NET_0_118089, S => \BIT_OS_SEL_6[1]\, Y => 
        HIEFFPLA_NET_0_118080);
    
    HIEFFPLA_INST_0_39605 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_5[3]\, B => 
        HIEFFPLA_NET_0_119520, S => HIEFFPLA_NET_0_119251, Y => 
        HIEFFPLA_NET_0_119972);
    
    HIEFFPLA_INST_0_39020 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_16[2]\, B => 
        HIEFFPLA_NET_0_119522, S => HIEFFPLA_NET_0_119257, Y => 
        HIEFFPLA_NET_0_120037);
    
    HIEFFPLA_INST_0_52266 : AND3A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[6]_net_1\, B => 
        HIEFFPLA_NET_0_117607, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[1]_net_1\, Y => 
        HIEFFPLA_NET_0_117597);
    
    \U_ELK3_CH/U_ELK1_SERDAT_SOURCE/SERDAT[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118101, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_15, Q => 
        \U_ELK3_CH/ELK_TX_DAT[2]\);
    
    \U50_PATTERNS/U105_PATT_ELINK_BLK/DPRT_512X9_SRAM_R0C0\ : 
        RAM4K9
      generic map(MEMORYFILE => "DPRT_512X9_SRAM_R0C0.mem")

      port map(ADDRA11 => AFLSDF_GND, ADDRA10 => AFLSDF_GND, 
        ADDRA9 => AFLSDF_GND, ADDRA8 => \GND\, ADDRA7 => 
        \U50_PATTERNS/ELINK_ADDRA_5[7]\, ADDRA6 => 
        \U50_PATTERNS/ELINK_ADDRA_5[6]\, ADDRA5 => 
        \U50_PATTERNS/ELINK_ADDRA_5[5]\, ADDRA4 => 
        \U50_PATTERNS/ELINK_ADDRA_5[4]\, ADDRA3 => 
        \U50_PATTERNS/ELINK_ADDRA_5[3]\, ADDRA2 => 
        \U50_PATTERNS/ELINK_ADDRA_5[2]\, ADDRA1 => 
        \U50_PATTERNS/ELINK_ADDRA_5[1]\, ADDRA0 => 
        \U50_PATTERNS/ELINK_ADDRA_5[0]\, ADDRB11 => AFLSDF_GND, 
        ADDRB10 => AFLSDF_GND, ADDRB9 => AFLSDF_GND, ADDRB8 => 
        \GND\, ADDRB7 => \ELKS_ADDRB[7]\, ADDRB6 => 
        \ELKS_ADDRB_0[6]\, ADDRB5 => \ELKS_ADDRB[5]\, ADDRB4 => 
        \ELKS_ADDRB_0[4]\, ADDRB3 => \ELKS_ADDRB[3]\, ADDRB2 => 
        \ELKS_ADDRB_0[2]\, ADDRB1 => \ELKS_ADDRB[1]\, ADDRB0 => 
        \ELKS_ADDRB[0]\, DINA8 => \GND\, DINA7 => 
        \U50_PATTERNS/ELINK_DINA_5[7]\, DINA6 => 
        \U50_PATTERNS/ELINK_DINA_5[6]\, DINA5 => 
        \U50_PATTERNS/ELINK_DINA_5[5]\, DINA4 => 
        \U50_PATTERNS/ELINK_DINA_5[4]\, DINA3 => 
        \U50_PATTERNS/ELINK_DINA_5[3]\, DINA2 => 
        \U50_PATTERNS/ELINK_DINA_5[2]\, DINA1 => 
        \U50_PATTERNS/ELINK_DINA_5[1]\, DINA0 => 
        \U50_PATTERNS/ELINK_DINA_5[0]\, DINB8 => \GND\, DINB7 => 
        \ELK_RX_SER_WORD_5[7]\, DINB6 => \ELK_RX_SER_WORD_5[6]\, 
        DINB5 => \ELK_RX_SER_WORD_5[5]\, DINB4 => 
        \ELK_RX_SER_WORD_5[4]\, DINB3 => \ELK_RX_SER_WORD_5[3]\, 
        DINB2 => \ELK_RX_SER_WORD_5[2]\, DINB1 => 
        \ELK_RX_SER_WORD_5[1]\, DINB0 => \ELK_RX_SER_WORD_5[0]\, 
        WIDTHA0 => \VCC\, WIDTHA1 => \VCC\, WIDTHB0 => \VCC\, 
        WIDTHB1 => \VCC\, PIPEA => \VCC\, PIPEB => \VCC\, WMODEA
         => \GND\, WMODEB => \GND\, BLKA => 
        \U50_PATTERNS/ELINK_BLKA[5]\, BLKB => ELKS_RAM_BLKB_EN, 
        WENA => \U50_PATTERNS/ELINK_RWA[5]\, WENB => ELKS_RWB, 
        CLKA => CLK60MHZ, CLKB => CLK_40M_GL, RESET => 
        P_USB_MASTER_EN_c_0, DOUTA8 => OPEN, DOUTA7 => 
        \U50_PATTERNS/ELINK_DOUTA_5[7]\, DOUTA6 => 
        \U50_PATTERNS/ELINK_DOUTA_5[6]\, DOUTA5 => 
        \U50_PATTERNS/ELINK_DOUTA_5[5]\, DOUTA4 => 
        \U50_PATTERNS/ELINK_DOUTA_5[4]\, DOUTA3 => 
        \U50_PATTERNS/ELINK_DOUTA_5[3]\, DOUTA2 => 
        \U50_PATTERNS/ELINK_DOUTA_5[2]\, DOUTA1 => 
        \U50_PATTERNS/ELINK_DOUTA_5[1]\, DOUTA0 => 
        \U50_PATTERNS/ELINK_DOUTA_5[0]\, DOUTB8 => OPEN, DOUTB7
         => \PATT_ELK_DAT_5[7]\, DOUTB6 => \PATT_ELK_DAT_5[6]\, 
        DOUTB5 => \PATT_ELK_DAT_5[5]\, DOUTB4 => 
        \PATT_ELK_DAT_5[4]\, DOUTB3 => \PATT_ELK_DAT_5[3]\, 
        DOUTB2 => \PATT_ELK_DAT_5[2]\, DOUTB1 => 
        \PATT_ELK_DAT_5[1]\, DOUTB0 => \PATT_ELK_DAT_5[0]\);
    
    HIEFFPLA_INST_0_60543 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_12[3]\, B => 
        HIEFFPLA_NET_0_117075, S => HIEFFPLA_NET_0_117133, Y => 
        HIEFFPLA_NET_0_116252);
    
    \U_EXEC_MASTER/PRESCALE[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117767, CLK => CLK_40M_GL, CLR
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i\, Q => 
        \U_EXEC_MASTER/PRESCALE[1]\);
    
    \U_ELK11_CH/U_SLAVE_1ELK/RECD_SER_WORD[1]\ : DFN1C0
      port map(D => \U_ELK11_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[1]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_11[1]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/Q[13]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[13]_net_1\, CLK => 
        CCC_160M_FXD, CLR => P_MASTER_POR_B_c_23, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/Q[13]_net_1\);
    
    \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[11]\ : DFN1C0
      port map(D => 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[11]_net_1\);
    
    HIEFFPLA_INST_0_57638 : NAND3A
      port map(A => HIEFFPLA_NET_0_116647, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_5[5]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_5[4]\, Y => 
        HIEFFPLA_NET_0_116645);
    
    HIEFFPLA_INST_0_52060 : MX2C
      port map(A => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[0]_net_1\, B => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[1]_net_1\, S => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[0]\, Y => 
        HIEFFPLA_NET_0_117644);
    
    HIEFFPLA_INST_0_56472 : AO1
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[4]_net_1\, B => 
        HIEFFPLA_NET_0_117428, C => HIEFFPLA_NET_0_116840, Y => 
        HIEFFPLA_NET_0_116856);
    
    \U50_PATTERNS/ELINKS_STRT_ADDR[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120107, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_17, Q => 
        \U50_PATTERNS/ELINKS_STRT_ADDR[4]\);
    
    HIEFFPLA_INST_0_62267 : AND2A
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[0]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_31[4]\, Y
         => HIEFFPLA_NET_0_116011);
    
    HIEFFPLA_INST_0_55214 : AND2B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[8]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[4]_net_1\, Y => 
        HIEFFPLA_NET_0_117087);
    
    HIEFFPLA_INST_0_42223 : NOR3A
      port map(A => HIEFFPLA_NET_0_119563, B => 
        \U50_PATTERNS/RD_USB_ADBUS[5]\, C => 
        \U50_PATTERNS/RD_USB_ADBUS[7]\, Y => 
        HIEFFPLA_NET_0_119600);
    
    \U_ELK16_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]\ : DFN1C0
      port map(D => \U_ELK16_CH/U_SLAVE_1ELK/Q[2]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]_net_1\);
    
    HIEFFPLA_INST_0_60459 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_11[2]\, B => 
        HIEFFPLA_NET_0_117131, S => HIEFFPLA_NET_0_117348, Y => 
        HIEFFPLA_NET_0_116263);
    
    HIEFFPLA_INST_0_55436 : AO1
      port map(A => HIEFFPLA_NET_0_117087, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[3]\, C => 
        HIEFFPLA_NET_0_117008, Y => HIEFFPLA_NET_0_117037);
    
    \U_TFC_CMD_TX/SER_OUT_FDEL\ : DFN1C0
      port map(D => \U_TFC_CMD_TX/SER_OUT_FI_net_1\, CLK => 
        CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        TFC_OUT_F);
    
    \U50_PATTERNS/ELINK_DINA_5[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119751, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_14, Q => 
        \U50_PATTERNS/ELINK_DINA_5[0]\);
    
    HIEFFPLA_INST_0_49323 : AND2
      port map(A => \U_ELK2_CH/ELK_TX_DAT[0]\, B => 
        \U_ELK2_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118157);
    
    HIEFFPLA_INST_0_47997 : MX2
      port map(A => HIEFFPLA_NET_0_118402, B => 
        HIEFFPLA_NET_0_118399, S => \BIT_OS_SEL_3[0]\, Y => 
        \U_ELK15_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[1]\);
    
    HIEFFPLA_INST_0_50800 : MX2
      port map(A => HIEFFPLA_NET_0_117902, B => 
        HIEFFPLA_NET_0_117888, S => \BIT_OS_SEL_6[1]\, Y => 
        HIEFFPLA_NET_0_117890);
    
    \U50_PATTERNS/U3_USB_DAT_BUS/_BIBUF_F_24U[4]_/U0/U1\ : 
        IOBI_IRC_OB_EB
      port map(D => \U50_PATTERNS/WR_USB_ADBUS[4]\, CLR => 
        \AFLSDF_INV_8\, E => \U50_PATTERNS/TrienAux\, ICLK => 
        CLK60MHZ, YIN => 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[4]\\\\/U0/NET3\, 
        DOUT => 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[4]\\\\/U0/NET1\, 
        EOUT => 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[4]\\\\/U0/NET2\, 
        Y => \U50_PATTERNS/RD_USB_ADBUS[4]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_115927, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_9, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[3]\);
    
    \U_ELK5_CH/U_SLAVE_1ELK/Q[13]\ : DFN1C0
      port map(D => \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[13]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/Q[13]_net_1\);
    
    HIEFFPLA_INST_0_51166 : MX2
      port map(A => HIEFFPLA_NET_0_117817, B => 
        HIEFFPLA_NET_0_117815, S => \BIT_OS_SEL_3[1]\, Y => 
        HIEFFPLA_NET_0_117818);
    
    HIEFFPLA_INST_0_50696 : MX2
      port map(A => \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\, B
         => \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\, S => 
        \BIT_OS_SEL_4[2]\, Y => HIEFFPLA_NET_0_117904);
    
    HIEFFPLA_INST_0_40387 : MX2
      port map(A => HIEFFPLA_NET_0_119576, B => 
        \U50_PATTERNS/ELINK_DINA_11[1]\, S => 
        HIEFFPLA_NET_0_119280, Y => HIEFFPLA_NET_0_119854);
    
    \U_ELK18_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0\ : DFN1C0
      port map(D => CLK_40M_GL, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_9, Q => 
        \U_ELK18_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0_net_1\);
    
    HIEFFPLA_INST_0_40151 : AOI1D
      port map(A => HIEFFPLA_NET_0_119389, B => 
        HIEFFPLA_NET_0_119464, C => 
        \U50_PATTERNS/SM_BANK_SEL[15]\, Y => 
        HIEFFPLA_NET_0_119889);
    
    \U50_PATTERNS/WR_XFER_TYPE[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118689, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c, Q => 
        \U50_PATTERNS/WR_XFER_TYPE[0]_net_1\);
    
    \U_ELK9_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117841, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_4, Q => 
        \U_ELK9_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]_net_1\);
    
    HIEFFPLA_INST_0_53624 : MX2
      port map(A => HIEFFPLA_NET_0_117363, B => 
        HIEFFPLA_NET_0_117398, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[1]_net_1\, Y
         => HIEFFPLA_NET_0_117381);
    
    HIEFFPLA_INST_0_45448 : AO1
      port map(A => HIEFFPLA_NET_0_119254, B => 
        \U50_PATTERNS/ELINK_DOUTA_6[1]\, C => 
        HIEFFPLA_NET_0_118819, Y => HIEFFPLA_NET_0_118912);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_11[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116551, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_8, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_11[3]\);
    
    \U_ELK12_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL\ : DFN1C0
      port map(D => \U_ELK12_CH/ELK_IN_R_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL_net_1\);
    
    HIEFFPLA_INST_0_37411 : MX2
      port map(A => \U200A_TFC/LOC_STOP_ADDR[1]\, B => 
        \TFC_STOP_ADDR[1]\, S => \U200A_TFC/GP_PG_SM_0[10]_net_1\, 
        Y => HIEFFPLA_NET_0_120289);
    
    HIEFFPLA_INST_0_55235 : AOI1D
      port map(A => HIEFFPLA_NET_0_117184, B => 
        HIEFFPLA_NET_0_117388, C => HIEFFPLA_NET_0_117213, Y => 
        HIEFFPLA_NET_0_117079);
    
    HIEFFPLA_INST_0_51001 : MX2
      port map(A => HIEFFPLA_NET_0_117865, B => 
        HIEFFPLA_NET_0_117860, S => \BIT_OS_SEL_5[0]\, Y => 
        \U_ELK8_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[3]\);
    
    \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[8]\ : DFN1C0
      port map(D => 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\);
    
    HIEFFPLA_INST_0_56365 : AO1
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[5]_net_1\, B => 
        HIEFFPLA_NET_0_117431, C => HIEFFPLA_NET_0_116861, Y => 
        HIEFFPLA_NET_0_116885);
    
    \U_ELK13_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]\ : DFN1C0
      port map(D => \U_ELK13_CH/U_SLAVE_1ELK/Q[6]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]_net_1\);
    
    \U50_PATTERNS/ELINK_ADDRA_1[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120002, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_20, Q => 
        \U50_PATTERNS/ELINK_ADDRA_1[5]\);
    
    HIEFFPLA_INST_0_41957 : AND3C
      port map(A => HIEFFPLA_NET_0_119265, B => 
        HIEFFPLA_NET_0_119261, C => 
        \U50_PATTERNS/SM_BANK_SEL[18]\, Y => 
        HIEFFPLA_NET_0_119646);
    
    \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[12]\ : DFN1C0
      port map(D => 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]_net_1\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[12]_net_1\);
    
    \U50_PATTERNS/ELINK_ADDRA_10[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120080, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_22, Q => 
        \U50_PATTERNS/ELINK_ADDRA_10[7]\);
    
    \U_EXEC_MASTER/USB_MASTER_EN/CNT_EN_60M2S\ : DFN1C0
      port map(D => 
        \U_EXEC_MASTER/USB_MASTER_EN/CNT_EN_60M1S_net_1\, CLK => 
        CLK60MHZ, CLR => P_MASTER_POR_B_c_23, Q => 
        \U_EXEC_MASTER/USB_MASTER_EN/CNT_EN_60M2S_net_1\);
    
    HIEFFPLA_INST_0_38490 : MX2
      port map(A => \U50_PATTERNS/ELINKS_STRT_ADDR_T[7]\, B => 
        \U50_PATTERNS/RD_USB_ADBUS[7]\, S => 
        HIEFFPLA_NET_0_119493, Y => HIEFFPLA_NET_0_120096);
    
    HIEFFPLA_INST_0_44888 : AO1
      port map(A => HIEFFPLA_NET_0_119015, B => 
        HIEFFPLA_NET_0_119456, C => HIEFFPLA_NET_0_119031, Y => 
        HIEFFPLA_NET_0_119027);
    
    ELK0_IN_R : DFN1C0
      port map(D => \AFLSDF_INV_62\, CLK => CCC_160M_ADJ, CLR => 
        DEV_RST_B_c, Q => \ELK0_IN_R\);
    
    \U_ELK10_CH/U_ELK1_CMD_TX/SER_OUT_RI\ : DFN1C0
      port map(D => 
        \U_ELK10_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_11, Q
         => \U_ELK10_CH/U_ELK1_CMD_TX/SER_OUT_RI_net_1\);
    
    \U50_PATTERNS/SI_CNT[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119333, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_5, Q => \U50_PATTERNS/SI_CNT[1]\);
    
    HIEFFPLA_INST_0_48409 : MX2
      port map(A => HIEFFPLA_NET_0_118316, B => 
        HIEFFPLA_NET_0_118312, S => \BIT_OS_SEL_1[1]\, Y => 
        HIEFFPLA_NET_0_118315);
    
    \U_EXEC_MASTER/MPOR_B_33\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117787, CLK => CLK_40M_GL, CLR
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_0\, Q => 
        P_MASTER_POR_B_c_33);
    
    HIEFFPLA_INST_0_111892 : NAND3C
      port map(A => HIEFFPLA_NET_0_115826, B => 
        HIEFFPLA_NET_0_118744, C => HIEFFPLA_NET_0_118753, Y => 
        HIEFFPLA_NET_0_118965);
    
    \U50_PATTERNS/WR_XFER_TYPE[4]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118685, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c, Q => 
        \U50_PATTERNS/WR_XFER_TYPE[4]_net_1\);
    
    HIEFFPLA_INST_0_47266 : MX2
      port map(A => HIEFFPLA_NET_0_118534, B => 
        HIEFFPLA_NET_0_118545, S => \BIT_OS_SEL_5[0]\, Y => 
        \U_ELK12_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[3]\);
    
    \U_ELK12_CH/U_ELK1_SERDAT_SOURCE/SERDAT[5]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118548, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_2, Q => 
        \U_ELK12_CH/ELK_TX_DAT[5]\);
    
    \U_ELK9_CH/U_SLAVE_1ELK/Q[3]\ : DFN1C0
      port map(D => \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/Q[3]_net_1\);
    
    HIEFFPLA_INST_0_42650 : AND3A
      port map(A => \U50_PATTERNS/REG_STATE_0[4]_net_1\, B => 
        HIEFFPLA_NET_0_119367, C => HIEFFPLA_NET_0_119021, Y => 
        HIEFFPLA_NET_0_119491);
    
    \U_ELK12_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]\ : DFN1C0
      port map(D => \U_ELK12_CH/U_SLAVE_1ELK/Q[12]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]_net_1\);
    
    \U_ELK11_CH/U_SLAVE_1ELK/Q[13]\ : DFN1C0
      port map(D => \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[13]_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/Q[13]_net_1\);
    
    \U_ELK12_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]\ : DFN1C0
      port map(D => \U_ELK12_CH/U_SLAVE_1ELK/Q[0]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]_net_1\);
    
    HIEFFPLA_INST_0_51356 : MX2
      port map(A => HIEFFPLA_NET_0_117775, B => 
        \U_EXEC_MASTER/DEL_CNT[3]\, S => HIEFFPLA_NET_0_117796, Y
         => HIEFFPLA_NET_0_117792);
    
    HIEFFPLA_INST_0_44533 : XO1
      port map(A => \ELKS_STRT_ADDR[5]\, B => 
        \U50_PATTERNS/U4C_REGCROSS/SAMP_TWO[5]_net_1\, C => 
        HIEFFPLA_NET_0_119099, Y => HIEFFPLA_NET_0_119100);
    
    HIEFFPLA_INST_0_42840 : AND3C
      port map(A => \U50_PATTERNS/REG_STATE[2]_net_1\, B => 
        \U50_PATTERNS/REG_STATE[0]_net_1\, C => 
        HIEFFPLA_NET_0_119436, Y => HIEFFPLA_NET_0_119452);
    
    \U50_PATTERNS/U4B_REGCROSS/LOCAL_REG_VAL[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119129, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_19, Q => \TFC_STOP_ADDR[4]\);
    
    HIEFFPLA_INST_0_37675 : AND3C
      port map(A => \U200B_ELINKS/GP_PG_SM[6]_net_1\, B => 
        \U200B_ELINKS/GP_PG_SM[7]_net_1\, C => 
        \U200B_ELINKS/GP_PG_SM[8]_net_1\, Y => 
        HIEFFPLA_NET_0_120233);
    
    \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[14]\ : DFN1C0
      port map(D => 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]_net_1\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[14]_net_1\);
    
    HIEFFPLA_INST_0_55528 : MX2
      port map(A => HIEFFPLA_NET_0_117024, B => 
        HIEFFPLA_NET_0_117012, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[2]\, Y => 
        HIEFFPLA_NET_0_117025);
    
    HIEFFPLA_INST_0_39731 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_7[1]\, B => 
        HIEFFPLA_NET_0_119523, S => HIEFFPLA_NET_0_119289, Y => 
        HIEFFPLA_NET_0_119958);
    
    \U_ELK14_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U0\ : IOPADP_BI
      port map(N2PIN => 
        \U_ELK14_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2_N2P\, D => 
        \U_ELK14_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, E => 
        \U_ELK14_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET2\, PAD => 
        ELK14_DAT_P, Y => 
        \U_ELK14_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\);
    
    \U50_PATTERNS/U4E_REGCROSS/SAMP_TWO[5]\ : DFN1C0
      port map(D => \U50_PATTERNS/U4E_REGCROSS/SAMP_ONE[5]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_24, Q => 
        \U50_PATTERNS/U4E_REGCROSS/SAMP_TWO[5]_net_1\);
    
    HIEFFPLA_INST_0_42344 : AND2A
      port map(A => \U50_PATTERNS/RD_USB_ADBUS[1]\, B => 
        \U50_PATTERNS/RD_USB_ADBUS[0]\, Y => 
        HIEFFPLA_NET_0_119563);
    
    HIEFFPLA_INST_0_51696 : MX2
      port map(A => \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[49]\, B
         => \U_MASTER_DES/PHASE_ADJ_160_L[3]\, S => 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM_0[4]_net_1\, Y => 
        HIEFFPLA_NET_0_117723);
    
    \U_EXEC_MASTER/MPOR_B_20\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117787, CLK => CLK_40M_GL, CLR
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_1\, Q => 
        P_MASTER_POR_B_c_20);
    
    HIEFFPLA_INST_0_59088 : MX2
      port map(A => HIEFFPLA_NET_0_116687, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_23[2]\, S => 
        HIEFFPLA_NET_0_117214, Y => HIEFFPLA_NET_0_116436);
    
    \U_ELK4_CH/U_SLAVE_1ELK/Q[3]\ : DFN1C0
      port map(D => \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/Q[3]_net_1\);
    
    HIEFFPLA_INST_0_56825 : AXOI4
      port map(A => HIEFFPLA_NET_0_117085, B => 
        HIEFFPLA_NET_0_117600, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_1[0]\, Y => 
        HIEFFPLA_NET_0_116788);
    
    HIEFFPLA_INST_0_43727 : NAND3C
      port map(A => HIEFFPLA_NET_0_119282, B => 
        HIEFFPLA_NET_0_119261, C => 
        \U50_PATTERNS/SM_BANK_SEL[19]\, Y => 
        HIEFFPLA_NET_0_119230);
    
    \U_ELK13_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]\ : DFN1C0
      port map(D => \U_ELK13_CH/U_SLAVE_1ELK/Q[14]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]_net_1\);
    
    HIEFFPLA_INST_0_52306 : NAND3A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[7]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[5]_net_1\, C => 
        HIEFFPLA_NET_0_117605, Y => HIEFFPLA_NET_0_117585);
    
    HIEFFPLA_INST_0_52180 : MX2
      port map(A => \U_MASTER_DES/AUX_SSHIFT\, B => 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM[2]_net_1\, S => 
        HIEFFPLA_NET_0_117628, Y => HIEFFPLA_NET_0_117615);
    
    \U_ELK15_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]\ : DFN1C0
      port map(D => \U_ELK15_CH/U_SLAVE_1ELK/Q[12]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]_net_1\);
    
    \U200B_ELINKS/GP_PG_SM[10]\ : DFN1P0
      port map(D => HIEFFPLA_NET_0_120227, CLK => CLK_40M_GL, PRE
         => P_MASTER_POR_B_c_34_0, Q => 
        \U200B_ELINKS/GP_PG_SM[10]_net_1\);
    
    \U_ELK15_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]\ : DFN1C0
      port map(D => \U_ELK15_CH/U_SLAVE_1ELK/Q[0]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]_net_1\);
    
    HIEFFPLA_INST_0_49401 : MX2
      port map(A => \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[3]_net_1\, B
         => \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\, S => 
        \BIT_OS_SEL_7[2]\, Y => HIEFFPLA_NET_0_118136);
    
    HIEFFPLA_INST_0_53703 : NAND3A
      port map(A => HIEFFPLA_NET_0_117390, B => 
        HIEFFPLA_NET_0_117325, C => HIEFFPLA_NET_0_116589, Y => 
        HIEFFPLA_NET_0_117369);
    
    HIEFFPLA_INST_0_62484 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_6[2]\, 
        B => HIEFFPLA_NET_0_117131, S => HIEFFPLA_NET_0_117132, Y
         => HIEFFPLA_NET_0_115983);
    
    HIEFFPLA_INST_0_53911 : AND3B
      port map(A => HIEFFPLA_NET_0_117390, B => 
        HIEFFPLA_NET_0_117392, C => HIEFFPLA_NET_0_117391, Y => 
        HIEFFPLA_NET_0_117334);
    
    HIEFFPLA_INST_0_49576 : MX2
      port map(A => 
        \U_ELK3_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]_net_1\, B => 
        \U_ELK3_CH/ELK_TX_DAT[2]\, S => 
        \U_ELK3_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118111);
    
    \U50_PATTERNS/TFC_ADDRA[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119205, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_9, Q => \U50_PATTERNS/TFC_ADDRA[2]\);
    
    HIEFFPLA_INST_0_61655 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_8[4]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_24[4]\, S
         => \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_4[4]_net_1\, 
        Y => HIEFFPLA_NET_0_116096);
    
    \U50_PATTERNS/CHKSUM[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120143, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_3, Q => \U50_PATTERNS/CHKSUM[0]\);
    
    HIEFFPLA_INST_0_40130 : AO1A
      port map(A => HIEFFPLA_NET_0_119872, B => 
        HIEFFPLA_NET_0_119240, C => HIEFFPLA_NET_0_119232, Y => 
        HIEFFPLA_NET_0_119897);
    
    \U50_PATTERNS/ELINK_DINA_7[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119730, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_17, Q => 
        \U50_PATTERNS/ELINK_DINA_7[5]\);
    
    HIEFFPLA_INST_0_51973 : MX2
      port map(A => HIEFFPLA_NET_0_117641, B => 
        HIEFFPLA_NET_0_117636, S => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[3]\, Y => 
        HIEFFPLA_NET_0_117658);
    
    HIEFFPLA_INST_0_44429 : XO1
      port map(A => \TFC_STOP_ADDR[5]\, B => 
        \U50_PATTERNS/U4B_REGCROSS/SAMP_TWO[5]_net_1\, C => 
        HIEFFPLA_NET_0_119120, Y => HIEFFPLA_NET_0_119121);
    
    HIEFFPLA_INST_0_59214 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_25[0]\, B => 
        HIEFFPLA_NET_0_116416, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_2[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116420);
    
    HIEFFPLA_INST_0_54902 : AOI1C
      port map(A => HIEFFPLA_NET_0_117184, B => 
        HIEFFPLA_NET_0_117388, C => HIEFFPLA_NET_0_117206, Y => 
        HIEFFPLA_NET_0_117175);
    
    HIEFFPLA_INST_0_44448 : MX2
      port map(A => \ELKS_STRT_ADDR[0]\, B => 
        \U50_PATTERNS/U4C_REGCROSS/SAMP_TWO[0]_net_1\, S => 
        HIEFFPLA_NET_0_119114, Y => HIEFFPLA_NET_0_119112);
    
    HIEFFPLA_INST_0_59480 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_11[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_27[1]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_5[4]_net_1\, Y
         => HIEFFPLA_NET_0_116389);
    
    \U50_PATTERNS/ELINK_ADDRA_11[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120077, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_2, Q => 
        \U50_PATTERNS/ELINK_ADDRA_11[2]\);
    
    HIEFFPLA_INST_0_60798 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_15[0]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_16[0]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[0]\, Y => 
        HIEFFPLA_NET_0_116218);
    
    HIEFFPLA_INST_0_52728 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_25[3]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_26[3]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_3[0]\, Y => 
        HIEFFPLA_NET_0_117521);
    
    \U50_PATTERNS/ELINK_ADDRA_8[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119944, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_8, Q => 
        \U50_PATTERNS/ELINK_ADDRA_8[7]\);
    
    HIEFFPLA_INST_0_56267 : NAND3C
      port map(A => HIEFFPLA_NET_0_116879, B => 
        HIEFFPLA_NET_0_116887, C => HIEFFPLA_NET_0_116895, Y => 
        HIEFFPLA_NET_0_116903);
    
    \U_ELK0_CMD_TX/SER_OUT_RI\ : DFI1C0
      port map(D => \U_ELK0_CMD_TX/SER_CMD_WORD_R[3]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_14, QN
         => \U_ELK0_CMD_TX/SER_OUT_RI_i\);
    
    HIEFFPLA_INST_0_37091 : AND2A
      port map(A => \TFC_STRT_ADDR[7]\, B => 
        HIEFFPLA_NET_0_120349, Y => HIEFFPLA_NET_0_120350);
    
    \U_ELK13_CH/U_SLAVE_1ELK/Q[7]\ : DFN1C0
      port map(D => \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/Q[7]_net_1\);
    
    \U50_PATTERNS/ELINK_ADDRA_1[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120000, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_20, Q => 
        \U50_PATTERNS/ELINK_ADDRA_1[7]\);
    
    \U50_PATTERNS/ELINK_ADDRA_6[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119964, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_4, Q => 
        \U50_PATTERNS/ELINK_ADDRA_6[3]\);
    
    \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[12]\ : DFN1C0
      port map(D => 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[12]_net_1\);
    
    \U50_PATTERNS/ELINK_ADDRA_0[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120095, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_18, Q => 
        \U50_PATTERNS/ELINK_ADDRA_0[0]\);
    
    HIEFFPLA_INST_0_49172 : MX2
      port map(A => \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\, B
         => \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\, S => 
        \BIT_OS_SEL[2]\, Y => HIEFFPLA_NET_0_118178);
    
    HIEFFPLA_INST_0_37835 : AND3
      port map(A => \U200B_ELINKS/GP_PG_SM[4]_net_1\, B => 
        HIEFFPLA_NET_0_120222, C => HIEFFPLA_NET_0_120190, Y => 
        HIEFFPLA_NET_0_120194);
    
    \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[3]\ : DFN1C0
      port map(D => \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\);
    
    HIEFFPLA_INST_0_57441 : AND3
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_4[5]\, B => 
        HIEFFPLA_NET_0_116684, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_4[6]\, Y => 
        HIEFFPLA_NET_0_116682);
    
    \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[6]\ : DFN1C0
      port map(D => 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\);
    
    \U50_PATTERNS/REG_STATE_0[5]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119008, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_22_0, Q => 
        \U50_PATTERNS/REG_STATE_0[5]_net_1\);
    
    \U200A_TFC/LOC_STOP_ADDR[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120288, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_1, Q => \U200A_TFC/LOC_STOP_ADDR[2]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/PHASE_ADJ[2]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[2]_net_1\, CLK
         => CLK_40M_GL, CLR => P_MASTER_POR_B_c, Q => 
        \U_MASTER_DES/PHASE_ADJ_160_L[2]\);
    
    \U_ELK15_CH/U_ELK1_SERDAT_SOURCE/SERDAT[5]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118413, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_8, Q => 
        \U_ELK15_CH/ELK_TX_DAT[5]\);
    
    \U50_PATTERNS/ELINK_DINA_4[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119758, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_12, Q => 
        \U50_PATTERNS/ELINK_DINA_4[1]\);
    
    \U50_PATTERNS/ELINK_ADDRA_8[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119947, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_8, Q => 
        \U50_PATTERNS/ELINK_ADDRA_8[4]\);
    
    HIEFFPLA_INST_0_49369 : NAND2B
      port map(A => \OP_MODE_c_1[1]\, B => \PATT_ELK_DAT_2[7]\, Y
         => HIEFFPLA_NET_0_118141);
    
    HIEFFPLA_INST_0_55371 : AND3
      port map(A => HIEFFPLA_NET_0_115906, B => 
        \U_MASTER_DES/CCC_RX_CLK_LOCK\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[3]_net_1\, Y => 
        HIEFFPLA_NET_0_117047);
    
    HIEFFPLA_INST_0_38450 : MX2
      port map(A => \U50_PATTERNS/ELINKS_STRT_ADDR_T[2]\, B => 
        \U50_PATTERNS/RD_USB_ADBUS[2]\, S => 
        HIEFFPLA_NET_0_119493, Y => HIEFFPLA_NET_0_120101);
    
    HIEFFPLA_INST_0_40900 : MX2
      port map(A => HIEFFPLA_NET_0_119575, B => 
        \U50_PATTERNS/ELINK_DINA_18[2]\, S => 
        HIEFFPLA_NET_0_119264, Y => HIEFFPLA_NET_0_119797);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_3[8]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116717, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_7, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_3[8]\);
    
    \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[6]\ : DFN1C0
      port map(D => \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_29[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116375, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_4, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_29[3]\);
    
    \U_ELK11_CH/U_SLAVE_1ELK/Q[5]\ : DFN1C0
      port map(D => \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/Q[5]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[10]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[8]_net_1\, CLK => 
        CCC_160M_ADJ, CLR => P_MASTER_POR_B_c_26, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[10]_net_1\);
    
    \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[12]\ : DFN1C0
      port map(D => 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[12]_net_1\);
    
    HIEFFPLA_INST_0_38012 : MX2
      port map(A => \U200B_ELINKS/LOC_STRT_ADDR[5]\, B => 
        \ELKS_STRT_ADDR[5]\, S => 
        \U200B_ELINKS/GP_PG_SM_0[10]_net_1\, Y => 
        HIEFFPLA_NET_0_120174);
    
    \U_ELK13_CH/U_ELK1_SERDAT_SOURCE/SERDAT[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118507, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_4, Q => 
        \U_ELK13_CH/ELK_TX_DAT[1]\);
    
    HIEFFPLA_INST_0_48883 : MX2
      port map(A => \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\, 
        B => \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\, S => 
        \BIT_OS_SEL[2]\, Y => HIEFFPLA_NET_0_118229);
    
    \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_SEL_0[0]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_BIT_OS_VAL[0]\, CLK
         => CLK_40M_GL, CLR => P_MASTER_POR_B_c_27_0, Q => 
        \BIT_OS_SEL_0[0]\);
    
    \U200A_TFC/LOC_DIR_MODE/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120292, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_15, Q => \U200A_TFC/N_232_li\);
    
    \U200B_ELINKS/LOC_STRT_ADDR[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120176, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_11, Q => 
        \U200B_ELINKS/LOC_STRT_ADDR[3]\);
    
    HIEFFPLA_INST_0_60504 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_11[3]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_12[3]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_4[0]\, Y => 
        HIEFFPLA_NET_0_116257);
    
    HIEFFPLA_INST_0_54967 : OR2A
      port map(A => HIEFFPLA_NET_0_117115, B => 
        HIEFFPLA_NET_0_117152, Y => HIEFFPLA_NET_0_117153);
    
    HIEFFPLA_INST_0_50168 : MX2
      port map(A => \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\, B
         => \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\, S => 
        \BIT_OS_SEL_6[2]\, Y => HIEFFPLA_NET_0_117998);
    
    HIEFFPLA_INST_0_47125 : AND2A
      port map(A => \OP_MODE_c_3[1]\, B => \PATT_ELK_DAT_12[4]\, 
        Y => HIEFFPLA_NET_0_118549);
    
    \U_ELK15_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118420, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_6, Q => 
        \U_ELK15_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]_net_1\);
    
    HIEFFPLA_INST_0_61271 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_4[0]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_20[0]\, S
         => \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_5[4]_net_1\, 
        Y => HIEFFPLA_NET_0_116150);
    
    HIEFFPLA_INST_0_62436 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_5[3]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_6[3]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_2[0]\, Y => 
        HIEFFPLA_NET_0_115990);
    
    HIEFFPLA_INST_0_62271 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_3[0]\, 
        B => HIEFFPLA_NET_0_117096, S => HIEFFPLA_NET_0_117178, Y
         => HIEFFPLA_NET_0_116010);
    
    HIEFFPLA_INST_0_51788 : MX2
      port map(A => \U_MASTER_DES/U13A_ADJ_160M/BITCNT[6]\, B => 
        HIEFFPLA_NET_0_117676, S => HIEFFPLA_NET_0_117630, Y => 
        HIEFFPLA_NET_0_117692);
    
    HIEFFPLA_INST_0_39119 : MX2
      port map(A => HIEFFPLA_NET_0_119518, B => 
        \U50_PATTERNS/ELINK_ADDRA_17[5]\, S => 
        HIEFFPLA_NET_0_119260, Y => HIEFFPLA_NET_0_120026);
    
    HIEFFPLA_INST_0_111912 : AOI1D
      port map(A => HIEFFPLA_NET_0_118692, B => 
        \U50_PATTERNS/WR_XFER_TYPE[1]_net_1\, C => 
        \U50_PATTERNS/ELK_N_ACTIVE_net_1\, Y => 
        HIEFFPLA_NET_0_115822);
    
    \U50_PATTERNS/U4E_REGCROSS/SAMP_TWO[1]\ : DFN1C0
      port map(D => \U50_PATTERNS/U4E_REGCROSS/SAMP_ONE[1]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_23, Q => 
        \U50_PATTERNS/U4E_REGCROSS/SAMP_TWO[1]_net_1\);
    
    HIEFFPLA_INST_0_51726 : NAND2B
      port map(A => 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM[4]_net_1\, B => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[8]_net_1\, Y => 
        HIEFFPLA_NET_0_117700);
    
    HIEFFPLA_INST_0_50110 : NAND2B
      port map(A => \OP_MODE_c_4[1]\, B => \PATT_ELK_DAT_5[1]\, Y
         => HIEFFPLA_NET_0_118012);
    
    \U_ELK17_CH/U_ELK1_SERDAT_SOURCE/SERDAT[7]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118321, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_12, Q => 
        \U_ELK17_CH/ELK_TX_DAT[7]\);
    
    HIEFFPLA_INST_0_46311 : NAND3B
      port map(A => HIEFFPLA_NET_0_118885, B => 
        HIEFFPLA_NET_0_118867, C => HIEFFPLA_NET_0_119427, Y => 
        HIEFFPLA_NET_0_118719);
    
    \U_ELK15_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2\ : IOPADN_BI
      port map(DB => \U_ELK15_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, 
        E => \U_ELK15_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET3\, PAD
         => ELK15_DAT_N, N2POUT => 
        \U_ELK15_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2_N2P\);
    
    \U50_PATTERNS/ELINK_ADDRA_17[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120027, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_11, Q => 
        \U50_PATTERNS/ELINK_ADDRA_17[4]\);
    
    HIEFFPLA_INST_0_54905 : AO1A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_0[6]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_0[8]_net_1\, C => 
        HIEFFPLA_NET_0_117173, Y => HIEFFPLA_NET_0_117174);
    
    \U_ELK16_CH/U_ELK1_CMD_TX/SER_OUT_FI\ : DFN1C0
      port map(D => 
        \U_ELK16_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_10, Q
         => \U_ELK16_CH/U_ELK1_CMD_TX/SER_OUT_FI_net_1\);
    
    \U_ELK3_CH/U_SLAVE_1ELK/Q[9]\ : DFN1C0
      port map(D => \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/Q[9]_net_1\);
    
    \U_ELK8_CH/U_SLAVE_1ELK/Q[2]\ : DFN1C0
      port map(D => \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/Q[2]_net_1\);
    
    HIEFFPLA_INST_0_47852 : MX2
      port map(A => 
        \U_ELK15_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]_net_1\, B => 
        \U_ELK15_CH/ELK_TX_DAT[3]\, S => 
        \U_ELK15_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118422);
    
    HIEFFPLA_INST_0_40648 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_14[6]\, B => 
        HIEFFPLA_NET_0_119566, S => HIEFFPLA_NET_0_119249, Y => 
        HIEFFPLA_NET_0_119825);
    
    HIEFFPLA_INST_0_43683 : NAND3C
      port map(A => \U50_PATTERNS/SM_BANK_SEL[1]\, B => 
        \U50_PATTERNS/SM_BANK_SEL[19]\, C => 
        \U50_PATTERNS/SM_BANK_SEL[2]\, Y => HIEFFPLA_NET_0_119242);
    
    \U_ELK12_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]\ : DFN1C0
      port map(D => \U_ELK12_CH/U_SLAVE_1ELK/Q[14]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]_net_1\);
    
    HIEFFPLA_INST_0_52438 : MX2
      port map(A => HIEFFPLA_NET_0_117515, B => 
        HIEFFPLA_NET_0_117511, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[3]\, Y => 
        HIEFFPLA_NET_0_117563);
    
    HIEFFPLA_INST_0_51507 : XOR2
      port map(A => \U_EXEC_MASTER/PRESCALE[1]\, B => 
        \U_EXEC_MASTER/PRESCALE[0]\, Y => HIEFFPLA_NET_0_117760);
    
    HIEFFPLA_INST_0_61115 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_3[0]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_19[0]\, S
         => \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_1[4]_net_1\, 
        Y => HIEFFPLA_NET_0_116171);
    
    HIEFFPLA_INST_0_54958 : AND2A
      port map(A => HIEFFPLA_NET_0_117218, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_3[6]_net_1\, Y => 
        HIEFFPLA_NET_0_117156);
    
    HIEFFPLA_INST_0_52386 : MX2
      port map(A => HIEFFPLA_NET_0_117526, B => 
        HIEFFPLA_NET_0_117482, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[1]\, Y => 
        HIEFFPLA_NET_0_117570);
    
    HIEFFPLA_INST_0_42914 : NAND3
      port map(A => \U50_PATTERNS/REG_STATE[4]_net_1\, B => 
        \U50_PATTERNS/REG_STATE[2]_net_1\, C => 
        \U50_PATTERNS/REG_STATE[3]_net_1\, Y => 
        HIEFFPLA_NET_0_119426);
    
    HIEFFPLA_INST_0_56389 : NAND3C
      port map(A => HIEFFPLA_NET_0_116832, B => 
        HIEFFPLA_NET_0_116848, C => HIEFFPLA_NET_0_116856, Y => 
        HIEFFPLA_NET_0_116880);
    
    HIEFFPLA_INST_0_112355 : AO1D
      port map(A => HIEFFPLA_NET_0_116740, B => 
        HIEFFPLA_NET_0_116708, C => HIEFFPLA_NET_0_116678, Y => 
        HIEFFPLA_NET_0_115815);
    
    HIEFFPLA_INST_0_45118 : MX2
      port map(A => HIEFFPLA_NET_0_118971, B => 
        \U50_PATTERNS/WR_USB_ADBUS[4]\, S => 
        HIEFFPLA_NET_0_119486, Y => HIEFFPLA_NET_0_118981);
    
    HIEFFPLA_INST_0_49588 : MX2
      port map(A => 
        \U_ELK3_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]_net_1\, B => 
        \U_ELK3_CH/ELK_TX_DAT[6]\, S => 
        \U_ELK3_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118109);
    
    HIEFFPLA_INST_0_39317 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_1[3]\, B => 
        HIEFFPLA_NET_0_119520, S => HIEFFPLA_NET_0_119243, Y => 
        HIEFFPLA_NET_0_120004);
    
    \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[14]\ : DFN1C0
      port map(D => 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[14]_net_1\);
    
    HIEFFPLA_INST_0_61196 : MX2
      port map(A => HIEFFPLA_NET_0_117190, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_20[0]\, S => 
        HIEFFPLA_NET_0_117141, Y => HIEFFPLA_NET_0_116160);
    
    \U_ELK15_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]\ : DFN1C0
      port map(D => \U_ELK15_CH/U_SLAVE_1ELK/Q[14]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]_net_1\);
    
    HIEFFPLA_INST_0_55157 : NAND3
      port map(A => HIEFFPLA_NET_0_117414, B => 
        HIEFFPLA_NET_0_117359, C => HIEFFPLA_NET_0_117085, Y => 
        HIEFFPLA_NET_0_117109);
    
    \U_ELK6_CH/U_SLAVE_1ELK/RECD_SER_WORD[6]\ : DFN1C0
      port map(D => \U_ELK6_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[6]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_6[6]\);
    
    HIEFFPLA_INST_0_50113 : AND2A
      port map(A => \OP_MODE_c_4[1]\, B => \PATT_ELK_DAT_5[4]\, Y
         => HIEFFPLA_NET_0_118009);
    
    HIEFFPLA_INST_0_42426 : AND2
      port map(A => HIEFFPLA_NET_0_119473, B => 
        \U50_PATTERNS/RD_XFER_TYPE[3]_net_1\, Y => 
        HIEFFPLA_NET_0_119538);
    
    HIEFFPLA_INST_0_38266 : MX2
      port map(A => \U50_PATTERNS/ELINKS_STOP_ADDR[3]\, B => 
        \U50_PATTERNS/ELINKS_STOP_ADDR_T[3]\, S => 
        HIEFFPLA_NET_0_119472, Y => HIEFFPLA_NET_0_120124);
    
    \U_ELK10_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]\ : DFN1C0
      port map(D => \U_ELK10_CH/U_SLAVE_1ELK/Q[5]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]_net_1\);
    
    \U_ELK3_CH/U_SLAVE_1ELK/Q[0]\ : DFN1C0
      port map(D => \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/Q[0]_net_1\);
    
    HIEFFPLA_INST_0_61415 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_22[1]\, B => 
        HIEFFPLA_NET_0_117167, S => HIEFFPLA_NET_0_117080, Y => 
        HIEFFPLA_NET_0_116129);
    
    HIEFFPLA_INST_0_51827 : AND2
      port map(A => \U_MASTER_DES/U13A_ADJ_160M/BITCNT[0]\, B => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[1]\, Y => 
        HIEFFPLA_NET_0_117684);
    
    \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[0]\ : DFN1C0
      port map(D => 
        \U_ELK3_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\);
    
    HIEFFPLA_INST_0_44784 : XOR2
      port map(A => \OP_MODE[0]\, B => 
        \U50_PATTERNS/U4E_REGCROSS/SAMP_TWO[0]_net_1\, Y => 
        HIEFFPLA_NET_0_119050);
    
    HIEFFPLA_INST_0_60107 : MX2
      port map(A => HIEFFPLA_NET_0_116677, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_6[1]\, S => 
        HIEFFPLA_NET_0_117211, Y => HIEFFPLA_NET_0_116309);
    
    HIEFFPLA_INST_0_52019 : AND2B
      port map(A => HIEFFPLA_NET_0_117639, B => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[1]\, Y => 
        HIEFFPLA_NET_0_117651);
    
    HIEFFPLA_INST_0_47331 : AND2
      port map(A => \U_ELK13_CH/ELK_TX_DAT[0]\, B => 
        \U_ELK13_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118517);
    
    HIEFFPLA_INST_0_43218 : AND3A
      port map(A => \U50_PATTERNS/REG_STATE_0[4]_net_1\, B => 
        \U50_PATTERNS/REG_STATE[3]_net_1\, C => 
        \U50_PATTERNS/REG_STATE_0[2]_net_1\, Y => 
        HIEFFPLA_NET_0_119345);
    
    \U_ELK14_CH/U_SLAVE_1ELK/RECD_SER_WORD[4]\ : DFN1C0
      port map(D => \U_ELK14_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[4]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_14[4]\);
    
    \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[14]\ : DFN1C0
      port map(D => \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\, 
        CLK => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[14]_net_1\);
    
    HIEFFPLA_INST_0_44694 : MX2
      port map(A => \OP_MODE_c[5]\, B => 
        \U50_PATTERNS/U4E_REGCROSS/SAMP_TWO[5]_net_1\, S => 
        HIEFFPLA_NET_0_119072, Y => HIEFFPLA_NET_0_119065);
    
    \U_MASTER_DES/U13C_MASTER_DESER/TUNE_CLKPHASE[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_115947, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_12, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/TUNE_CLKPHASE[2]\);
    
    \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[8]\ : DFN1C0
      port map(D => \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\);
    
    \U50_PATTERNS/ELINK_DINA_9[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119714, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_20, Q => 
        \U50_PATTERNS/ELINK_DINA_9[5]\);
    
    HIEFFPLA_INST_0_62887 : MX2
      port map(A => HIEFFPLA_NET_0_115897, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[11]\, S => 
        HIEFFPLA_NET_0_117073, Y => HIEFFPLA_NET_0_115932);
    
    HIEFFPLA_INST_0_43112 : AOI1C
      port map(A => HIEFFPLA_NET_0_118694, B => 
        \U50_PATTERNS/REG_STATE[3]_net_1\, C => 
        HIEFFPLA_NET_0_118996, Y => HIEFFPLA_NET_0_119373);
    
    HIEFFPLA_INST_0_47868 : AND2A
      port map(A => \OP_MODE_c_6[1]\, B => \PATT_ELK_DAT_15[0]\, 
        Y => HIEFFPLA_NET_0_118418);
    
    HIEFFPLA_INST_0_37819 : AND2
      port map(A => \U200B_ELINKS/N_232_li\, B => 
        \U200B_ELINKS/GP_PG_SM[9]_net_1\, Y => 
        HIEFFPLA_NET_0_120199);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_1[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116474, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_17, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_1[1]\);
    
    AFLSDF_INV_6 : INV
      port map(A => P_USB_MASTER_EN_c_22, Y => \AFLSDF_INV_6\);
    
    \U_ELK14_CH/U_ELK1_SERDAT_SOURCE/SERDAT[4]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118459, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_6, Q => 
        \U_ELK14_CH/ELK_TX_DAT[4]\);
    
    HIEFFPLA_INST_0_44568 : MX2
      port map(A => \ELKS_STOP_ADDR[2]\, B => 
        \U50_PATTERNS/U4D_REGCROSS/SAMP_TWO[2]_net_1\, S => 
        HIEFFPLA_NET_0_119093, Y => HIEFFPLA_NET_0_119089);
    
    \U_ELK15_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118423, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_6, Q => 
        \U_ELK15_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]_net_1\);
    
    HIEFFPLA_INST_0_46155 : AO1
      port map(A => HIEFFPLA_NET_0_119263, B => 
        \U50_PATTERNS/ELINK_DOUTA_8[0]\, C => 
        HIEFFPLA_NET_0_118929, Y => HIEFFPLA_NET_0_118754);
    
    HIEFFPLA_INST_0_50105 : MX2
      port map(A => 
        \U_ELK5_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]_net_1\, B => 
        \U_ELK5_CH/ELK_TX_DAT[7]\, S => 
        \U_ELK5_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118015);
    
    \U_ELK5_CH/U_SLAVE_1ELK/RECD_SER_WORD[3]\ : DFN1C0
      port map(D => \U_ELK5_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[3]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_5[3]\);
    
    \U_ELK12_CH/U_ELK1_SERDAT_SOURCE/SERDAT[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118552, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_2, Q => 
        \U_ELK12_CH/ELK_TX_DAT[1]\);
    
    HIEFFPLA_INST_0_50479 : MX2
      port map(A => HIEFFPLA_NET_0_117936, B => 
        HIEFFPLA_NET_0_117945, S => \BIT_OS_SEL[0]\, Y => 
        \U_ELK6_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[0]\);
    
    HIEFFPLA_INST_0_39434 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_3[0]\, B => 
        HIEFFPLA_NET_0_119524, S => HIEFFPLA_NET_0_119247, Y => 
        HIEFFPLA_NET_0_119991);
    
    \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[12]\ : DFN1C0
      port map(D => \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\, 
        CLK => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\);
    
    HIEFFPLA_INST_0_60259 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_8[3]\, B => 
        HIEFFPLA_NET_0_116815, S => HIEFFPLA_NET_0_117160, Y => 
        HIEFFPLA_NET_0_116290);
    
    HIEFFPLA_INST_0_57452 : AND3B
      port map(A => HIEFFPLA_NET_0_116740, B => 
        HIEFFPLA_NET_0_116686, C => HIEFFPLA_NET_0_116620, Y => 
        HIEFFPLA_NET_0_116679);
    
    HIEFFPLA_INST_0_50413 : MX2
      port map(A => \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[3]_net_1\, B
         => \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\, S => 
        \BIT_OS_SEL_5[2]\, Y => HIEFFPLA_NET_0_117954);
    
    \U_ELK15_CH/U_SLAVE_1ELK/Q[4]\ : DFN1C0
      port map(D => \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/Q[4]_net_1\);
    
    \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[4]\ : DFN1C0
      port map(D => 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\);
    
    \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[14]\ : DFN1C0
      port map(D => 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]_net_1\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[14]_net_1\);
    
    HIEFFPLA_INST_0_62959 : MX2
      port map(A => HIEFFPLA_NET_0_115888, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[6]\, S => 
        HIEFFPLA_NET_0_117073, Y => HIEFFPLA_NET_0_115924);
    
    HIEFFPLA_INST_0_55520 : MX2
      port map(A => HIEFFPLA_NET_0_116986, B => 
        HIEFFPLA_NET_0_117033, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[2]\, Y => 
        HIEFFPLA_NET_0_117026);
    
    HIEFFPLA_INST_0_52502 : MX2
      port map(A => HIEFFPLA_NET_0_117499, B => 
        HIEFFPLA_NET_0_117495, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_1[3]\, Y => 
        HIEFFPLA_NET_0_117555);
    
    HIEFFPLA_INST_0_60834 : MX2
      port map(A => HIEFFPLA_NET_0_117181, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_16[2]\, S => 
        HIEFFPLA_NET_0_117142, Y => HIEFFPLA_NET_0_116213);
    
    HIEFFPLA_INST_0_49628 : MX2
      port map(A => \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[2]_net_1\, B
         => \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\, S => 
        \BIT_OS_SEL_7[2]\, Y => HIEFFPLA_NET_0_118094);
    
    \U_ELK5_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]\ : DFN1C0
      port map(D => \U_ELK5_CH/U_SLAVE_1ELK/Q[7]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]_net_1\);
    
    \U_ELK19_CH/U_ELK1_SERDAT_SOURCE/SERDAT[4]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118234, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_15, Q => 
        \U_ELK19_CH/ELK_TX_DAT[4]\);
    
    HIEFFPLA_INST_0_56771 : NAND3
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_0[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_0[2]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_0[3]\, Y => 
        HIEFFPLA_NET_0_116802);
    
    \U_ELK9_CH/U_ELK1_SERDAT_SOURCE/SERDAT[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117832, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_7, Q => 
        \U_ELK9_CH/ELK_TX_DAT[1]\);
    
    HIEFFPLA_INST_0_62649 : MX2
      port map(A => HIEFFPLA_NET_0_117131, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_9[2]\, S => 
        HIEFFPLA_NET_0_117183, Y => HIEFFPLA_NET_0_115963);
    
    \U_ELK19_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]\ : DFN1C0
      port map(D => \U_ELK19_CH/U_SLAVE_1ELK/Q[13]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]_net_1\);
    
    HIEFFPLA_INST_0_53387 : MX2
      port map(A => HIEFFPLA_NET_0_117292, B => 
        HIEFFPLA_NET_0_117314, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[2]_net_1\, Y
         => HIEFFPLA_NET_0_117417);
    
    HIEFFPLA_INST_0_51595 : AX1C
      port map(A => HIEFFPLA_NET_0_117748, B => 
        HIEFFPLA_NET_0_117753, C => HIEFFPLA_NET_0_117732, Y => 
        HIEFFPLA_NET_0_117737);
    
    HIEFFPLA_INST_0_50316 : MX2
      port map(A => \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\, 
        B => \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[14]_net_1\, S => 
        \BIT_OS_SEL_7[2]\, Y => HIEFFPLA_NET_0_117978);
    
    HIEFFPLA_INST_0_61562 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_7[0]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_23[0]\, S
         => \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[4]_net_1\, 
        Y => HIEFFPLA_NET_0_116109);
    
    HIEFFPLA_INST_0_40057 : MX2
      port map(A => HIEFFPLA_NET_0_119884, B => 
        \U50_PATTERNS/ELINK_BLKA[7]\, S => 
        \U50_PATTERNS/SM_BANK_SEL[20]\, Y => 
        HIEFFPLA_NET_0_119918);
    
    \U_ELK3_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118109, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_16, Q => 
        \U_ELK3_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]_net_1\);
    
    \U200B_ELINKS/RX_SER_WORD_1DEL[2]\ : DFN1C0
      port map(D => \ELK_RX_SER_WORD_0[2]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c_23, Q => 
        \U200B_ELINKS/RX_SER_WORD_1DEL[2]_net_1\);
    
    \U_ELK13_CH/U_SLAVE_1ELK/Q[10]\ : DFN1C0
      port map(D => \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/Q[10]_net_1\);
    
    HIEFFPLA_INST_0_48993 : MX2
      port map(A => HIEFFPLA_NET_0_118230, B => 
        HIEFFPLA_NET_0_118228, S => \BIT_OS_SEL_2[0]\, Y => 
        \U_ELK19_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[1]\);
    
    HIEFFPLA_INST_0_48120 : NAND2B
      port map(A => \OP_MODE_c_2[1]\, B => \PATT_ELK_DAT_16[3]\, 
        Y => HIEFFPLA_NET_0_118370);
    
    \U_ELK15_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118426, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_9, Q => 
        \U_ELK15_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]_net_1\);
    
    HIEFFPLA_INST_0_46588 : MX2
      port map(A => 
        \U_ELK10_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]_net_1\, B => 
        \U_ELK10_CH/ELK_TX_DAT[2]\, S => 
        \U_ELK10_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118651);
    
    \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[10]\ : DFN1C0
      port map(D => \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\);
    
    \U50_PATTERNS/TFC_RWA/U1\ : DFN1P0
      port map(D => HIEFFPLA_NET_0_119189, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_3, Q => \U50_PATTERNS/TFC_RWA\);
    
    HIEFFPLA_INST_0_49118 : AND2A
      port map(A => \OP_MODE_c_5[1]\, B => \PATT_ELK_DAT_1[5]\, Y
         => HIEFFPLA_NET_0_118188);
    
    HIEFFPLA_INST_0_51116 : MX2
      port map(A => \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\, B
         => \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[13]_net_1\, S => 
        \BIT_OS_SEL_3[2]\, Y => HIEFFPLA_NET_0_117825);
    
    HIEFFPLA_INST_0_44846 : MX2
      port map(A => USB_RD_BI, B => HIEFFPLA_NET_0_119035, S => 
        HIEFFPLA_NET_0_119033, Y => HIEFFPLA_NET_0_119036);
    
    \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[2]\ : DFN1C0
      port map(D => \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\);
    
    \U_EXEC_MASTER/DEV_RST_0B\ : DFN1C0
      port map(D => \VCC\, CLK => CCC_160M_FXD, CLR => 
        DEV_RST_B_c, Q => \U_EXEC_MASTER/DEV_RST_0B_net_1\);
    
    \U50_PATTERNS/ELINK_ADDRA_5[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119971, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_3, Q => 
        \U50_PATTERNS/ELINK_ADDRA_5[4]\);
    
    HIEFFPLA_INST_0_62460 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_5[2]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_6[2]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_2[0]\, Y => 
        HIEFFPLA_NET_0_115986);
    
    HIEFFPLA_INST_0_49266 : MX2
      port map(A => HIEFFPLA_NET_0_118177, B => 
        HIEFFPLA_NET_0_118176, S => \BIT_OS_SEL_2[0]\, Y => 
        \U_ELK1_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[4]\);
    
    HIEFFPLA_INST_0_55363 : AND3B
      port map(A => HIEFFPLA_NET_0_117046, B => 
        HIEFFPLA_NET_0_117049, C => HIEFFPLA_NET_0_115909, Y => 
        HIEFFPLA_NET_0_117050);
    
    HIEFFPLA_INST_0_38346 : MX2
      port map(A => \U50_PATTERNS/ELINKS_STOP_ADDR_T[5]\, B => 
        \U50_PATTERNS/RD_USB_ADBUS[5]\, S => 
        HIEFFPLA_NET_0_119413, Y => HIEFFPLA_NET_0_120114);
    
    \U_ELK11_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]\ : DFN1C0
      port map(D => \U_ELK11_CH/U_SLAVE_1ELK/Q[2]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_13[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116539, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_12, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_13[3]\);
    
    \U_EXEC_MASTER/MPOR_B_16\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117787, CLK => CLK_40M_GL, CLR
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_1\, Q => 
        P_MASTER_POR_B_c_16);
    
    \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[5]\ : DFN1C0
      port map(D => \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\);
    
    HIEFFPLA_INST_0_42503 : MX2
      port map(A => \U50_PATTERNS/REG_ADDR[7]\, B => 
        HIEFFPLA_NET_0_119502, S => HIEFFPLA_NET_0_119007, Y => 
        HIEFFPLA_NET_0_119526);
    
    HIEFFPLA_INST_0_37163 : AND3B
      port map(A => HIEFFPLA_NET_0_120259, B => 
        \U200A_TFC/GP_PG_SM[10]_net_1\, C => 
        HIEFFPLA_NET_0_120325, Y => HIEFFPLA_NET_0_120336);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_26[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116080, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_12, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_26[0]\);
    
    \U_ELK15_CH/U_ELK1_SERDAT_SOURCE/SERDAT[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118417, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_8, Q => 
        \U_ELK15_CH/ELK_TX_DAT[1]\);
    
    HIEFFPLA_INST_0_54317 : MX2
      port map(A => HIEFFPLA_NET_0_116206, B => 
        HIEFFPLA_NET_0_116096, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_2[3]_net_1\, Y
         => HIEFFPLA_NET_0_117281);
    
    \U50_PATTERNS/ELINK_ADDRA_18[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120021, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_12, Q => 
        \U50_PATTERNS/ELINK_ADDRA_18[2]\);
    
    \U_ELK17_CH/U_SLAVE_1ELK/RECD_SER_WORD[2]\ : DFN1C0
      port map(D => \U_ELK17_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[2]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_17[2]\);
    
    HIEFFPLA_INST_0_56418 : AND3
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[4]_net_1\, B => 
        HIEFFPLA_NET_0_117427, C => HIEFFPLA_NET_0_117423, Y => 
        HIEFFPLA_NET_0_116871);
    
    HIEFFPLA_INST_0_38050 : AND3B
      port map(A => \U200B_ELINKS/LOC_STRT_ADDR[6]\, B => 
        HIEFFPLA_NET_0_120190, C => HIEFFPLA_NET_0_120234, Y => 
        HIEFFPLA_NET_0_120165);
    
    \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[10]\ : DFN1C0
      port map(D => \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\);
    
    \U50_PATTERNS/ELINKS_STRT_ADDR_T[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120101, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_21, Q => 
        \U50_PATTERNS/ELINKS_STRT_ADDR_T[2]\);
    
    HIEFFPLA_INST_0_62896 : MX2
      port map(A => HIEFFPLA_NET_0_115895, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[12]\, S => 
        HIEFFPLA_NET_0_117073, Y => HIEFFPLA_NET_0_115931);
    
    HIEFFPLA_INST_0_51705 : NAND2B
      port map(A => 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM[4]_net_1\, B => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[0]_net_1\, Y => 
        HIEFFPLA_NET_0_117721);
    
    HIEFFPLA_INST_0_45673 : AO1A
      port map(A => HIEFFPLA_NET_0_119475, B => 
        \U50_PATTERNS/ELINKS_STOP_ADDR[4]\, C => 
        HIEFFPLA_NET_0_118771, Y => HIEFFPLA_NET_0_118867);
    
    HIEFFPLA_INST_0_62562 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_7[1]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_8[1]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[0]\, Y => 
        HIEFFPLA_NET_0_115974);
    
    HIEFFPLA_INST_0_50459 : MX2
      port map(A => \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\, B
         => \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[12]_net_1\, S => 
        \BIT_OS_SEL_5[2]\, Y => HIEFFPLA_NET_0_117947);
    
    \U_ELK8_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]\ : DFN1C0
      port map(D => \U_ELK8_CH/U_SLAVE_1ELK/Q[7]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]_net_1\);
    
    HIEFFPLA_INST_0_161265 : DFN1C0
      port map(D => \U_ELK9_CH/ELK_TX_DAT[5]\, CLK => 
        CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_0, Q => 
        HIEFFPLA_NET_0_161290);
    
    HIEFFPLA_INST_0_37982 : MX2
      port map(A => \U200B_ELINKS/LOC_STRT_ADDR[0]\, B => 
        \ELKS_STRT_ADDR[0]\, S => 
        \U200B_ELINKS/GP_PG_SM_0[10]_net_1\, Y => 
        HIEFFPLA_NET_0_120179);
    
    HIEFFPLA_INST_0_38741 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_12[3]\, B => 
        HIEFFPLA_NET_0_119520, S => HIEFFPLA_NET_0_119295, Y => 
        HIEFFPLA_NET_0_120068);
    
    HIEFFPLA_INST_0_63004 : NOR3B
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[7]\, 
        B => HIEFFPLA_NET_0_115904, C => HIEFFPLA_NET_0_115907, Y
         => HIEFFPLA_NET_0_115917);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_16[4]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116211, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_5, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_16[4]\);
    
    \U50_PATTERNS/U110_PATT_ELINK_BLK/DPRT_512X9_SRAM_R0C0\ : 
        RAM4K9
      generic map(MEMORYFILE => "DPRT_512X9_SRAM_R0C0.mem")

      port map(ADDRA11 => AFLSDF_GND, ADDRA10 => AFLSDF_GND, 
        ADDRA9 => AFLSDF_GND, ADDRA8 => \GND\, ADDRA7 => 
        \U50_PATTERNS/ELINK_ADDRA_10[7]\, ADDRA6 => 
        \U50_PATTERNS/ELINK_ADDRA_10[6]\, ADDRA5 => 
        \U50_PATTERNS/ELINK_ADDRA_10[5]\, ADDRA4 => 
        \U50_PATTERNS/ELINK_ADDRA_10[4]\, ADDRA3 => 
        \U50_PATTERNS/ELINK_ADDRA_10[3]\, ADDRA2 => 
        \U50_PATTERNS/ELINK_ADDRA_10[2]\, ADDRA1 => 
        \U50_PATTERNS/ELINK_ADDRA_10[1]\, ADDRA0 => 
        \U50_PATTERNS/ELINK_ADDRA_10[0]\, ADDRB11 => AFLSDF_GND, 
        ADDRB10 => AFLSDF_GND, ADDRB9 => AFLSDF_GND, ADDRB8 => 
        \GND\, ADDRB7 => \ELKS_ADDRB[7]\, ADDRB6 => 
        \ELKS_ADDRB_0[6]\, ADDRB5 => \ELKS_ADDRB[5]\, ADDRB4 => 
        \ELKS_ADDRB_0[4]\, ADDRB3 => \ELKS_ADDRB[3]\, ADDRB2 => 
        \ELKS_ADDRB_0[2]\, ADDRB1 => \ELKS_ADDRB[1]\, ADDRB0 => 
        \ELKS_ADDRB[0]\, DINA8 => \GND\, DINA7 => 
        \U50_PATTERNS/ELINK_DINA_10[7]\, DINA6 => 
        \U50_PATTERNS/ELINK_DINA_10[6]\, DINA5 => 
        \U50_PATTERNS/ELINK_DINA_10[5]\, DINA4 => 
        \U50_PATTERNS/ELINK_DINA_10[4]\, DINA3 => 
        \U50_PATTERNS/ELINK_DINA_10[3]\, DINA2 => 
        \U50_PATTERNS/ELINK_DINA_10[2]\, DINA1 => 
        \U50_PATTERNS/ELINK_DINA_10[1]\, DINA0 => 
        \U50_PATTERNS/ELINK_DINA_10[0]\, DINB8 => \GND\, DINB7
         => \ELK_RX_SER_WORD_10[7]\, DINB6 => 
        \ELK_RX_SER_WORD_10[6]\, DINB5 => \ELK_RX_SER_WORD_10[5]\, 
        DINB4 => \ELK_RX_SER_WORD_10[4]\, DINB3 => 
        \ELK_RX_SER_WORD_10[3]\, DINB2 => \ELK_RX_SER_WORD_10[2]\, 
        DINB1 => \ELK_RX_SER_WORD_10[1]\, DINB0 => 
        \ELK_RX_SER_WORD_10[0]\, WIDTHA0 => \VCC\, WIDTHA1 => 
        \VCC\, WIDTHB0 => \VCC\, WIDTHB1 => \VCC\, PIPEA => \VCC\, 
        PIPEB => \VCC\, WMODEA => \GND\, WMODEB => \GND\, BLKA
         => \U50_PATTERNS/ELINK_BLKA[10]\, BLKB => 
        ELKS_RAM_BLKB_EN, WENA => \U50_PATTERNS/ELINK_RWA[10]\, 
        WENB => ELKS_RWB, CLKA => CLK60MHZ, CLKB => CLK_40M_GL, 
        RESET => P_USB_MASTER_EN_c_0, DOUTA8 => OPEN, DOUTA7 => 
        \U50_PATTERNS/ELINK_DOUTA_10[7]\, DOUTA6 => 
        \U50_PATTERNS/ELINK_DOUTA_10[6]\, DOUTA5 => 
        \U50_PATTERNS/ELINK_DOUTA_10[5]\, DOUTA4 => 
        \U50_PATTERNS/ELINK_DOUTA_10[4]\, DOUTA3 => 
        \U50_PATTERNS/ELINK_DOUTA_10[3]\, DOUTA2 => 
        \U50_PATTERNS/ELINK_DOUTA_10[2]\, DOUTA1 => 
        \U50_PATTERNS/ELINK_DOUTA_10[1]\, DOUTA0 => 
        \U50_PATTERNS/ELINK_DOUTA_10[0]\, DOUTB8 => OPEN, DOUTB7
         => \PATT_ELK_DAT_10[7]\, DOUTB6 => \PATT_ELK_DAT_10[6]\, 
        DOUTB5 => \PATT_ELK_DAT_10[5]\, DOUTB4 => 
        \PATT_ELK_DAT_10[4]\, DOUTB3 => \PATT_ELK_DAT_10[3]\, 
        DOUTB2 => \PATT_ELK_DAT_10[2]\, DOUTB1 => 
        \PATT_ELK_DAT_10[1]\, DOUTB0 => \PATT_ELK_DAT_10[0]\);
    
    \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[13]\ : DFN1C0
      port map(D => 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[13]_net_1\);
    
    \U_ELK11_CH/U_SLAVE_1ELK/RECD_SER_WORD[7]\ : DFN1C0
      port map(D => \U_ELK11_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[7]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_11[7]\);
    
    \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[10]\ : DFN1C0
      port map(D => \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\);
    
    HIEFFPLA_INST_0_51720 : NAND2B
      port map(A => 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM_0[4]_net_1\, B => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[73]_net_1\, Y => 
        HIEFFPLA_NET_0_117706);
    
    HIEFFPLA_INST_0_56330 : AO1
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[5]_net_1\, B => 
        HIEFFPLA_NET_0_117429, C => HIEFFPLA_NET_0_116868, Y => 
        HIEFFPLA_NET_0_116892);
    
    HIEFFPLA_INST_0_42125 : MX2
      port map(A => \U50_PATTERNS/OP_MODE[4]\, B => 
        \U50_PATTERNS/OP_MODE_T[4]\, S => HIEFFPLA_NET_0_119472, 
        Y => HIEFFPLA_NET_0_119613);
    
    \U50_PATTERNS/WR_XFER_TYPE[5]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118684, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c, Q => 
        \U50_PATTERNS/WR_XFER_TYPE[5]_net_1\);
    
    \U_ELK9_CH/U_ELK1_SERDAT_SOURCE/SERDAT[4]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117829, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_7, Q => 
        \U_ELK9_CH/ELK_TX_DAT[4]\);
    
    \U_ELK10_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118645, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_3, Q => 
        \U_ELK10_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]_net_1\);
    
    \U_ELK11_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL\ : DFN1C0
      port map(D => \U_ELK11_CH/ELK_IN_R_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL_net_1\);
    
    HIEFFPLA_INST_0_52582 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_9[0]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_10[0]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[0]\, Y => 
        HIEFFPLA_NET_0_117544);
    
    \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[2]\ : DFN1C0
      port map(D => \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\);
    
    \U_ELK14_CH/U_SLAVE_1ELK/RECD_SER_WORD[2]\ : DFN1C0
      port map(D => \U_ELK14_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[2]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_14[2]\);
    
    \U_ELK19_CH/U_SLAVE_1ELK/RECD_SER_WORD[0]\ : DFN1C0
      port map(D => \U_ELK19_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[0]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_19[0]\);
    
    \U50_PATTERNS/ELINK_BLKA[5]/U1\ : DFN1P0
      port map(D => HIEFFPLA_NET_0_119920, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_19, Q => 
        \U50_PATTERNS/ELINK_BLKA[5]\);
    
    HIEFFPLA_INST_0_52188 : MX2
      port map(A => \U_MASTER_DES/AUX_SUPDATE\, B => 
        HIEFFPLA_NET_0_117613, S => HIEFFPLA_NET_0_117628, Y => 
        HIEFFPLA_NET_0_117614);
    
    HIEFFPLA_INST_0_44875 : AND3C
      port map(A => \U50_PATTERNS/REG_STATE[3]_net_1\, B => 
        \U50_PATTERNS/USB_RXF_B\, C => 
        \U50_PATTERNS/REG_STATE[4]_net_1\, Y => 
        HIEFFPLA_NET_0_119030);
    
    \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[3]\ : DFN1C0
      port map(D => 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[3]_net_1\);
    
    HIEFFPLA_INST_0_47132 : MX2
      port map(A => HIEFFPLA_NET_0_118543, B => 
        HIEFFPLA_NET_0_118539, S => \BIT_OS_SEL_4[1]\, Y => 
        HIEFFPLA_NET_0_118545);
    
    HIEFFPLA_INST_0_41833 : AOI1B
      port map(A => HIEFFPLA_NET_0_119389, B => 
        \U50_PATTERNS/SM_BANK_SEL[6]\, C => HIEFFPLA_NET_0_119658, 
        Y => HIEFFPLA_NET_0_119687);
    
    \U_ELK5_CH/U_SLAVE_1ELK/Q[12]\ : DFN1C0
      port map(D => \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/Q[12]_net_1\);
    
    HIEFFPLA_INST_0_44840 : NAND3B
      port map(A => \U50_PATTERNS/REG_STATE[3]_net_1\, B => 
        HIEFFPLA_NET_0_119450, C => 
        \U50_PATTERNS/REG_STATE[2]_net_1\, Y => 
        HIEFFPLA_NET_0_119037);
    
    \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[11]\ : DFN1C0
      port map(D => \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\);
    
    HIEFFPLA_INST_0_41868 : AOI1B
      port map(A => HIEFFPLA_NET_0_119389, B => 
        \U50_PATTERNS/SM_BANK_SEL[18]\, C => 
        HIEFFPLA_NET_0_119649, Y => HIEFFPLA_NET_0_119679);
    
    \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[14]\ : DFN1C0
      port map(D => \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\, 
        CLK => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[14]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/RECD_SER_WORD[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_116901, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_29, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/RECD_SER_WORD[3]_net_1\);
    
    HIEFFPLA_INST_0_60079 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_6[1]\, B => 
        HIEFFPLA_NET_0_116309, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_0[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116313);
    
    HIEFFPLA_INST_0_39587 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_5[1]\, B => 
        HIEFFPLA_NET_0_119523, S => HIEFFPLA_NET_0_119251, Y => 
        HIEFFPLA_NET_0_119974);
    
    HIEFFPLA_INST_0_61301 : MX2
      port map(A => HIEFFPLA_NET_0_117190, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_21[0]\, S => 
        HIEFFPLA_NET_0_117144, Y => HIEFFPLA_NET_0_116145);
    
    HIEFFPLA_INST_0_44344 : MX2
      port map(A => \TFC_STOP_ADDR[0]\, B => 
        \U50_PATTERNS/U4B_REGCROSS/SAMP_TWO[0]_net_1\, S => 
        HIEFFPLA_NET_0_119135, Y => HIEFFPLA_NET_0_119133);
    
    \U_ELK18_CH/U_SLAVE_1ELK/RECD_SER_WORD[1]\ : DFN1C0
      port map(D => \U_ELK18_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[1]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_18[1]\);
    
    HIEFFPLA_INST_0_61724 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_25[2]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_26[2]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_4[0]\, Y => 
        HIEFFPLA_NET_0_116087);
    
    HIEFFPLA_INST_0_52776 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_3[3]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_4[3]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[0]\, Y => 
        HIEFFPLA_NET_0_117513);
    
    HIEFFPLA_INST_0_44421 : XO1
      port map(A => \U50_PATTERNS/U4B_REGCROSS/SAMP_TWO[2]_net_1\, 
        B => \TFC_STOP_ADDR[2]\, C => HIEFFPLA_NET_0_119119, Y
         => HIEFFPLA_NET_0_119123);
    
    HIEFFPLA_INST_0_60477 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_11[4]\, B => 
        HIEFFPLA_NET_0_117100, S => HIEFFPLA_NET_0_117348, Y => 
        HIEFFPLA_NET_0_116261);
    
    HIEFFPLA_INST_0_40133 : AOI1C
      port map(A => \U50_PATTERNS/ELINK_BLKA[1]\, B => 
        HIEFFPLA_NET_0_119648, C => HIEFFPLA_NET_0_119895, Y => 
        HIEFFPLA_NET_0_119896);
    
    HIEFFPLA_INST_0_56423 : AND3
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[5]_net_1\, B => 
        HIEFFPLA_NET_0_117427, C => HIEFFPLA_NET_0_117423, Y => 
        HIEFFPLA_NET_0_116870);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_30[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116353, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_18, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_30[3]\);
    
    \U50_PATTERNS/ELINK_ADDRA_4[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119983, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_2, Q => 
        \U50_PATTERNS/ELINK_ADDRA_4[0]\);
    
    HIEFFPLA_INST_0_45063 : AO1
      port map(A => \U50_PATTERNS/REG_STATE[4]_net_1\, B => 
        HIEFFPLA_NET_0_119368, C => HIEFFPLA_NET_0_118988, Y => 
        HIEFFPLA_NET_0_118989);
    
    HIEFFPLA_INST_0_41548 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_8[2]\, B => 
        HIEFFPLA_NET_0_119575, S => HIEFFPLA_NET_0_119291, Y => 
        HIEFFPLA_NET_0_119725);
    
    HIEFFPLA_INST_0_57444 : NAND2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_4[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_4[2]\, Y => 
        HIEFFPLA_NET_0_116681);
    
    \U50_PATTERNS/ELINK_DINA_17[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119805, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_19, Q => 
        \U50_PATTERNS/ELINK_DINA_17[2]\);
    
    HIEFFPLA_INST_0_42263 : AO18
      port map(A => HIEFFPLA_NET_0_119559, B => 
        \U50_PATTERNS/RD_USB_ADBUS[5]\, C => 
        \U50_PATTERNS/RD_USB_ADBUS[4]\, Y => 
        HIEFFPLA_NET_0_119587);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_12[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116547, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_10, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_12[1]\);
    
    \U50_PATTERNS/TFC_STRT_ADDR[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119171, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_13, Q => 
        \U50_PATTERNS/TFC_STRT_ADDR[1]\);
    
    HIEFFPLA_INST_0_59594 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_13[2]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_29[2]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[4]_net_1\, Y => 
        HIEFFPLA_NET_0_116373);
    
    HIEFFPLA_INST_0_47804 : MX2
      port map(A => HIEFFPLA_NET_0_118429, B => 
        HIEFFPLA_NET_0_118454, S => \BIT_OS_SEL_2[1]\, Y => 
        HIEFFPLA_NET_0_118431);
    
    HIEFFPLA_INST_0_45971 : NAND3C
      port map(A => HIEFFPLA_NET_0_118944, B => 
        HIEFFPLA_NET_0_118954, C => HIEFFPLA_NET_0_118699, Y => 
        HIEFFPLA_NET_0_118799);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_26[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116404, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_21, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_26[2]\);
    
    \U_ELK1_CH/U_SLAVE_1ELK/RECD_SER_WORD[2]\ : DFN1C0
      port map(D => \U_ELK1_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[2]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_1[2]\);
    
    HIEFFPLA_INST_0_37252 : NOR3B
      port map(A => HIEFFPLA_NET_0_120268, B => 
        HIEFFPLA_NET_0_120273, C => HIEFFPLA_NET_0_120313, Y => 
        HIEFFPLA_NET_0_120314);
    
    \U200A_TFC/RX_SER_WORD_1DEL[1]\ : DFN1C0
      port map(D => \TFC_RX_SER_WORD[1]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_30, Q => 
        \U200A_TFC/RX_SER_WORD_1DEL[1]_net_1\);
    
    HIEFFPLA_INST_0_49865 : AND2A
      port map(A => \OP_MODE_c_1[1]\, B => \PATT_ELK_DAT_4[5]\, Y
         => HIEFFPLA_NET_0_118053);
    
    HIEFFPLA_INST_0_47764 : MX2
      port map(A => HIEFFPLA_NET_0_118440, B => 
        HIEFFPLA_NET_0_118453, S => \BIT_OS_SEL_4[0]\, Y => 
        \U_ELK14_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[3]\);
    
    HIEFFPLA_INST_0_40522 : MX2
      port map(A => HIEFFPLA_NET_0_119578, B => 
        \U50_PATTERNS/ELINK_DINA_13[0]\, S => 
        HIEFFPLA_NET_0_119285, Y => HIEFFPLA_NET_0_119839);
    
    HIEFFPLA_INST_0_48222 : MX2
      port map(A => HIEFFPLA_NET_0_118357, B => 
        HIEFFPLA_NET_0_118353, S => \BIT_OS_SEL_2[1]\, Y => 
        HIEFFPLA_NET_0_118351);
    
    \U50_PATTERNS/ELINK_RWA[4]/U1\ : DFN1P0
      port map(D => HIEFFPLA_NET_0_119697, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_6, Q => \U50_PATTERNS/ELINK_RWA[4]\);
    
    \U50_PATTERNS/ELINK_DINA_13[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119838, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_14, Q => 
        \U50_PATTERNS/ELINK_DINA_13[1]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_4[7]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116689, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_9, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_4[7]\);
    
    HIEFFPLA_INST_0_52430 : MX2
      port map(A => HIEFFPLA_NET_0_117516, B => 
        HIEFFPLA_NET_0_117512, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[3]\, Y => 
        HIEFFPLA_NET_0_117564);
    
    HIEFFPLA_INST_0_42710 : XNOR2
      port map(A => \U50_PATTERNS/REG_STATE[0]_net_1\, B => 
        \U50_PATTERNS/REG_STATE_0[2]_net_1\, Y => 
        HIEFFPLA_NET_0_119477);
    
    \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[78]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117703, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_34, Q => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[78]_net_1\);
    
    \U_ELK4_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]\ : DFN1C0
      port map(D => \U_ELK4_CH/U_SLAVE_1ELK/Q[0]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]_net_1\);
    
    HIEFFPLA_INST_0_41512 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_7[6]\, B => 
        HIEFFPLA_NET_0_119566, S => HIEFFPLA_NET_0_119289, Y => 
        HIEFFPLA_NET_0_119729);
    
    HIEFFPLA_INST_0_42868 : NAND2
      port map(A => \U50_PATTERNS/REG_STATE[2]_net_1\, B => 
        \U50_PATTERNS/REG_STATE[3]_net_1\, Y => 
        HIEFFPLA_NET_0_119442);
    
    HIEFFPLA_INST_0_37321 : AO1E
      port map(A => \OP_MODE_c[2]\, B => HIEFFPLA_NET_0_120293, C
         => \U200A_TFC/GP_PG_SM[2]_net_1\, Y => 
        HIEFFPLA_NET_0_120295);
    
    \U_ELK13_CH/U_ELK1_SERDAT_SOURCE/SERDAT[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118508, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_4, Q => 
        \U_ELK13_CH/ELK_TX_DAT[0]\);
    
    HIEFFPLA_INST_0_48889 : MX2
      port map(A => HIEFFPLA_NET_0_118219, B => 
        HIEFFPLA_NET_0_118215, S => \BIT_OS_SEL_0[1]\, Y => 
        HIEFFPLA_NET_0_118228);
    
    HIEFFPLA_INST_0_59281 : AND2
      port map(A => HIEFFPLA_NET_0_116740, B => 
        HIEFFPLA_NET_0_117394, Y => HIEFFPLA_NET_0_116410);
    
    HIEFFPLA_INST_0_54857 : AO1A
      port map(A => \OP_MODE_c[5]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_0[8]_net_1\, C => 
        HIEFFPLA_NET_0_115917, Y => HIEFFPLA_NET_0_117188);
    
    \U_ELK4_CH/U_SLAVE_1ELK/RECD_SER_WORD[1]\ : DFN1C0
      port map(D => \U_ELK4_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[1]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_4[1]\);
    
    \U_ELK11_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118605, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_11, Q => 
        \U_ELK11_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]_net_1\);
    
    \U50_PATTERNS/ELINK_DINA_2[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119768, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_9, Q => 
        \U50_PATTERNS/ELINK_DINA_2[7]\);
    
    HIEFFPLA_INST_0_56539 : AND3A
      port map(A => HIEFFPLA_NET_0_117430, B => \BIT_OS_SEL_1[2]\, 
        C => \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[11]_net_1\, 
        Y => HIEFFPLA_NET_0_116843);
    
    HIEFFPLA_INST_0_51234 : MX2
      port map(A => HIEFFPLA_NET_0_117824, B => 
        HIEFFPLA_NET_0_117822, S => \BIT_OS_SEL_4[0]\, Y => 
        \U_ELK9_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[1]\);
    
    \U_ELK13_CH/ELK_IN_R\ : DFN1C0
      port map(D => \U_ELK13_CH/ELK_IN_DDR_R\, CLK => 
        CCC_160M_ADJ, CLR => DEV_RST_B_c, Q => 
        \U_ELK13_CH/ELK_IN_R_net_1\);
    
    HIEFFPLA_INST_0_45827 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_14[7]\, C => 
        \U50_PATTERNS/SM_BANK_SEL[5]\, Y => HIEFFPLA_NET_0_118830);
    
    \U_EXEC_MASTER/CCC_1_LOCK_STAT_1D\ : DFN1C0
      port map(D => \U_EXEC_MASTER/CCC_1_LOCK_STAT_0D_net_1\, CLK
         => CLK_40M_GL, CLR => 
        \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i\, Q => 
        \U_EXEC_MASTER/CCC_1_LOCK_STAT_1D_net_1\);
    
    HIEFFPLA_INST_0_37429 : MX2
      port map(A => \U200A_TFC/LOC_STOP_ADDR[4]\, B => 
        \TFC_STOP_ADDR[4]\, S => \U200A_TFC/GP_PG_SM_0[10]_net_1\, 
        Y => HIEFFPLA_NET_0_120286);
    
    HIEFFPLA_INST_0_37304 : AO1D
      port map(A => \OP_MODE_c[2]\, B => HIEFFPLA_NET_0_120293, C
         => HIEFFPLA_NET_0_120329, Y => HIEFFPLA_NET_0_120299);
    
    \U_ELK15_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL\ : DFN1C0
      port map(D => \U_ELK15_CH/ELK_IN_R_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL_net_1\);
    
    \U_ELK0_CMD_TX/SER_CMD_WORD_R[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118664, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_14, Q => 
        \U_ELK0_CMD_TX/SER_CMD_WORD_R[1]_net_1\);
    
    HIEFFPLA_INST_0_39524 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_4[2]\, B => 
        HIEFFPLA_NET_0_119522, S => HIEFFPLA_NET_0_119284, Y => 
        HIEFFPLA_NET_0_119981);
    
    HIEFFPLA_INST_0_60866 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_17[0]\, B => 
        HIEFFPLA_NET_0_117190, S => HIEFFPLA_NET_0_117169, Y => 
        HIEFFPLA_NET_0_116205);
    
    \U_ELK10_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]\ : DFN1C0
      port map(D => \U_ELK10_CH/U_SLAVE_1ELK/Q[13]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]_net_1\);
    
    HIEFFPLA_INST_0_42642 : AND3
      port map(A => HIEFFPLA_NET_0_119400, B => 
        HIEFFPLA_NET_0_119371, C => 
        \U50_PATTERNS/REG_STATE_0[1]_net_1\, Y => 
        HIEFFPLA_NET_0_119493);
    
    \U_ELK18_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]\ : DFN1C0
      port map(D => \U_ELK18_CH/U_SLAVE_1ELK/Q[13]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]_net_1\);
    
    HIEFFPLA_INST_0_111349 : NAND3C
      port map(A => HIEFFPLA_NET_0_116806, B => 
        HIEFFPLA_NET_0_116742, C => HIEFFPLA_NET_0_116687, Y => 
        HIEFFPLA_NET_0_115840);
    
    \U_ELK5_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL\ : DFN1C0
      port map(D => 
        \U_ELK5_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL_net_1\);
    
    \U_ELK4_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]\ : DFN1C0
      port map(D => \U_ELK4_CH/U_SLAVE_1ELK/Q[12]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]_net_1\);
    
    \U50_PATTERNS/ELINK_ADDRA_17[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120026, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_11, Q => 
        \U50_PATTERNS/ELINK_ADDRA_17[5]\);
    
    HIEFFPLA_INST_0_55444 : MX2
      port map(A => HIEFFPLA_NET_0_116979, B => 
        HIEFFPLA_NET_0_117032, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[2]\, Y => 
        HIEFFPLA_NET_0_117036);
    
    \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[3]\ : DFN1C0
      port map(D => 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[3]_net_1\);
    
    HIEFFPLA_INST_0_51651 : AND2A
      port map(A => HIEFFPLA_NET_0_117753, B => 
        \U_EXEC_MASTER/USB_MASTER_EN/CNT_EN_60M2S_net_1\, Y => 
        HIEFFPLA_NET_0_117731);
    
    \U50_PATTERNS/U113_PATT_ELINK_BLK/DPRT_512X9_SRAM_R0C0\ : 
        RAM4K9
      generic map(MEMORYFILE => "DPRT_512X9_SRAM_R0C0.mem")

      port map(ADDRA11 => AFLSDF_GND, ADDRA10 => AFLSDF_GND, 
        ADDRA9 => AFLSDF_GND, ADDRA8 => \GND\, ADDRA7 => 
        \U50_PATTERNS/ELINK_ADDRA_13[7]\, ADDRA6 => 
        \U50_PATTERNS/ELINK_ADDRA_13[6]\, ADDRA5 => 
        \U50_PATTERNS/ELINK_ADDRA_13[5]\, ADDRA4 => 
        \U50_PATTERNS/ELINK_ADDRA_13[4]\, ADDRA3 => 
        \U50_PATTERNS/ELINK_ADDRA_13[3]\, ADDRA2 => 
        \U50_PATTERNS/ELINK_ADDRA_13[2]\, ADDRA1 => 
        \U50_PATTERNS/ELINK_ADDRA_13[1]\, ADDRA0 => 
        \U50_PATTERNS/ELINK_ADDRA_13[0]\, ADDRB11 => AFLSDF_GND, 
        ADDRB10 => AFLSDF_GND, ADDRB9 => AFLSDF_GND, ADDRB8 => 
        \GND\, ADDRB7 => \ELKS_ADDRB[7]\, ADDRB6 => 
        \ELKS_ADDRB_0[6]\, ADDRB5 => \ELKS_ADDRB[5]\, ADDRB4 => 
        \ELKS_ADDRB_0[4]\, ADDRB3 => \ELKS_ADDRB[3]\, ADDRB2 => 
        \ELKS_ADDRB_0[2]\, ADDRB1 => \ELKS_ADDRB[1]\, ADDRB0 => 
        \ELKS_ADDRB[0]\, DINA8 => \GND\, DINA7 => 
        \U50_PATTERNS/ELINK_DINA_13[7]\, DINA6 => 
        \U50_PATTERNS/ELINK_DINA_13[6]\, DINA5 => 
        \U50_PATTERNS/ELINK_DINA_13[5]\, DINA4 => 
        \U50_PATTERNS/ELINK_DINA_13[4]\, DINA3 => 
        \U50_PATTERNS/ELINK_DINA_13[3]\, DINA2 => 
        \U50_PATTERNS/ELINK_DINA_13[2]\, DINA1 => 
        \U50_PATTERNS/ELINK_DINA_13[1]\, DINA0 => 
        \U50_PATTERNS/ELINK_DINA_13[0]\, DINB8 => \GND\, DINB7
         => \ELK_RX_SER_WORD_13[7]\, DINB6 => 
        \ELK_RX_SER_WORD_13[6]\, DINB5 => \ELK_RX_SER_WORD_13[5]\, 
        DINB4 => \ELK_RX_SER_WORD_13[4]\, DINB3 => 
        \ELK_RX_SER_WORD_13[3]\, DINB2 => \ELK_RX_SER_WORD_13[2]\, 
        DINB1 => \ELK_RX_SER_WORD_13[1]\, DINB0 => 
        \ELK_RX_SER_WORD_13[0]\, WIDTHA0 => \VCC\, WIDTHA1 => 
        \VCC\, WIDTHB0 => \VCC\, WIDTHB1 => \VCC\, PIPEA => \VCC\, 
        PIPEB => \VCC\, WMODEA => \GND\, WMODEB => \GND\, BLKA
         => \U50_PATTERNS/ELINK_BLKA[13]\, BLKB => 
        ELKS_RAM_BLKB_EN, WENA => \U50_PATTERNS/ELINK_RWA[13]\, 
        WENB => ELKS_RWB, CLKA => CLK60MHZ, CLKB => CLK_40M_GL, 
        RESET => P_USB_MASTER_EN_c_0, DOUTA8 => OPEN, DOUTA7 => 
        \U50_PATTERNS/ELINK_DOUTA_13[7]\, DOUTA6 => 
        \U50_PATTERNS/ELINK_DOUTA_13[6]\, DOUTA5 => 
        \U50_PATTERNS/ELINK_DOUTA_13[5]\, DOUTA4 => 
        \U50_PATTERNS/ELINK_DOUTA_13[4]\, DOUTA3 => 
        \U50_PATTERNS/ELINK_DOUTA_13[3]\, DOUTA2 => 
        \U50_PATTERNS/ELINK_DOUTA_13[2]\, DOUTA1 => 
        \U50_PATTERNS/ELINK_DOUTA_13[1]\, DOUTA0 => 
        \U50_PATTERNS/ELINK_DOUTA_13[0]\, DOUTB8 => OPEN, DOUTB7
         => \PATT_ELK_DAT_13[7]\, DOUTB6 => \PATT_ELK_DAT_13[6]\, 
        DOUTB5 => \PATT_ELK_DAT_13[5]\, DOUTB4 => 
        \PATT_ELK_DAT_13[4]\, DOUTB3 => \PATT_ELK_DAT_13[3]\, 
        DOUTB2 => \PATT_ELK_DAT_13[2]\, DOUTB1 => 
        \PATT_ELK_DAT_13[1]\, DOUTB0 => \PATT_ELK_DAT_13[0]\);
    
    \U_ELK3_CH/U_ELK1_SERDAT_SOURCE/SERDAT[5]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118098, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_15, Q => 
        \U_ELK3_CH/ELK_TX_DAT[5]\);
    
    HIEFFPLA_INST_0_62723 : XNOR3
      port map(A => HIEFFPLA_NET_0_115955, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_CLKPHASE[3]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_SEQCNT[4]\, Y => 
        HIEFFPLA_NET_0_115953);
    
    HIEFFPLA_INST_0_43897 : AO1D
      port map(A => HIEFFPLA_NET_0_119389, B => 
        HIEFFPLA_NET_0_119464, C => 
        \U50_PATTERNS/SM_BANK_SEL_0[21]\, Y => 
        HIEFFPLA_NET_0_119198);
    
    HIEFFPLA_INST_0_57615 : NAND2B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_5[4]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_5[5]\, Y => 
        HIEFFPLA_NET_0_116652);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_1[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116168, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_8, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_1[2]\);
    
    \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[9]\ : DFN1C0
      port map(D => 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\);
    
    \U_ELK3_CH/U_ELK1_CMD_TX/SER_OUT_FDEL\ : DFN1P0
      port map(D => \U_ELK3_CH/U_ELK1_CMD_TX/SER_OUT_FI_i\, CLK
         => CCC_160M_FXD, PRE => MASTER_SALT_POR_B_i_0_i_5, Q => 
        \U_ELK3_CH/ELK_OUT_F_i_0\);
    
    HIEFFPLA_INST_0_60191 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_7[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_23[1]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_4[4]_net_1\, Y
         => HIEFFPLA_NET_0_116298);
    
    HIEFFPLA_INST_0_58701 : AND2
      port map(A => HIEFFPLA_NET_0_116740, B => 
        HIEFFPLA_NET_0_117204, Y => HIEFFPLA_NET_0_116485);
    
    HIEFFPLA_INST_0_58225 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_12[0]\, B => 
        HIEFFPLA_NET_0_116680, S => HIEFFPLA_NET_0_117089, Y => 
        HIEFFPLA_NET_0_116548);
    
    HIEFFPLA_INST_0_56279 : NAND3C
      port map(A => HIEFFPLA_NET_0_116877, B => 
        HIEFFPLA_NET_0_116885, C => HIEFFPLA_NET_0_116893, Y => 
        HIEFFPLA_NET_0_116901);
    
    HIEFFPLA_INST_0_54261 : MX2
      port map(A => HIEFFPLA_NET_0_116150, B => 
        HIEFFPLA_NET_0_116050, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_2[3]_net_1\, Y
         => HIEFFPLA_NET_0_117288);
    
    \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_115941, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_24_0, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[1]_net_1\);
    
    HIEFFPLA_INST_0_61109 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_3[4]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_19[4]\, S
         => \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_1[4]_net_1\, 
        Y => HIEFFPLA_NET_0_116172);
    
    \U_ELK13_CH/U_SLAVE_1ELK/RECD_SER_WORD[7]\ : DFN1C0
      port map(D => \U_ELK13_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[7]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_13[7]\);
    
    HIEFFPLA_INST_0_49393 : MX2
      port map(A => HIEFFPLA_NET_0_118138, B => 
        HIEFFPLA_NET_0_118135, S => \BIT_OS_SEL[1]\, Y => 
        HIEFFPLA_NET_0_118137);
    
    HIEFFPLA_INST_0_52618 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_5[2]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_6[2]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_2[0]\, Y => 
        HIEFFPLA_NET_0_117538);
    
    HIEFFPLA_INST_0_58485 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_31[0]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_15[0]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_3[4]_net_1\, Y
         => HIEFFPLA_NET_0_116516);
    
    HIEFFPLA_INST_0_54914 : AOI1C
      port map(A => HIEFFPLA_NET_0_117184, B => 
        HIEFFPLA_NET_0_117388, C => HIEFFPLA_NET_0_117218, Y => 
        HIEFFPLA_NET_0_117171);
    
    HIEFFPLA_INST_0_46345 : NAND3C
      port map(A => HIEFFPLA_NET_0_118858, B => 
        HIEFFPLA_NET_0_118863, C => HIEFFPLA_NET_0_118868, Y => 
        HIEFFPLA_NET_0_118711);
    
    HIEFFPLA_INST_0_37976 : MX2
      port map(A => \U200B_ELINKS/LOC_STOP_ADDR[7]\, B => 
        \ELKS_STOP_ADDR[7]\, S => 
        \U200B_ELINKS/GP_PG_SM_0[10]_net_1\, Y => 
        HIEFFPLA_NET_0_120180);
    
    \U_ELK18_CH/U_SLAVE_1ELK/Q[11]\ : DFN1C0
      port map(D => \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/Q[11]_net_1\);
    
    HIEFFPLA_INST_0_56240 : AND2
      port map(A => DCB_SALT_SEL_c, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/RECD_SER_WORD[3]_net_1\, 
        Y => \ELK_RX_SER_WORD_0[3]\);
    
    HIEFFPLA_INST_0_40864 : MX2
      port map(A => HIEFFPLA_NET_0_119566, B => 
        \U50_PATTERNS/ELINK_DINA_17[6]\, S => 
        HIEFFPLA_NET_0_119260, Y => HIEFFPLA_NET_0_119801);
    
    \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[5]\ : DFN1C0
      port map(D => \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\);
    
    HIEFFPLA_INST_0_62110 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_2[1]\, 
        B => HIEFFPLA_NET_0_117167, S => HIEFFPLA_NET_0_117176, Y
         => HIEFFPLA_NET_0_116034);
    
    HIEFFPLA_INST_0_53348 : MX2
      port map(A => HIEFFPLA_NET_0_117278, B => 
        HIEFFPLA_NET_0_117268, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[2]_net_1\, Y
         => HIEFFPLA_NET_0_117421);
    
    \U50_PATTERNS/RD_XFER_TYPE[5]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119544, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c, Q => 
        \U50_PATTERNS/RD_XFER_TYPE[5]_net_1\);
    
    HIEFFPLA_INST_0_53335 : AND2A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_SEL[3]_net_1\, B
         => \BIT_OS_SEL[2]\, Y => HIEFFPLA_NET_0_117424);
    
    \U_ELK5_CH/U_ELK1_CMD_TX/SER_OUT_RI\ : DFN1C0
      port map(D => 
        \U_ELK5_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_14, Q
         => \U_ELK5_CH/U_ELK1_CMD_TX/SER_OUT_RI_net_1\);
    
    \U_ELK3_CH/U_SLAVE_1ELK/RECD_SER_WORD[1]\ : DFN1C0
      port map(D => \U_ELK3_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[1]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_3[1]\);
    
    \U50_PATTERNS/U4A_REGCROSS/SAMP_ONE[6]\ : DFN1C0
      port map(D => \U50_PATTERNS/TFC_STRT_ADDR[6]\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_32_0, Q => 
        \U50_PATTERNS/U4A_REGCROSS/SAMP_ONE[6]_net_1\);
    
    \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[13]\ : DFN1C0
      port map(D => \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\, 
        CLK => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[13]_net_1\);
    
    \U50_PATTERNS/U4B_REGCROSS/SAMP_ONE[3]\ : DFN1C0
      port map(D => \U50_PATTERNS/TFC_STOP_ADDR[3]\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_25, Q => 
        \U50_PATTERNS/U4B_REGCROSS/SAMP_ONE[3]_net_1\);
    
    HIEFFPLA_INST_0_50162 : MX2
      port map(A => \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\, B
         => \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\, S => 
        \BIT_OS_SEL_6[2]\, Y => HIEFFPLA_NET_0_117999);
    
    \U_ELK1_CH/U_ELK1_CMD_TX/SER_OUT_RI\ : DFI1C0
      port map(D => 
        \U_ELK1_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_14, QN
         => \U_ELK1_CH/U_ELK1_CMD_TX/SER_OUT_RI_i\);
    
    \U_ELK13_CH/U_SLAVE_1ELK/Q[6]\ : DFN1C0
      port map(D => \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/Q[6]_net_1\);
    
    \U_ELK11_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]\ : DFN1C0
      port map(D => \U_ELK11_CH/U_SLAVE_1ELK/Q[12]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]_net_1\);
    
    \U50_PATTERNS/WR_USB_ADBUS[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118980, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_15, Q => 
        \U50_PATTERNS/WR_USB_ADBUS[5]\);
    
    HIEFFPLA_INST_0_52990 : MX2
      port map(A => HIEFFPLA_NET_0_117463, B => 
        HIEFFPLA_NET_0_117459, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[2]\, Y => 
        HIEFFPLA_NET_0_117479);
    
    HIEFFPLA_INST_0_40513 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_12[7]\, B => 
        HIEFFPLA_NET_0_119560, S => HIEFFPLA_NET_0_119295, Y => 
        HIEFFPLA_NET_0_119840);
    
    \U50_PATTERNS/ELINK_DINA_2[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119774, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_9, Q => 
        \U50_PATTERNS/ELINK_DINA_2[1]\);
    
    HIEFFPLA_INST_0_57953 : NAND2A
      port map(A => HIEFFPLA_NET_0_116589, B => 
        HIEFFPLA_NET_0_116620, Y => HIEFFPLA_NET_0_116593);
    
    HIEFFPLA_INST_0_52278 : AND3A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[6]_net_1\, B => 
        HIEFFPLA_NET_0_117606, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[1]_net_1\, Y => 
        HIEFFPLA_NET_0_117592);
    
    HIEFFPLA_INST_0_48626 : MX2
      port map(A => HIEFFPLA_NET_0_118265, B => 
        HIEFFPLA_NET_0_118262, S => \BIT_OS_SEL_1[1]\, Y => 
        HIEFFPLA_NET_0_118275);
    
    \P_OP_MODE5_AAE_pad/U0/U0\ : IOPAD_TRI_U
      port map(D => \P_OP_MODE5_AAE_pad/U0/NET1\, E => 
        \P_OP_MODE5_AAE_pad/U0/NET2\, PAD => P_OP_MODE5_AAE);
    
    HIEFFPLA_INST_0_56186 : XA1C
      port map(A => HIEFFPLA_NET_0_116940, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/MAX_CNT[5]\, C => 
        HIEFFPLA_NET_0_117112, Y => HIEFFPLA_NET_0_116934);
    
    HIEFFPLA_INST_0_44938 : MX2
      port map(A => USB_SIWU_BI, B => HIEFFPLA_NET_0_119329, S
         => HIEFFPLA_NET_0_119443, Y => HIEFFPLA_NET_0_119013);
    
    HIEFFPLA_INST_0_39959 : MX2
      port map(A => HIEFFPLA_NET_0_119909, B => 
        \U50_PATTERNS/ELINK_BLKA[12]\, S => 
        \U50_PATTERNS/SM_BANK_SEL[20]\, Y => 
        HIEFFPLA_NET_0_119932);
    
    HIEFFPLA_INST_0_48866 : NAND2B
      port map(A => \OP_MODE_c_5[1]\, B => \PATT_ELK_DAT_19[2]\, 
        Y => HIEFFPLA_NET_0_118236);
    
    HIEFFPLA_INST_0_54721 : AND3
      port map(A => HIEFFPLA_NET_0_117236, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[0]_net_1\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[3]_net_1\, Y => 
        HIEFFPLA_NET_0_117217);
    
    \P_MASTER_POR_B_pad/U0/U0\ : IOPAD_TRI_U
      port map(D => \P_MASTER_POR_B_pad/U0/NET1\, E => 
        \P_MASTER_POR_B_pad/U0/NET2\, PAD => P_MASTER_POR_B);
    
    HIEFFPLA_INST_0_37616 : XO1A
      port map(A => HIEFFPLA_NET_0_120226, B => \ELKS_ADDRB[0]\, 
        C => \U200B_ELINKS/GP_PG_SM[10]_net_1\, Y => 
        HIEFFPLA_NET_0_120246);
    
    \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[4]\ : DFN1C0
      port map(D => \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\);
    
    \U_ELK4_CH/U_ELK1_CMD_TX/SER_OUT_RDEL\ : DFN1P0
      port map(D => \U_ELK4_CH/U_ELK1_CMD_TX/SER_OUT_RI_i\, CLK
         => CCC_160M_FXD, PRE => MASTER_SALT_POR_B_i_0_i_13, Q
         => \U_ELK4_CH/ELK_OUT_R_i_0\);
    
    \U_ELK18_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2\ : IOPADN_BI
      port map(DB => \U_ELK18_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, 
        E => \U_ELK18_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET3\, PAD
         => ELK18_DAT_N, N2POUT => 
        \U_ELK18_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2_N2P\);
    
    \U_ELK12_CH/U_SLAVE_1ELK/Q[8]\ : DFN1C0
      port map(D => \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/Q[8]_net_1\);
    
    HIEFFPLA_INST_0_58634 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_18[0]\, B => 
        HIEFFPLA_NET_0_116491, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_2[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116495);
    
    HIEFFPLA_INST_0_59751 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_30[3]\, B => 
        HIEFFPLA_NET_0_116347, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_2[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116353);
    
    HIEFFPLA_INST_0_47620 : NAND2B
      port map(A => \OP_MODE_c_2[1]\, B => \PATT_ELK_DAT_14[1]\, 
        Y => HIEFFPLA_NET_0_118462);
    
    \U50_PATTERNS/U4C_REGCROSS/SYNC_SM[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119104, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_32, Q => 
        \U50_PATTERNS/U4C_REGCROSS/SYNC_SM[0]_net_1\);
    
    \U_ELK2_CH/U_SLAVE_1ELK/RECD_SER_WORD[7]\ : DFN1C0
      port map(D => \U_ELK2_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[7]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_2[7]\);
    
    \U_ELK12_CH/U_ELK1_SERDAT_SOURCE/SERDAT[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118553, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_2, Q => 
        \U_ELK12_CH/ELK_TX_DAT[0]\);
    
    \U_DDR_TFC/BIBUF_LVDS_0/U0/U2\ : IOPADN_BI
      port map(DB => \U_DDR_TFC/BIBUF_LVDS_0/U0/NET1\, E => 
        \U_DDR_TFC/BIBUF_LVDS_0/U0/NET3\, PAD => TFC_DAT_0N, 
        N2POUT => \U_DDR_TFC/BIBUF_LVDS_0/U0/U2_N2P\);
    
    HIEFFPLA_INST_0_58893 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_4[0]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_20[0]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_2[4]_net_1\, Y
         => HIEFFPLA_NET_0_116462);
    
    HIEFFPLA_INST_0_55348 : AND3
      port map(A => HIEFFPLA_NET_0_117104, B => 
        HIEFFPLA_NET_0_117048, C => HIEFFPLA_NET_0_115910, Y => 
        HIEFFPLA_NET_0_117054);
    
    HIEFFPLA_INST_0_61265 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_19[4]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_20[4]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_4[0]\, Y => 
        HIEFFPLA_NET_0_116151);
    
    HIEFFPLA_INST_0_44991 : AO1
      port map(A => \U50_PATTERNS/USB_TXE_B\, B => 
        HIEFFPLA_NET_0_119381, C => HIEFFPLA_NET_0_119457, Y => 
        HIEFFPLA_NET_0_119005);
    
    HIEFFPLA_INST_0_60792 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_31[4]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_15[4]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[4]_net_1\, Y
         => HIEFFPLA_NET_0_116219);
    
    HIEFFPLA_INST_0_53304 : AND2A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_0[8]_net_1\, B => 
        HIEFFPLA_NET_0_116976, Y => HIEFFPLA_NET_0_117436);
    
    HIEFFPLA_INST_0_54397 : MX2
      port map(A => HIEFFPLA_NET_0_116210, B => 
        HIEFFPLA_NET_0_116100, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_2[3]_net_1\, Y
         => HIEFFPLA_NET_0_117271);
    
    HIEFFPLA_INST_0_45497 : AND3A
      port map(A => HIEFFPLA_NET_0_119437, B => 
        \U50_PATTERNS/WR_XFER_TYPE[3]_net_1\, C => 
        HIEFFPLA_NET_0_119367, Y => HIEFFPLA_NET_0_118902);
    
    HIEFFPLA_INST_0_38118 : AX1C
      port map(A => \ELKS_ADDRB[4]\, B => HIEFFPLA_NET_0_120146, 
        C => \ELKS_ADDRB[5]\, Y => HIEFFPLA_NET_0_120148);
    
    HIEFFPLA_INST_0_45407 : NAND2A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_9[4]\, Y => 
        HIEFFPLA_NET_0_118919);
    
    HIEFFPLA_INST_0_62977 : MX2
      port map(A => HIEFFPLA_NET_0_115886, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[8]\, S => 
        HIEFFPLA_NET_0_117073, Y => HIEFFPLA_NET_0_115922);
    
    HIEFFPLA_INST_0_45882 : AO1
      port map(A => HIEFFPLA_NET_0_119246, B => 
        \U50_PATTERNS/ELINK_DOUTA_3[7]\, C => 
        HIEFFPLA_NET_0_118774, Y => HIEFFPLA_NET_0_118821);
    
    HIEFFPLA_INST_0_43050 : AO1
      port map(A => HIEFFPLA_NET_0_119453, B => 
        HIEFFPLA_NET_0_119373, C => HIEFFPLA_NET_0_119383, Y => 
        HIEFFPLA_NET_0_119391);
    
    HIEFFPLA_INST_0_41688 : MX2
      port map(A => HIEFFPLA_NET_0_119689, B => 
        \U50_PATTERNS/ELINK_RWA[11]\, S => 
        \U50_PATTERNS/SM_BANK_SEL_0[20]\, Y => 
        HIEFFPLA_NET_0_119709);
    
    \U_ELK10_CH/U_SLAVE_1ELK/RECD_SER_WORD[6]\ : DFN1C0
      port map(D => \U_ELK10_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[6]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_10[6]\);
    
    HIEFFPLA_INST_0_50471 : MX2
      port map(A => HIEFFPLA_NET_0_117957, B => 
        HIEFFPLA_NET_0_117954, S => \BIT_OS_SEL_5[1]\, Y => 
        HIEFFPLA_NET_0_117945);
    
    \U50_PATTERNS/REG_ADDR[8]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119525, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_10, Q => \U50_PATTERNS/REG_ADDR[8]\);
    
    HIEFFPLA_INST_0_63102 : XA1B
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[6]\, 
        B => HIEFFPLA_NET_0_115881, C => HIEFFPLA_NET_0_117078, Y
         => HIEFFPLA_NET_0_115888);
    
    HIEFFPLA_INST_0_56401 : NAND3C
      port map(A => HIEFFPLA_NET_0_116828, B => 
        HIEFFPLA_NET_0_116844, C => HIEFFPLA_NET_0_116852, Y => 
        HIEFFPLA_NET_0_116876);
    
    HIEFFPLA_INST_0_39533 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_4[3]\, B => 
        HIEFFPLA_NET_0_119520, S => HIEFFPLA_NET_0_119284, Y => 
        HIEFFPLA_NET_0_119980);
    
    HIEFFPLA_INST_0_39236 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_19[2]\, B => 
        HIEFFPLA_NET_0_119522, S => HIEFFPLA_NET_0_119293, Y => 
        HIEFFPLA_NET_0_120013);
    
    \U_EXEC_MASTER/MPOR_B_1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117787, CLK => CLK_40M_GL, CLR
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_2\, Q => 
        P_MASTER_POR_B_c_1);
    
    HIEFFPLA_INST_0_50294 : MX2
      port map(A => HIEFFPLA_NET_0_117979, B => 
        HIEFFPLA_NET_0_118001, S => \BIT_OS_SEL_5[1]\, Y => 
        HIEFFPLA_NET_0_117981);
    
    \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[7]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[5]_net_1\, CLK => 
        CCC_160M_ADJ, CLR => P_MASTER_POR_B_c_34_0, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[7]_net_1\);
    
    HIEFFPLA_INST_0_49708 : MX2
      port map(A => HIEFFPLA_NET_0_118089, B => 
        HIEFFPLA_NET_0_118087, S => \BIT_OS_SEL[1]\, Y => 
        HIEFFPLA_NET_0_118082);
    
    HIEFFPLA_INST_0_53899 : AND3A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[0]_net_1\, B
         => HIEFFPLA_NET_0_117236, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_1[3]_net_1\, Y
         => HIEFFPLA_NET_0_117337);
    
    HIEFFPLA_INST_0_61247 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_19[2]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_20[2]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_4[0]\, Y => 
        HIEFFPLA_NET_0_116154);
    
    HIEFFPLA_INST_0_45817 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/SM_BANK_SEL[18]\, C => 
        \U50_PATTERNS/ELINK_DOUTA_1[4]\, Y => 
        HIEFFPLA_NET_0_118833);
    
    HIEFFPLA_INST_0_51727 : NAND2B
      port map(A => 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM[4]_net_1\, B => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[9]_net_1\, Y => 
        HIEFFPLA_NET_0_117699);
    
    HIEFFPLA_INST_0_49582 : MX2
      port map(A => 
        \U_ELK3_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]_net_1\, B => 
        \U_ELK3_CH/ELK_TX_DAT[4]\, S => 
        \U_ELK3_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118110);
    
    HIEFFPLA_INST_0_46367 : AO1
      port map(A => HIEFFPLA_NET_0_119476, B => 
        \U50_PATTERNS/CHKSUM[6]\, C => HIEFFPLA_NET_0_118855, Y
         => HIEFFPLA_NET_0_118706);
    
    HIEFFPLA_INST_0_56410 : NAND3C
      port map(A => HIEFFPLA_NET_0_116825, B => 
        HIEFFPLA_NET_0_116841, C => HIEFFPLA_NET_0_116849, Y => 
        HIEFFPLA_NET_0_116873);
    
    \U_ELK18_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL\ : DFN1C0
      port map(D => \U_ELK18_CH/ELK_IN_R_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL_net_1\);
    
    HIEFFPLA_INST_0_51101 : MX2
      port map(A => HIEFFPLA_NET_0_117836, B => 
        \U_ELK9_CH/ELK_TX_DAT[7]\, S => 
        \U_ELK9_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_117835);
    
    HIEFFPLA_INST_0_111246 : MX2A
      port map(A => HIEFFPLA_NET_0_115847, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_7[3]\, S => 
        HIEFFPLA_NET_0_117212, Y => HIEFFPLA_NET_0_116294);
    
    \U_EXEC_MASTER/MPOR_SALT_B_15\ : DFI1P0
      port map(D => HIEFFPLA_NET_0_117781, CLK => CLK_40M_GL, PRE
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_2\, QN => 
        MASTER_SALT_POR_B_i_0_i_15);
    
    \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[6]\ : DFN1C0
      port map(D => \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\);
    
    HIEFFPLA_INST_0_54101 : MX2
      port map(A => HIEFFPLA_NET_0_117362, B => 
        HIEFFPLA_NET_0_117197, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[1]_net_1\, Y
         => HIEFFPLA_NET_0_117308);
    
    HIEFFPLA_INST_0_52564 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_1[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_2[1]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[0]\, Y => 
        HIEFFPLA_NET_0_117547);
    
    HIEFFPLA_INST_0_43455 : MX2
      port map(A => \U50_PATTERNS/SM_BANK_SEL[21]\, B => 
        HIEFFPLA_NET_0_119018, S => HIEFFPLA_NET_0_118691, Y => 
        HIEFFPLA_NET_0_119309);
    
    HIEFFPLA_INST_0_51770 : MX2
      port map(A => \U_MASTER_DES/U13A_ADJ_160M/BITCNT[4]\, B => 
        HIEFFPLA_NET_0_117678, S => HIEFFPLA_NET_0_117630, Y => 
        HIEFFPLA_NET_0_117694);
    
    \U_ELK9_CH/U_SLAVE_1ELK/RECD_SER_WORD[5]\ : DFN1C0
      port map(D => \U_ELK9_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[5]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_9[5]\);
    
    HIEFFPLA_INST_0_52770 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_3[2]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_4[2]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[0]\, Y => 
        HIEFFPLA_NET_0_117514);
    
    \U50_PATTERNS/ELINK_ADDRA_3[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119985, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_1, Q => 
        \U50_PATTERNS/ELINK_ADDRA_3[6]\);
    
    \U50_PATTERNS/ELINK_ADDRA_14[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120051, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_5, Q => 
        \U50_PATTERNS/ELINK_ADDRA_14[4]\);
    
    HIEFFPLA_INST_0_55232 : AO1A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[6]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[8]_net_1\, C => 
        HIEFFPLA_NET_0_117079, Y => HIEFFPLA_NET_0_117080);
    
    \U_ELK13_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]\ : DFN1C0
      port map(D => \U_ELK13_CH/U_SLAVE_1ELK/Q[3]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]_net_1\);
    
    \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[0]\ : DFN1C0
      port map(D => 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[0]_net_1\);
    
    HIEFFPLA_INST_0_62604 : MX2
      port map(A => HIEFFPLA_NET_0_117131, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_8[2]\, S => 
        HIEFFPLA_NET_0_117153, Y => HIEFFPLA_NET_0_115968);
    
    HIEFFPLA_INST_0_59662 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_2[2]\, B => 
        HIEFFPLA_NET_0_116359, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_1[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116365);
    
    HIEFFPLA_INST_0_37447 : MX2
      port map(A => \U200A_TFC/LOC_STOP_ADDR[7]\, B => 
        \TFC_STOP_ADDR[7]\, S => \U200A_TFC/GP_PG_SM_0[10]_net_1\, 
        Y => HIEFFPLA_NET_0_120283);
    
    \U_ELK3_CH/U_SLAVE_1ELK/RECD_SER_WORD[0]\ : DFN1C0
      port map(D => \U_ELK3_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[0]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_3[0]\);
    
    \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[0]\ : DFN1C0
      port map(D => 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[0]_net_1\);
    
    HIEFFPLA_INST_0_62265 : AND2A
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[0]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_31[2]\, Y
         => HIEFFPLA_NET_0_116013);
    
    HIEFFPLA_INST_0_48123 : AND2A
      port map(A => \OP_MODE_c_2[1]\, B => \PATT_ELK_DAT_16[6]\, 
        Y => HIEFFPLA_NET_0_118367);
    
    HIEFFPLA_INST_0_51174 : MX2
      port map(A => \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[3]_net_1\, B
         => \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\, S => 
        \BIT_OS_SEL_2[2]\, Y => HIEFFPLA_NET_0_117817);
    
    \U50_PATTERNS/U4B_REGCROSS/SAMP_TWO[5]\ : DFN1C0
      port map(D => \U50_PATTERNS/U4B_REGCROSS/SAMP_ONE[5]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_29, Q => 
        \U50_PATTERNS/U4B_REGCROSS/SAMP_TWO[5]_net_1\);
    
    HIEFFPLA_INST_0_52174 : MX2
      port map(A => 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM[5]_net_1\, B => 
        \U_MASTER_DES/CCC2_CONFIG_TRIG\, S => 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM[6]_net_1\, Y => 
        HIEFFPLA_NET_0_117616);
    
    HIEFFPLA_INST_0_48985 : MX2
      port map(A => HIEFFPLA_NET_0_118206, B => 
        HIEFFPLA_NET_0_118230, S => \BIT_OS_SEL_2[0]\, Y => 
        \U_ELK19_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[0]\);
    
    HIEFFPLA_INST_0_50407 : MX2
      port map(A => \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[2]_net_1\, B
         => \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\, S => 
        \BIT_OS_SEL_5[2]\, Y => HIEFFPLA_NET_0_117955);
    
    \U50_PATTERNS/ELINK_ADDRA_2[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119995, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_21, Q => 
        \U50_PATTERNS/ELINK_ADDRA_2[4]\);
    
    HIEFFPLA_INST_0_51152 : MX2
      port map(A => HIEFFPLA_NET_0_117811, B => 
        HIEFFPLA_NET_0_117825, S => \BIT_OS_SEL_3[1]\, Y => 
        HIEFFPLA_NET_0_117820);
    
    HIEFFPLA_INST_0_111348 : MX2A
      port map(A => HIEFFPLA_NET_0_115840, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_20[3]\, S => 
        HIEFFPLA_NET_0_117203, Y => HIEFFPLA_NET_0_116457);
    
    HIEFFPLA_INST_0_37229 : AOI1
      port map(A => \U200A_TFC/GP_PG_SM[0]_net_1\, B => 
        HIEFFPLA_NET_0_120309, C => HIEFFPLA_NET_0_120301, Y => 
        HIEFFPLA_NET_0_120319);
    
    \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[4]\\\\/U0/U0\ : 
        IOPAD_BI_U
      port map(D => 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[4]\\\\/U0/NET1\, 
        E => 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[4]\\\\/U0/NET2\, 
        Y => 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[4]\\\\/U0/NET3\, 
        PAD => BIDIR_USB_ADBUS(4));
    
    \U50_PATTERNS/ELINK_DINA_11[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119849, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_11, Q => 
        \U50_PATTERNS/ELINK_DINA_11[6]\);
    
    HIEFFPLA_INST_0_44126 : MX2
      port map(A => \U50_PATTERNS/TFC_STRT_ADDR[2]\, B => 
        \U50_PATTERNS/TFC_STRT_ADDR_T[2]\, S => 
        HIEFFPLA_NET_0_119472, Y => HIEFFPLA_NET_0_119170);
    
    HIEFFPLA_INST_0_48860 : MX2
      port map(A => 
        \U_ELK19_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]_net_1\, B => 
        \U_ELK19_CH/ELK_TX_DAT[7]\, S => 
        \U_ELK19_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118240);
    
    \U_ELK15_CH/U_ELK1_SERDAT_SOURCE/SERDAT[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118418, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_7, Q => 
        \U_ELK15_CH/ELK_TX_DAT[0]\);
    
    HIEFFPLA_INST_0_40001 : MX2
      port map(A => HIEFFPLA_NET_0_119899, B => 
        \U50_PATTERNS/ELINK_BLKA[18]\, S => 
        \U50_PATTERNS/SM_BANK_SEL[20]\, Y => 
        HIEFFPLA_NET_0_119926);
    
    HIEFFPLA_INST_0_37181 : AND3
      port map(A => HIEFFPLA_NET_0_120334, B => 
        HIEFFPLA_NET_0_120324, C => HIEFFPLA_NET_0_120332, Y => 
        HIEFFPLA_NET_0_120331);
    
    \U_ELK5_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]\ : DFN1C0
      port map(D => \U_ELK5_CH/U_SLAVE_1ELK/Q[14]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]_net_1\);
    
    \U200B_ELINKS/ADDR_POINTER_0[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120169, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_31_0, Q => \ELKS_ADDRB_0[2]\);
    
    HIEFFPLA_INST_0_63243 : AND2A
      port map(A => \OP_MODE_c_0[1]\, B => \PATT_TFC_DAT[6]\, Y
         => \U_TFC_SERDAT_SOURCE/N_SERDAT[6]\);
    
    HIEFFPLA_INST_0_59070 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_23[3]\, B => 
        HIEFFPLA_NET_0_116435, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_1[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116439);
    
    HIEFFPLA_INST_0_40756 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_16[2]\, B => 
        HIEFFPLA_NET_0_119575, S => HIEFFPLA_NET_0_119257, Y => 
        HIEFFPLA_NET_0_119813);
    
    \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[11]\ : DFN1C0
      port map(D => \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\);
    
    HIEFFPLA_INST_0_42292 : NAND3B
      port map(A => \U50_PATTERNS/RD_USB_ADBUS[3]\, B => 
        \U50_PATTERNS/RD_USB_ADBUS[2]\, C => 
        \U50_PATTERNS/RD_USB_ADBUS[5]\, Y => 
        HIEFFPLA_NET_0_119580);
    
    HIEFFPLA_INST_0_60178 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_7[3]\, B => 
        HIEFFPLA_NET_0_116294, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_0[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116300);
    
    HIEFFPLA_INST_0_52102 : AND2A
      port map(A => \U_MASTER_DES/U13A_ADJ_160M/BITCNT[4]\, B => 
        HIEFFPLA_NET_0_117668, Y => HIEFFPLA_NET_0_117636);
    
    \U50_PATTERNS/WR_USB_ADBUS[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118985, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_15, Q => 
        \U50_PATTERNS/WR_USB_ADBUS[0]\);
    
    \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[7]\ : DFN1C0
      port map(D => 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\);
    
    HIEFFPLA_INST_0_47710 : MX2
      port map(A => HIEFFPLA_NET_0_118454, B => 
        HIEFFPLA_NET_0_118451, S => \BIT_OS_SEL_2[1]\, Y => 
        HIEFFPLA_NET_0_118443);
    
    HIEFFPLA_INST_0_46475 : AOI1D
      port map(A => HIEFFPLA_NET_0_119571, B => 
        HIEFFPLA_NET_0_119583, C => 
        \U50_PATTERNS/WR_XFER_TYPE[5]_net_1\, Y => 
        HIEFFPLA_NET_0_118683);
    
    \U_ELK12_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL\ : DFN1C0
      port map(D => \U_ELK12_CH/ELK_IN_F_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL_net_1\);
    
    \U_ELK11_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]\ : DFN1C0
      port map(D => \U_ELK11_CH/U_SLAVE_1ELK/Q[14]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]_net_1\);
    
    HIEFFPLA_INST_0_47180 : MX2
      port map(A => HIEFFPLA_NET_0_118530, B => 
        HIEFFPLA_NET_0_118543, S => \BIT_OS_SEL_4[1]\, Y => 
        HIEFFPLA_NET_0_118538);
    
    HIEFFPLA_INST_0_51146 : MX2
      port map(A => \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[1]_net_1\, B
         => \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\, S => 
        \BIT_OS_SEL_2[2]\, Y => HIEFFPLA_NET_0_117821);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_31[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116340, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_20, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_31[3]\);
    
    \U50_PATTERNS/U117_PATT_ELINK_BLK/DPRT_512X9_SRAM_R0C0\ : 
        RAM4K9
      generic map(MEMORYFILE => "DPRT_512X9_SRAM_R0C0.mem")

      port map(ADDRA11 => AFLSDF_GND, ADDRA10 => AFLSDF_GND, 
        ADDRA9 => AFLSDF_GND, ADDRA8 => \GND\, ADDRA7 => 
        \U50_PATTERNS/ELINK_ADDRA_17[7]\, ADDRA6 => 
        \U50_PATTERNS/ELINK_ADDRA_17[6]\, ADDRA5 => 
        \U50_PATTERNS/ELINK_ADDRA_17[5]\, ADDRA4 => 
        \U50_PATTERNS/ELINK_ADDRA_17[4]\, ADDRA3 => 
        \U50_PATTERNS/ELINK_ADDRA_17[3]\, ADDRA2 => 
        \U50_PATTERNS/ELINK_ADDRA_17[2]\, ADDRA1 => 
        \U50_PATTERNS/ELINK_ADDRA_17[1]\, ADDRA0 => 
        \U50_PATTERNS/ELINK_ADDRA_17[0]\, ADDRB11 => AFLSDF_GND, 
        ADDRB10 => AFLSDF_GND, ADDRB9 => AFLSDF_GND, ADDRB8 => 
        \GND\, ADDRB7 => \ELKS_ADDRB[7]\, ADDRB6 => 
        \ELKS_ADDRB[6]\, ADDRB5 => \ELKS_ADDRB[5]\, ADDRB4 => 
        \ELKS_ADDRB[4]\, ADDRB3 => \ELKS_ADDRB[3]\, ADDRB2 => 
        \ELKS_ADDRB[2]\, ADDRB1 => \ELKS_ADDRB[1]\, ADDRB0 => 
        \ELKS_ADDRB[0]\, DINA8 => \GND\, DINA7 => 
        \U50_PATTERNS/ELINK_DINA_17[7]\, DINA6 => 
        \U50_PATTERNS/ELINK_DINA_17[6]\, DINA5 => 
        \U50_PATTERNS/ELINK_DINA_17[5]\, DINA4 => 
        \U50_PATTERNS/ELINK_DINA_17[4]\, DINA3 => 
        \U50_PATTERNS/ELINK_DINA_17[3]\, DINA2 => 
        \U50_PATTERNS/ELINK_DINA_17[2]\, DINA1 => 
        \U50_PATTERNS/ELINK_DINA_17[1]\, DINA0 => 
        \U50_PATTERNS/ELINK_DINA_17[0]\, DINB8 => \GND\, DINB7
         => \ELK_RX_SER_WORD_17[7]\, DINB6 => 
        \ELK_RX_SER_WORD_17[6]\, DINB5 => \ELK_RX_SER_WORD_17[5]\, 
        DINB4 => \ELK_RX_SER_WORD_17[4]\, DINB3 => 
        \ELK_RX_SER_WORD_17[3]\, DINB2 => \ELK_RX_SER_WORD_17[2]\, 
        DINB1 => \ELK_RX_SER_WORD_17[1]\, DINB0 => 
        \ELK_RX_SER_WORD_17[0]\, WIDTHA0 => \VCC\, WIDTHA1 => 
        \VCC\, WIDTHB0 => \VCC\, WIDTHB1 => \VCC\, PIPEA => \VCC\, 
        PIPEB => \VCC\, WMODEA => \GND\, WMODEB => \GND\, BLKA
         => \U50_PATTERNS/ELINK_BLKA[17]\, BLKB => 
        ELKS_RAM_BLKB_EN, WENA => \U50_PATTERNS/ELINK_RWA[17]\, 
        WENB => ELKS_RWB, CLKA => CLK60MHZ, CLKB => CLK_40M_GL, 
        RESET => P_USB_MASTER_EN_c_0, DOUTA8 => OPEN, DOUTA7 => 
        \U50_PATTERNS/ELINK_DOUTA_17[7]\, DOUTA6 => 
        \U50_PATTERNS/ELINK_DOUTA_17[6]\, DOUTA5 => 
        \U50_PATTERNS/ELINK_DOUTA_17[5]\, DOUTA4 => 
        \U50_PATTERNS/ELINK_DOUTA_17[4]\, DOUTA3 => 
        \U50_PATTERNS/ELINK_DOUTA_17[3]\, DOUTA2 => 
        \U50_PATTERNS/ELINK_DOUTA_17[2]\, DOUTA1 => 
        \U50_PATTERNS/ELINK_DOUTA_17[1]\, DOUTA0 => 
        \U50_PATTERNS/ELINK_DOUTA_17[0]\, DOUTB8 => OPEN, DOUTB7
         => \PATT_ELK_DAT_17[7]\, DOUTB6 => \PATT_ELK_DAT_17[6]\, 
        DOUTB5 => \PATT_ELK_DAT_17[5]\, DOUTB4 => 
        \PATT_ELK_DAT_17[4]\, DOUTB3 => \PATT_ELK_DAT_17[3]\, 
        DOUTB2 => \PATT_ELK_DAT_17[2]\, DOUTB1 => 
        \PATT_ELK_DAT_17[1]\, DOUTB0 => \PATT_ELK_DAT_17[0]\);
    
    \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[10]\ : DFN1C0
      port map(D => 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\);
    
    \U50_PATTERNS/ELINK_ADDRA_19[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120013, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_13, Q => 
        \U50_PATTERNS/ELINK_ADDRA_19[2]\);
    
    HIEFFPLA_INST_0_55754 : MX2
      port map(A => HIEFFPLA_NET_0_116973, B => 
        HIEFFPLA_NET_0_116960, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[4]\, Y => 
        HIEFFPLA_NET_0_116994);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_8[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_115969, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_19, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_8[1]\);
    
    HIEFFPLA_INST_0_40828 : MX2
      port map(A => HIEFFPLA_NET_0_119575, B => 
        \U50_PATTERNS/ELINK_DINA_17[2]\, S => 
        HIEFFPLA_NET_0_119260, Y => HIEFFPLA_NET_0_119805);
    
    HIEFFPLA_INST_0_47642 : MX2
      port map(A => HIEFFPLA_NET_0_118451, B => 
        HIEFFPLA_NET_0_118448, S => \BIT_OS_SEL_2[1]\, Y => 
        HIEFFPLA_NET_0_118453);
    
    \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[14]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_WRD_40M_FIXED[14]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_33, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[14]_net_1\);
    
    \U_ELK10_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL\ : DFN1C0
      port map(D => 
        \U_ELK10_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL_net_1\);
    
    HIEFFPLA_INST_0_46582 : AND2A
      port map(A => \OP_MODE_c_4[1]\, B => \PATT_ELK_DAT_0[6]\, Y
         => HIEFFPLA_NET_0_118654);
    
    AFLSDF_INV_12 : INV
      port map(A => DCB_SALT_SEL_c, Y => \AFLSDF_INV_12\);
    
    \U_ELK3_CH/U_SLAVE_1ELK/RECD_SER_WORD[6]\ : DFN1C0
      port map(D => \U_ELK3_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[6]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_3[6]\);
    
    HIEFFPLA_INST_0_41818 : AOI1B
      port map(A => HIEFFPLA_NET_0_119389, B => 
        \U50_PATTERNS/SM_BANK_SEL[9]\, C => HIEFFPLA_NET_0_119663, 
        Y => HIEFFPLA_NET_0_119690);
    
    \P_USB_TXE_B_pad/U0/U0\ : IOPAD_IN_U
      port map(PAD => P_USB_TXE_B, Y => \P_USB_TXE_B_pad/U0/NET1\);
    
    \U_ELK8_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]\ : DFN1C0
      port map(D => \U_ELK8_CH/U_SLAVE_1ELK/Q[10]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]_net_1\);
    
    \U50_PATTERNS/U0_PATT_TFC_BLK/DPRT_512X9_SRAM_R0C0\ : RAM4K9
      generic map(MEMORYFILE => "DPRT_512X9_SRAM_R0C0.mem")

      port map(ADDRA11 => AFLSDF_GND, ADDRA10 => AFLSDF_GND, 
        ADDRA9 => AFLSDF_GND, ADDRA8 => \GND\, ADDRA7 => 
        \U50_PATTERNS/TFC_ADDRA[7]\, ADDRA6 => 
        \U50_PATTERNS/TFC_ADDRA[6]\, ADDRA5 => 
        \U50_PATTERNS/TFC_ADDRA[5]\, ADDRA4 => 
        \U50_PATTERNS/TFC_ADDRA[4]\, ADDRA3 => 
        \U50_PATTERNS/TFC_ADDRA[3]\, ADDRA2 => 
        \U50_PATTERNS/TFC_ADDRA[2]\, ADDRA1 => 
        \U50_PATTERNS/TFC_ADDRA[1]\, ADDRA0 => 
        \U50_PATTERNS/TFC_ADDRA[0]\, ADDRB11 => AFLSDF_GND, 
        ADDRB10 => AFLSDF_GND, ADDRB9 => AFLSDF_GND, ADDRB8 => 
        \GND\, ADDRB7 => \TFC_ADDRB[7]\, ADDRB6 => \TFC_ADDRB[6]\, 
        ADDRB5 => \TFC_ADDRB[5]\, ADDRB4 => \TFC_ADDRB[4]\, 
        ADDRB3 => \TFC_ADDRB[3]\, ADDRB2 => \TFC_ADDRB[2]\, 
        ADDRB1 => \TFC_ADDRB[1]\, ADDRB0 => \TFC_ADDRB[0]\, DINA8
         => \GND\, DINA7 => \U50_PATTERNS/TFC_DINA[7]\, DINA6 => 
        \U50_PATTERNS/TFC_DINA[6]\, DINA5 => 
        \U50_PATTERNS/TFC_DINA[5]\, DINA4 => 
        \U50_PATTERNS/TFC_DINA[4]\, DINA3 => 
        \U50_PATTERNS/TFC_DINA[3]\, DINA2 => 
        \U50_PATTERNS/TFC_DINA[2]\, DINA1 => 
        \U50_PATTERNS/TFC_DINA[1]\, DINA0 => 
        \U50_PATTERNS/TFC_DINA[0]\, DINB8 => \GND\, DINB7 => 
        \TFC_RX_SER_WORD[7]\, DINB6 => \TFC_RX_SER_WORD[6]\, 
        DINB5 => \TFC_RX_SER_WORD[5]\, DINB4 => 
        \TFC_RX_SER_WORD[4]\, DINB3 => \TFC_RX_SER_WORD[3]\, 
        DINB2 => \TFC_RX_SER_WORD[2]\, DINB1 => 
        \TFC_RX_SER_WORD[1]\, DINB0 => \TFC_RX_SER_WORD[0]\, 
        WIDTHA0 => \VCC\, WIDTHA1 => \VCC\, WIDTHB0 => \VCC\, 
        WIDTHB1 => \VCC\, PIPEA => \VCC\, PIPEB => \VCC\, WMODEA
         => \GND\, WMODEB => \GND\, BLKA => 
        \U50_PATTERNS/TFC_BLKA\, BLKB => TFC_RAM_BLKB_EN, WENA
         => \U50_PATTERNS/TFC_RWA\, WENB => TFC_RWB, CLKA => 
        CLK60MHZ, CLKB => CLK_40M_GL, RESET => 
        P_USB_MASTER_EN_c_0, DOUTA8 => OPEN, DOUTA7 => 
        \U50_PATTERNS/TFC_DOUTA[7]\, DOUTA6 => 
        \U50_PATTERNS/TFC_DOUTA[6]\, DOUTA5 => 
        \U50_PATTERNS/TFC_DOUTA[5]\, DOUTA4 => 
        \U50_PATTERNS/TFC_DOUTA[4]\, DOUTA3 => 
        \U50_PATTERNS/TFC_DOUTA[3]\, DOUTA2 => 
        \U50_PATTERNS/TFC_DOUTA[2]\, DOUTA1 => 
        \U50_PATTERNS/TFC_DOUTA[1]\, DOUTA0 => 
        \U50_PATTERNS/TFC_DOUTA[0]\, DOUTB8 => OPEN, DOUTB7 => 
        \PATT_TFC_DAT[7]\, DOUTB6 => \PATT_TFC_DAT[6]\, DOUTB5
         => \PATT_TFC_DAT[5]\, DOUTB4 => \PATT_TFC_DAT[4]\, 
        DOUTB3 => \PATT_TFC_DAT[3]\, DOUTB2 => \PATT_TFC_DAT[2]\, 
        DOUTB1 => \PATT_TFC_DAT[1]\, DOUTB0 => \PATT_TFC_DAT[0]\);
    
    HIEFFPLA_INST_0_37522 : NAND3C
      port map(A => \U200A_TFC/RX_SER_WORD_3DEL_i_0[3]\, B => 
        \U200A_TFC/RX_SER_WORD_3DEL_i_0[2]\, C => 
        HIEFFPLA_NET_0_120267, Y => HIEFFPLA_NET_0_120268);
    
    \U_ELK18_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]\ : DFN1C0
      port map(D => \U_ELK18_CH/U_SLAVE_1ELK/Q[7]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]_net_1\);
    
    HIEFFPLA_INST_0_47202 : MX2
      port map(A => \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\, 
        B => \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[12]_net_1\, S => 
        \BIT_OS_SEL_4[2]\, Y => HIEFFPLA_NET_0_118535);
    
    HIEFFPLA_INST_0_43642 : NAND3C
      port map(A => HIEFFPLA_NET_0_119273, B => 
        \U50_PATTERNS/SM_BANK_SEL[5]\, C => 
        \U50_PATTERNS/SM_BANK_SEL[8]\, Y => HIEFFPLA_NET_0_119256);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_7[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_115977, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_17_0, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_7[3]\);
    
    \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[10]\ : DFN1C0
      port map(D => 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]_net_1\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\);
    
    \U_ELK16_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U3\ : IOBI_ID_OD_EB
      port map(DR => \U_ELK16_CH/ELK_OUT_R\, DF => 
        \U_ELK16_CH/ELK_OUT_F\, CLR => \GND\, E => 
        \AFLSDF_INV_27\, ICLK => CCC_160M_ADJ, OCLK => 
        CCC_160M_FXD, YIN => 
        \U_ELK16_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\, DOUT => 
        OPEN, EOUT => 
        \U_ELK16_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET3\, YR => OPEN, 
        YF => OPEN);
    
    \U50_PATTERNS/ELINK_DINA_2[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119775, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_9, Q => 
        \U50_PATTERNS/ELINK_DINA_2[0]\);
    
    HIEFFPLA_INST_0_52295 : AND3A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[4]_net_1\, B => 
        HIEFFPLA_NET_0_117598, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[5]_net_1\, Y => 
        HIEFFPLA_NET_0_117588);
    
    HIEFFPLA_INST_0_52236 : AND2A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[2]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[3]_net_1\, Y => 
        HIEFFPLA_NET_0_117603);
    
    \U_ELK10_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]\ : DFN1C0
      port map(D => \U_ELK10_CH/U_SLAVE_1ELK/Q[4]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]_net_1\);
    
    HIEFFPLA_INST_0_50611 : AND2A
      port map(A => \OP_MODE_c_4[1]\, B => \PATT_ELK_DAT_7[4]\, Y
         => HIEFFPLA_NET_0_117919);
    
    HIEFFPLA_INST_0_49764 : MX2
      port map(A => HIEFFPLA_NET_0_118086, B => 
        HIEFFPLA_NET_0_118082, S => \BIT_OS_SEL_1[0]\, Y => 
        \U_ELK3_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[4]\);
    
    HIEFFPLA_INST_0_43119 : AND3B
      port map(A => \U50_PATTERNS/REG_STATE[1]_net_1\, B => 
        \U50_PATTERNS/REG_STATE[3]_net_1\, C => 
        \U50_PATTERNS/REG_STATE[0]_net_1\, Y => 
        HIEFFPLA_NET_0_119369);
    
    \U_ELK2_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118152, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_8, Q => 
        \U_ELK2_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]_net_1\);
    
    HIEFFPLA_INST_0_46625 : NAND2B
      port map(A => \OP_MODE_c_3[1]\, B => \PATT_ELK_DAT_10[2]\, 
        Y => HIEFFPLA_NET_0_118641);
    
    HIEFFPLA_INST_0_45316 : AO1A
      port map(A => HIEFFPLA_NET_0_118824, B => 
        \U50_PATTERNS/SM_BANK_SEL[15]\, C => 
        HIEFFPLA_NET_0_118816, Y => HIEFFPLA_NET_0_118943);
    
    HIEFFPLA_INST_0_55354 : AND3A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[5]_net_1\, B => 
        HIEFFPLA_NET_0_115906, C => 
        \U_MASTER_DES/CCC_RX_CLK_LOCK\, Y => 
        HIEFFPLA_NET_0_117053);
    
    \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[2]\ : DFN1C0
      port map(D => 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[2]_net_1\);
    
    \U_ELK0_SERDAT_SOURCE/SERDAT[4]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118656, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_10, Q => \ELK0_TX_DAT[4]\);
    
    HIEFFPLA_INST_0_59700 : MX2
      port map(A => HIEFFPLA_NET_0_116687, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_2[2]\, S => 
        HIEFFPLA_NET_0_117206, Y => HIEFFPLA_NET_0_116359);
    
    HIEFFPLA_INST_0_53287 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_SEQCNT[3]\, B => 
        HIEFFPLA_NET_0_117434, S => HIEFFPLA_NET_0_117062, Y => 
        HIEFFPLA_NET_0_117439);
    
    HIEFFPLA_INST_0_44973 : AND3C
      port map(A => HIEFFPLA_NET_0_119635, B => 
        HIEFFPLA_NET_0_119399, C => HIEFFPLA_NET_0_119005, Y => 
        HIEFFPLA_NET_0_119008);
    
    HIEFFPLA_INST_0_38274 : MX2
      port map(A => \U50_PATTERNS/ELINKS_STOP_ADDR[4]\, B => 
        \U50_PATTERNS/ELINKS_STOP_ADDR_T[4]\, S => 
        HIEFFPLA_NET_0_119472, Y => HIEFFPLA_NET_0_120123);
    
    HIEFFPLA_INST_0_46800 : MX2
      port map(A => HIEFFPLA_NET_0_118627, B => 
        HIEFFPLA_NET_0_118610, S => \BIT_OS_SEL_0[0]\, Y => 
        \U_ELK10_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[7]\);
    
    HIEFFPLA_INST_0_44330 : XOR2
      port map(A => \TFC_STRT_ADDR[2]\, B => 
        \U50_PATTERNS/U4A_REGCROSS/SAMP_TWO[2]_net_1\, Y => 
        HIEFFPLA_NET_0_119139);
    
    \U_ELK2_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]\ : DFN1C0
      port map(D => \U_ELK2_CH/U_SLAVE_1ELK/Q[0]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]_net_1\);
    
    \U_ELK0_SERDAT_SOURCE/SERDAT[5]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118655, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_10, Q => \ELK0_TX_DAT[5]\);
    
    \U50_PATTERNS/ELINK_DINA_3[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119762, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_11, Q => 
        \U50_PATTERNS/ELINK_DINA_3[5]\);
    
    HIEFFPLA_INST_0_46304 : NAND3C
      port map(A => HIEFFPLA_NET_0_119620, B => 
        HIEFFPLA_NET_0_119625, C => HIEFFPLA_NET_0_118886, Y => 
        HIEFFPLA_NET_0_118721);
    
    \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[8]\ : DFN1C0
      port map(D => \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\);
    
    HIEFFPLA_INST_0_48377 : MX2
      port map(A => HIEFFPLA_NET_0_118317, B => 
        HIEFFPLA_NET_0_118314, S => \BIT_OS_SEL_1[1]\, Y => 
        HIEFFPLA_NET_0_118320);
    
    HIEFFPLA_INST_0_49363 : NAND2B
      port map(A => \OP_MODE_c_1[1]\, B => \PATT_ELK_DAT_2[1]\, Y
         => HIEFFPLA_NET_0_118147);
    
    HIEFFPLA_INST_0_57278 : NAND3B
      port map(A => HIEFFPLA_NET_0_116715, B => 
        HIEFFPLA_NET_0_116710, C => HIEFFPLA_NET_0_116713, Y => 
        HIEFFPLA_NET_0_116708);
    
    HIEFFPLA_INST_0_53965 : MX2
      port map(A => HIEFFPLA_NET_0_116318, B => 
        HIEFFPLA_NET_0_116374, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[3]_net_1\, Y
         => HIEFFPLA_NET_0_117326);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_14[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116525, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_13, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_14[3]\);
    
    \P_CCC_160M_ADJ_pad/U0/U1\ : IOTRI_OB_EB
      port map(D => CCC_160M_ADJ, E => \VCC\, DOUT => 
        \P_CCC_160M_ADJ_pad/U0/NET1\, EOUT => 
        \P_CCC_160M_ADJ_pad/U0/NET2\);
    
    HIEFFPLA_INST_0_54994 : NAND2B
      port map(A => HIEFFPLA_NET_0_117182, B => 
        HIEFFPLA_NET_0_117145, Y => HIEFFPLA_NET_0_117146);
    
    HIEFFPLA_INST_0_54031 : MX2
      port map(A => HIEFFPLA_NET_0_116200, B => 
        HIEFFPLA_NET_0_116084, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[3]_net_1\, Y
         => HIEFFPLA_NET_0_117317);
    
    \U_EXEC_MASTER/PRESCALE[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117768, CLK => CLK_40M_GL, CLR
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i\, Q => 
        \U_EXEC_MASTER/PRESCALE[0]\);
    
    HIEFFPLA_INST_0_42311 : AND2A
      port map(A => HIEFFPLA_NET_0_119275, B => 
        \U50_PATTERNS/RD_USB_ADBUS[2]\, Y => 
        HIEFFPLA_NET_0_119575);
    
    \U_ELK5_CH/U_SLAVE_1ELK/RECD_SER_WORD[2]\ : DFN1C0
      port map(D => \U_ELK5_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[2]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_5[2]\);
    
    HIEFFPLA_INST_0_58157 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_10[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_26[1]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_2[4]_net_1\, Y
         => HIEFFPLA_NET_0_116557);
    
    HIEFFPLA_INST_0_55452 : MX2
      port map(A => HIEFFPLA_NET_0_116974, B => 
        HIEFFPLA_NET_0_117030, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[2]\, Y => 
        HIEFFPLA_NET_0_117035);
    
    \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_1S\ : DFN1C0
      port map(D => 
        \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_S_net_1\, CLK => 
        CLK60MHZ, CLR => P_MASTER_POR_B_c_22_0, Q => 
        \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_1S_net_1\);
    
    \U50_PATTERNS/ELINK_ADDRA_2[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119999, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_21, Q => 
        \U50_PATTERNS/ELINK_ADDRA_2[0]\);
    
    HIEFFPLA_INST_0_57047 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_2[4]\, B => 
        HIEFFPLA_NET_0_116731, S => HIEFFPLA_NET_0_117601, Y => 
        HIEFFPLA_NET_0_116751);
    
    HIEFFPLA_INST_0_41723 : MX2
      port map(A => HIEFFPLA_NET_0_119684, B => 
        \U50_PATTERNS/ELINK_RWA[16]\, S => 
        \U50_PATTERNS/SM_BANK_SEL_0[20]\, Y => 
        HIEFFPLA_NET_0_119704);
    
    \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[6]\ : DFN1C0
      port map(D => \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\);
    
    HIEFFPLA_INST_0_41629 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_9[3]\, B => 
        HIEFFPLA_NET_0_119574, S => HIEFFPLA_NET_0_119292, Y => 
        HIEFFPLA_NET_0_119716);
    
    HIEFFPLA_INST_0_57863 : NAND2A
      port map(A => HIEFFPLA_NET_0_116618, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_6[7]\, Y => 
        HIEFFPLA_NET_0_116604);
    
    HIEFFPLA_INST_0_50728 : MX2
      port map(A => HIEFFPLA_NET_0_117891, B => 
        HIEFFPLA_NET_0_117900, S => \BIT_OS_SEL_5[0]\, Y => 
        \U_ELK7_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[0]\);
    
    HIEFFPLA_INST_0_42620 : AOI1A
      port map(A => HIEFFPLA_NET_0_119521, B => 
        \U50_PATTERNS/REG_ADDR[5]\, C => 
        \U50_PATTERNS/REG_ADDR[6]\, Y => HIEFFPLA_NET_0_119498);
    
    \U50_PATTERNS/TFC_STOP_ADDR_T[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119180, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_15, Q => 
        \U50_PATTERNS/TFC_STOP_ADDR_T[0]\);
    
    HIEFFPLA_INST_0_50744 : MX2
      port map(A => HIEFFPLA_NET_0_117914, B => 
        HIEFFPLA_NET_0_117911, S => \BIT_OS_SEL_5[0]\, Y => 
        \U_ELK7_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[2]\);
    
    TFC_IN_R : DFN1C0
      port map(D => TFC_IN_DDR_R, CLK => CCC_160M_ADJ, CLR => 
        DEV_RST_B_c, Q => \TFC_IN_R\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[10]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_WRD_40M_FIXED[10]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_32_0, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[10]_net_1\);
    
    HIEFFPLA_INST_0_57259 : NAND2B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_3[7]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_3[6]\, Y => 
        HIEFFPLA_NET_0_116715);
    
    HIEFFPLA_INST_0_51718 : NAND2B
      port map(A => 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM[4]_net_1\, B => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[71]_net_1\, Y => 
        HIEFFPLA_NET_0_117708);
    
    HIEFFPLA_INST_0_56143 : NAND3A
      port map(A => HIEFFPLA_NET_0_116940, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/MAX_CNT[6]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/MAX_CNT[5]\, Y => 
        HIEFFPLA_NET_0_116945);
    
    \U_ELK3_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118111, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_16, Q => 
        \U_ELK3_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]_net_1\);
    
    HIEFFPLA_INST_0_63217 : AND2
      port map(A => \TFC_TX_DAT[1]\, B => 
        \U_TFC_CMD_TX/START_RISE_net_1\, Y => 
        \U_TFC_CMD_TX/N_SER_CMD_WORD_R[0]\);
    
    HIEFFPLA_INST_0_54229 : MX2
      port map(A => HIEFFPLA_NET_0_116567, B => 
        HIEFFPLA_NET_0_116289, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_1[3]_net_1\, Y
         => HIEFFPLA_NET_0_117292);
    
    \U50_PATTERNS/ELINK_ADDRA_16[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120039, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_8, Q => 
        \U50_PATTERNS/ELINK_ADDRA_16[0]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/TUNE_CLKPHASE[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_115946, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_13, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/TUNE_CLKPHASE[3]\);
    
    HIEFFPLA_INST_0_63057 : AND2B
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[8]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[12]\, Y => 
        HIEFFPLA_NET_0_115899);
    
    HIEFFPLA_INST_0_61916 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_27[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_28[1]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[0]\, Y => 
        HIEFFPLA_NET_0_116060);
    
    HIEFFPLA_INST_0_49009 : MX2
      port map(A => HIEFFPLA_NET_0_118227, B => 
        HIEFFPLA_NET_0_118223, S => \BIT_OS_SEL_2[0]\, Y => 
        \U_ELK19_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[3]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_SEL_2[1]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_BIT_OS_VAL[1]\, CLK
         => CLK_40M_GL, CLR => P_MASTER_POR_B_c_27_0, Q => 
        \BIT_OS_SEL_2[1]\);
    
    \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[2]\ : DFN1C0
      port map(D => \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\);
    
    HIEFFPLA_INST_0_47989 : MX2
      port map(A => HIEFFPLA_NET_0_118386, B => 
        HIEFFPLA_NET_0_118402, S => \BIT_OS_SEL_3[0]\, Y => 
        \U_ELK15_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[0]\);
    
    \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[11]\ : DFN1C0
      port map(D => 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[11]_net_1\);
    
    \U_ELK11_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2\ : IOPADN_BI
      port map(DB => \U_ELK11_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, 
        E => \U_ELK11_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET3\, PAD
         => ELK11_DAT_N, N2POUT => 
        \U_ELK11_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2_N2P\);
    
    HIEFFPLA_INST_0_53647 : AND2A
      port map(A => HIEFFPLA_NET_0_117377, B => 
        HIEFFPLA_NET_0_117334, Y => HIEFFPLA_NET_0_117378);
    
    HIEFFPLA_INST_0_40198 : AOI1D
      port map(A => HIEFFPLA_NET_0_119389, B => 
        HIEFFPLA_NET_0_119464, C => \U50_PATTERNS/SM_BANK_SEL[1]\, 
        Y => HIEFFPLA_NET_0_119875);
    
    \U_ELK6_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]\ : DFN1C0
      port map(D => \U_ELK6_CH/U_SLAVE_1ELK/Q[5]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]_net_1\);
    
    HIEFFPLA_INST_0_44214 : MX2
      port map(A => \U50_PATTERNS/TFC_STRT_ADDR_T[5]\, B => 
        \U50_PATTERNS/RD_USB_ADBUS[5]\, S => 
        HIEFFPLA_NET_0_119491, Y => HIEFFPLA_NET_0_119159);
    
    HIEFFPLA_INST_0_60816 : MX2
      port map(A => HIEFFPLA_NET_0_117190, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_16[0]\, S => 
        HIEFFPLA_NET_0_117142, Y => HIEFFPLA_NET_0_116215);
    
    HIEFFPLA_INST_0_55659 : MX2
      port map(A => HIEFFPLA_NET_0_115986, B => 
        HIEFFPLA_NET_0_116237, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_2[3]\, Y => 
        HIEFFPLA_NET_0_117007);
    
    HIEFFPLA_INST_0_47429 : MX2
      port map(A => \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\, 
        B => \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\, S => 
        \BIT_OS_SEL_3[2]\, Y => HIEFFPLA_NET_0_118493);
    
    HIEFFPLA_INST_0_42165 : MX2
      port map(A => \U50_PATTERNS/OP_MODE_T[1]\, B => 
        \U50_PATTERNS/RD_USB_ADBUS[1]\, S => 
        HIEFFPLA_NET_0_119440, Y => HIEFFPLA_NET_0_119608);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_16[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116215, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_5, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_16[0]\);
    
    \U50_PATTERNS/SM_BANK_SEL[17]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119314, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_1_0, Q => 
        \U50_PATTERNS/SM_BANK_SEL[17]\);
    
    HIEFFPLA_INST_0_60859 : AND2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[4]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_16[1]\, Y => 
        HIEFFPLA_NET_0_116209);
    
    HIEFFPLA_INST_0_49547 : MX2
      port map(A => HIEFFPLA_NET_0_118114, B => 
        HIEFFPLA_NET_0_118138, S => \BIT_OS_SEL[1]\, Y => 
        HIEFFPLA_NET_0_118116);
    
    HIEFFPLA_INST_0_41539 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_8[1]\, B => 
        HIEFFPLA_NET_0_119576, S => HIEFFPLA_NET_0_119291, Y => 
        HIEFFPLA_NET_0_119726);
    
    \U_ELK9_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U1\ : IOBI_ID_OD_EB
      port map(DR => \U_ELK9_CH/ELK_OUT_R\, DF => 
        \U_ELK9_CH/ELK_OUT_F\, CLR => \GND\, E => \AFLSDF_INV_50\, 
        ICLK => CCC_160M_ADJ, OCLK => CCC_160M_FXD, YIN => 
        \U_ELK9_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\, DOUT => 
        \U_ELK9_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, EOUT => 
        \U_ELK9_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET2\, YR => 
        \U_ELK9_CH/ELK_IN_DDR_R\, YF => \U_ELK9_CH/ELK_IN_DDR_F\);
    
    \U_ELK15_CH/U_SLAVE_1ELK/Q[12]\ : DFN1C0
      port map(D => \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/Q[12]_net_1\);
    
    HIEFFPLA_INST_0_59600 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_13[3]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_29[3]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[4]_net_1\, Y => 
        HIEFFPLA_NET_0_116372);
    
    \U50_PATTERNS/RD_XFER_TYPE[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119546, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c, Q => 
        \U50_PATTERNS/RD_XFER_TYPE[3]_net_1\);
    
    \U_ELK6_CH/U_SLAVE_1ELK/Q[0]\ : DFN1C0
      port map(D => \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/Q[0]_net_1\);
    
    \U50_PATTERNS/ELINK_DINA_4[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119755, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_13, Q => 
        \U50_PATTERNS/ELINK_DINA_4[4]\);
    
    HIEFFPLA_INST_0_47282 : MX2
      port map(A => HIEFFPLA_NET_0_118542, B => 
        HIEFFPLA_NET_0_118536, S => \BIT_OS_SEL_5[0]\, Y => 
        \U_ELK12_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[5]\);
    
    \U50_PATTERNS/SM_BANK_SEL[18]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119313, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_1_0, Q => 
        \U50_PATTERNS/SM_BANK_SEL[18]\);
    
    HIEFFPLA_INST_0_37710 : AND3B
      port map(A => \U200B_ELINKS/GP_PG_SM[0]_net_1\, B => 
        \U200B_ELINKS/GP_PG_SM[1]_net_1\, C => 
        HIEFFPLA_NET_0_120226, Y => HIEFFPLA_NET_0_120223);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_17[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116498, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_18, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_17[3]\);
    
    HIEFFPLA_INST_0_55342 : NAND3C
      port map(A => HIEFFPLA_NET_0_117047, B => 
        HIEFFPLA_NET_0_117050, C => HIEFFPLA_NET_0_117052, Y => 
        HIEFFPLA_NET_0_117055);
    
    \U50_PATTERNS/ELINKS_STOP_ADDR_T[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120117, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_7, Q => 
        \U50_PATTERNS/ELINKS_STOP_ADDR_T[2]\);
    
    HIEFFPLA_INST_0_58449 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_15[0]\, B => 
        HIEFFPLA_NET_0_116680, S => HIEFFPLA_NET_0_117098, Y => 
        HIEFFPLA_NET_0_116520);
    
    HIEFFPLA_INST_0_55989 : MX2
      port map(A => HIEFFPLA_NET_0_116961, B => 
        HIEFFPLA_NET_0_116992, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[4]\, Y => 
        HIEFFPLA_NET_0_116964);
    
    HIEFFPLA_INST_0_44642 : XOR2
      port map(A => \ELKS_STOP_ADDR[1]\, B => 
        \U50_PATTERNS/U4D_REGCROSS/SAMP_TWO[1]_net_1\, Y => 
        HIEFFPLA_NET_0_119076);
    
    \U50_PATTERNS/U4A_REGCROSS/SAMP_TWO[3]\ : DFN1C0
      port map(D => \U50_PATTERNS/U4A_REGCROSS/SAMP_ONE[3]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_22, Q => 
        \U50_PATTERNS/U4A_REGCROSS/SAMP_TWO[3]_net_1\);
    
    HIEFFPLA_INST_0_54932 : XO1A
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[3]\, 
        B => HIEFFPLA_NET_0_115870, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_0[8]_net_1\, Y => 
        HIEFFPLA_NET_0_117168);
    
    HIEFFPLA_INST_0_57001 : AOI1A
      port map(A => HIEFFPLA_NET_0_116777, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_1[6]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_1[7]\, Y => 
        HIEFFPLA_NET_0_116756);
    
    HIEFFPLA_INST_0_42908 : NAND3A
      port map(A => HIEFFPLA_NET_0_119430, B => 
        HIEFFPLA_NET_0_119378, C => HIEFFPLA_NET_0_119431, Y => 
        HIEFFPLA_NET_0_119427);
    
    \U50_PATTERNS/ELINK_DINA_11[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119852, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_11, Q => 
        \U50_PATTERNS/ELINK_DINA_11[3]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_4[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116693, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_9, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_4[3]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_3[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116724, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_7, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_3[1]\);
    
    \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[8]\ : DFN1C0
      port map(D => 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\);
    
    \U200B_ELINKS/RX_SER_WORD_3DEL[6]\ : DFN1C0
      port map(D => \U200B_ELINKS/RX_SER_WORD_2DEL[6]_net_1\, CLK
         => CLK_40M_GL, CLR => P_MASTER_POR_B_c_31_0, Q => 
        \U200B_ELINKS/RX_SER_WORD_3DEL[6]_net_1\);
    
    HIEFFPLA_INST_0_56443 : AND3
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[9]_net_1\, B => 
        HIEFFPLA_NET_0_117427, C => HIEFFPLA_NET_0_117423, Y => 
        HIEFFPLA_NET_0_116866);
    
    HIEFFPLA_INST_0_57174 : AXOI4
      port map(A => HIEFFPLA_NET_0_117085, B => 
        HIEFFPLA_NET_0_117120, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_3[0]\, Y => 
        HIEFFPLA_NET_0_116725);
    
    \U_ELK15_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118427, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_9, Q => 
        \U_ELK15_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_0[4]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116820, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_3, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_0[4]\);
    
    HIEFFPLA_INST_0_59159 : AND3A
      port map(A => HIEFFPLA_NET_0_116424, B => 
        HIEFFPLA_NET_0_116422, C => HIEFFPLA_NET_0_117249, Y => 
        HIEFFPLA_NET_0_116427);
    
    HIEFFPLA_INST_0_57712 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_6[1]\, B => 
        HIEFFPLA_NET_0_116615, S => HIEFFPLA_NET_0_117599, Y => 
        HIEFFPLA_NET_0_116631);
    
    HIEFFPLA_INST_0_111825 : AX1E
      port map(A => 
        \U_EXEC_MASTER/USB_MASTER_EN/T_CNT60M[1]_net_1\, B => 
        \U_EXEC_MASTER/USB_MASTER_EN/T_CNT60M[0]_net_1\, C => 
        \U_EXEC_MASTER/USB_MASTER_EN/T_CNT60M[2]_net_1\, Y => 
        HIEFFPLA_NET_0_115827);
    
    \U_MASTER_DES/U13C_MASTER_DESER/ARB_WRD_40M_FIXED[13]\ : 
        DFN1C0
      port map(D => \U_MASTER_DES/U13C_MASTER_DESER/Q[13]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_28, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_WRD_40M_FIXED[13]_net_1\);
    
    HIEFFPLA_INST_0_39506 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_4[0]\, B => 
        HIEFFPLA_NET_0_119524, S => HIEFFPLA_NET_0_119284, Y => 
        HIEFFPLA_NET_0_119983);
    
    HIEFFPLA_INST_0_45378 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_14[4]\, C => 
        \U50_PATTERNS/SM_BANK_SEL[5]\, Y => HIEFFPLA_NET_0_118926);
    
    \U_ELK7_CH/U_ELK1_SERDAT_SOURCE/SERDAT[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117922, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_3, Q => 
        \U_ELK7_CH/ELK_TX_DAT[1]\);
    
    \U_ELK17_CH/U_SLAVE_1ELK/RECD_SER_WORD[7]\ : DFN1C0
      port map(D => \U_ELK17_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[7]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_17[7]\);
    
    \U50_PATTERNS/U4E_REGCROSS/SAMP_ONE[3]\ : DFN1C0
      port map(D => \U50_PATTERNS/OP_MODE[3]\, CLK => CLK_40M_GL, 
        CLR => P_MASTER_POR_B_c, Q => 
        \U50_PATTERNS/U4E_REGCROSS/SAMP_ONE[3]_net_1\);
    
    \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[6]\ : DFN1C0
      port map(D => \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\);
    
    HIEFFPLA_INST_0_52958 : MX2
      port map(A => HIEFFPLA_NET_0_117471, B => 
        HIEFFPLA_NET_0_117467, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[4]\, Y => 
        HIEFFPLA_NET_0_117483);
    
    \U50_PATTERNS/ELINK_ADDRA_19[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120015, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_13, Q => 
        \U50_PATTERNS/ELINK_ADDRA_19[0]\);
    
    HIEFFPLA_INST_0_37453 : MX2
      port map(A => \U200A_TFC/LOC_STRT_ADDR[0]\, B => 
        \TFC_STRT_ADDR[0]\, S => \U200A_TFC/GP_PG_SM_0[10]_net_1\, 
        Y => HIEFFPLA_NET_0_120282);
    
    \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[8]\ : DFN1C0
      port map(D => 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\);
    
    HIEFFPLA_INST_0_50112 : NAND2B
      port map(A => \OP_MODE_c_4[1]\, B => \PATT_ELK_DAT_5[3]\, Y
         => HIEFFPLA_NET_0_118010);
    
    \U_ELK19_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]\ : DFN1C0
      port map(D => \U_ELK19_CH/U_SLAVE_1ELK/Q[6]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]_net_1\);
    
    \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[9]\ : DFN1C0
      port map(D => 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\);
    
    HIEFFPLA_INST_0_56216 : AND3A
      port map(A => \ELK_RX_SER_WORD_0[6]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/RECD_SER_WORD[3]_net_1\, 
        C => \ELK_RX_SER_WORD_0[7]\, Y => HIEFFPLA_NET_0_116928);
    
    HIEFFPLA_INST_0_54726 : NAND3B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[1]_net_1\, B => 
        HIEFFPLA_NET_0_117245, C => HIEFFPLA_NET_0_117251, Y => 
        HIEFFPLA_NET_0_117216);
    
    HIEFFPLA_INST_0_56465 : AOI1D
      port map(A => HIEFFPLA_NET_0_117432, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_SEL[3]_net_1\, C
         => \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[6]_net_1\, Y
         => HIEFFPLA_NET_0_116858);
    
    HIEFFPLA_INST_0_56621 : AND3
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[13]_net_1\, B
         => HIEFFPLA_NET_0_117424, C => HIEFFPLA_NET_0_117427, Y
         => HIEFFPLA_NET_0_116826);
    
    HIEFFPLA_INST_0_48230 : MX2
      port map(A => HIEFFPLA_NET_0_118363, B => 
        HIEFFPLA_NET_0_118360, S => \BIT_OS_SEL_1[1]\, Y => 
        HIEFFPLA_NET_0_118350);
    
    HIEFFPLA_INST_0_38543 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_0[5]\, B => 
        HIEFFPLA_NET_0_119518, S => HIEFFPLA_NET_0_119272, Y => 
        HIEFFPLA_NET_0_120090);
    
    HIEFFPLA_INST_0_48708 : MX2
      port map(A => \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\, 
        B => \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[12]_net_1\, S => 
        \BIT_OS_SEL_0[2]\, Y => HIEFFPLA_NET_0_118263);
    
    \U_ELK9_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]\ : DFN1C0
      port map(D => \U_ELK9_CH/U_SLAVE_1ELK/Q[7]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]_net_1\);
    
    HIEFFPLA_INST_0_50495 : MX2
      port map(A => HIEFFPLA_NET_0_117959, B => 
        HIEFFPLA_NET_0_117956, S => \BIT_OS_SEL[0]\, Y => 
        \U_ELK6_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[2]\);
    
    HIEFFPLA_INST_0_49572 : AND2
      port map(A => \U_ELK3_CH/ELK_TX_DAT[0]\, B => 
        \U_ELK3_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118112);
    
    AFLSDF_INV_35 : INV
      port map(A => DCB_SALT_SEL_c, Y => \AFLSDF_INV_35\);
    
    HIEFFPLA_INST_0_47079 : MX2
      port map(A => \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\, 
        B => \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[14]_net_1\, S => 
        \BIT_OS_SEL_7[2]\, Y => HIEFFPLA_NET_0_118563);
    
    HIEFFPLA_INST_0_41899 : AND2
      port map(A => HIEFFPLA_NET_0_119389, B => 
        \U50_PATTERNS/SM_BANK_SEL[12]\, Y => 
        HIEFFPLA_NET_0_119669);
    
    HIEFFPLA_INST_0_55204 : AND2A
      port map(A => HIEFFPLA_NET_0_117205, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[6]_net_1\, Y => 
        HIEFFPLA_NET_0_117092);
    
    HIEFFPLA_INST_0_38804 : MX2
      port map(A => HIEFFPLA_NET_0_119522, B => 
        \U50_PATTERNS/ELINK_ADDRA_13[2]\, S => 
        HIEFFPLA_NET_0_119285, Y => HIEFFPLA_NET_0_120061);
    
    HIEFFPLA_INST_0_54341 : MX2
      port map(A => HIEFFPLA_NET_0_116515, B => 
        HIEFFPLA_NET_0_116298, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_2[3]_net_1\, Y
         => HIEFFPLA_NET_0_117278);
    
    HIEFFPLA_INST_0_53903 : AND3A
      port map(A => HIEFFPLA_NET_0_117238, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[0]_net_1\, C
         => \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_1[3]_net_1\, 
        Y => HIEFFPLA_NET_0_117336);
    
    HIEFFPLA_INST_0_43255 : AND3B
      port map(A => HIEFFPLA_NET_0_119581, B => 
        HIEFFPLA_NET_0_119450, C => HIEFFPLA_NET_0_119600, Y => 
        HIEFFPLA_NET_0_119336);
    
    HIEFFPLA_INST_0_40666 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_15[0]\, B => 
        HIEFFPLA_NET_0_119578, S => HIEFFPLA_NET_0_119297, Y => 
        HIEFFPLA_NET_0_119823);
    
    HIEFFPLA_INST_0_40360 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_10[6]\, B => 
        HIEFFPLA_NET_0_119566, S => HIEFFPLA_NET_0_119239, Y => 
        HIEFFPLA_NET_0_119857);
    
    \U_EXEC_MASTER/MPOR_B_24_0\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117787, CLK => CLK_40M_GL, CLR
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_0\, Q => 
        P_MASTER_POR_B_c_24_0);
    
    \U50_PATTERNS/OP_MODE[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119615, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_15, Q => \U50_PATTERNS/OP_MODE[2]\);
    
    HIEFFPLA_INST_0_50836 : AND2
      port map(A => \U_ELK8_CH/ELK_TX_DAT[1]\, B => 
        \U_ELK8_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_117883);
    
    HIEFFPLA_INST_0_56404 : NAND3C
      port map(A => HIEFFPLA_NET_0_116827, B => 
        HIEFFPLA_NET_0_116843, C => HIEFFPLA_NET_0_116851, Y => 
        HIEFFPLA_NET_0_116875);
    
    \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[8]\ : DFN1C0
      port map(D => \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\);
    
    HIEFFPLA_INST_0_54047 : MX2
      port map(A => HIEFFPLA_NET_0_117248, B => 
        HIEFFPLA_NET_0_117313, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[2]_net_1\, Y
         => HIEFFPLA_NET_0_117315);
    
    HIEFFPLA_INST_0_51936 : AND3A
      port map(A => \U_MASTER_DES/U13A_ADJ_160M/BITCNT[0]\, B => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[34]_net_1\, C => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[1]\, Y => 
        HIEFFPLA_NET_0_117662);
    
    HIEFFPLA_INST_0_45307 : AO1A
      port map(A => HIEFFPLA_NET_0_118834, B => 
        \U50_PATTERNS/SM_BANK_SEL[7]\, C => HIEFFPLA_NET_0_118945, 
        Y => HIEFFPLA_NET_0_118946);
    
    HIEFFPLA_INST_0_62264 : AND2A
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[0]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_31[1]\, Y
         => HIEFFPLA_NET_0_116014);
    
    HIEFFPLA_INST_0_54935 : AND2A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_0[8]_net_1\, B => 
        HIEFFPLA_NET_0_115868, Y => HIEFFPLA_NET_0_117166);
    
    HIEFFPLA_INST_0_39137 : MX2
      port map(A => HIEFFPLA_NET_0_119516, B => 
        \U50_PATTERNS/ELINK_ADDRA_17[7]\, S => 
        HIEFFPLA_NET_0_119260, Y => HIEFFPLA_NET_0_120024);
    
    \U_ELK8_CH/U_SLAVE_1ELK/RECD_SER_WORD[3]\ : DFN1C0
      port map(D => \U_ELK8_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[3]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_8[3]\);
    
    \U50_PATTERNS/ELINKS_STOP_ADDR[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120122, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_14, Q => 
        \U50_PATTERNS/ELINKS_STOP_ADDR[5]\);
    
    HIEFFPLA_INST_0_62529 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_7[2]\, 
        B => HIEFFPLA_NET_0_117131, S => HIEFFPLA_NET_0_117174, Y
         => HIEFFPLA_NET_0_115978);
    
    \U_ELK19_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118247, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_7, Q => 
        \U_ELK19_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]_net_1\);
    
    \U0B_TX40M_REFCLK/_OUTBUF_LVDS[0]_/U0/U3\ : IOTRI_OB_EB
      port map(D => CLK_40M_BUF_RECD, E => \VCC\, DOUT => OPEN, 
        EOUT => OPEN);
    
    HIEFFPLA_INST_0_53522 : NAND3
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[4]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[2]_net_1\, C => 
        HIEFFPLA_NET_0_117318, Y => HIEFFPLA_NET_0_117395);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_27[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116392, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_2, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_27[2]\);
    
    \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[0]\ : DFN1C0
      port map(D => 
        \U_ELK11_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\);
    
    HIEFFPLA_INST_0_45274 : AO1
      port map(A => HIEFFPLA_NET_0_119263, B => 
        \U50_PATTERNS/ELINK_DOUTA_8[5]\, C => 
        HIEFFPLA_NET_0_118840, Y => HIEFFPLA_NET_0_118953);
    
    \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117042, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_17, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[3]\);
    
    \U_ELK16_CH/U_ELK1_CMD_TX/SER_OUT_RDEL\ : DFN1C0
      port map(D => \U_ELK16_CH/U_ELK1_CMD_TX/SER_OUT_RI_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_16, Q
         => \U_ELK16_CH/ELK_OUT_R\);
    
    HIEFFPLA_INST_0_61835 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_10[4]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_26[4]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_4[4]_net_1\, Y
         => HIEFFPLA_NET_0_116071);
    
    HIEFFPLA_INST_0_43739 : AND3A
      port map(A => \U50_PATTERNS/RD_USB_ADBUS[2]\, B => 
        HIEFFPLA_NET_0_119594, C => 
        \U50_PATTERNS/RD_USB_ADBUS[3]\, Y => 
        HIEFFPLA_NET_0_119226);
    
    HIEFFPLA_INST_0_50061 : MX2
      port map(A => \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[0]_net_1\, B
         => \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\, S => 
        \BIT_OS_SEL_6[2]\, Y => HIEFFPLA_NET_0_118024);
    
    HIEFFPLA_INST_0_46283 : NAND3C
      port map(A => HIEFFPLA_NET_0_118871, B => 
        HIEFFPLA_NET_0_118889, C => HIEFFPLA_NET_0_118897, Y => 
        HIEFFPLA_NET_0_118725);
    
    HIEFFPLA_INST_0_50089 : AND2
      port map(A => \U_ELK5_CH/ELK_TX_DAT[1]\, B => 
        \U_ELK5_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118018);
    
    \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[4]\ : DFN1C0
      port map(D => 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\);
    
    HIEFFPLA_INST_0_51674 : XOR2
      port map(A => \U_GEN_REF_CLK/GEN_40M_REFCNT[1]_net_1\, B
         => \U_GEN_REF_CLK/GEN_40M_REFCNT[0]_net_1\, Y => 
        HIEFFPLA_NET_0_117727);
    
    HIEFFPLA_INST_0_53765 : AO1A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_0[6]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_0[8]_net_1\, C => 
        HIEFFPLA_NET_0_117355, Y => HIEFFPLA_NET_0_117356);
    
    HIEFFPLA_INST_0_43036 : AO1A
      port map(A => HIEFFPLA_NET_0_119017, B => 
        HIEFFPLA_NET_0_119448, C => HIEFFPLA_NET_0_119404, Y => 
        HIEFFPLA_NET_0_119395);
    
    \U_TFC_SERDAT_SOURCE/SERDAT[6]\ : DFN1C0
      port map(D => \U_TFC_SERDAT_SOURCE/N_SERDAT[6]\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \TFC_TX_DAT[6]\);
    
    HIEFFPLA_INST_0_43631 : NAND3C
      port map(A => HIEFFPLA_NET_0_119234, B => 
        HIEFFPLA_NET_0_119259, C => HIEFFPLA_NET_0_119279, Y => 
        HIEFFPLA_NET_0_119262);
    
    HIEFFPLA_INST_0_56861 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_1[4]\, B => 
        HIEFFPLA_NET_0_116763, S => HIEFFPLA_NET_0_117600, Y => 
        HIEFFPLA_NET_0_116784);
    
    HIEFFPLA_INST_0_58578 : AND3
      port map(A => HIEFFPLA_NET_0_117215, B => 
        HIEFFPLA_NET_0_116649, C => HIEFFPLA_NET_0_116620, Y => 
        HIEFFPLA_NET_0_116502);
    
    \U_EXEC_MASTER/MPOR_B_17\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117787, CLK => CLK_40M_GL, CLR
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_1\, Q => 
        P_MASTER_POR_B_c_17);
    
    \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[10]\ : DFN1C0
      port map(D => \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\);
    
    HIEFFPLA_INST_0_50108 : AND2
      port map(A => CLK_40M_GL, B => 
        \U_ELK5_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0_net_1\, Y => 
        HIEFFPLA_NET_0_118014);
    
    \U50_PATTERNS/ELINK_ADDRA_6[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119966, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_4, Q => 
        \U50_PATTERNS/ELINK_ADDRA_6[1]\);
    
    \U50_PATTERNS/ELINK_ADDRA_10[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120085, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_22, Q => 
        \U50_PATTERNS/ELINK_ADDRA_10[2]\);
    
    HIEFFPLA_INST_0_50891 : MX2
      port map(A => HIEFFPLA_NET_0_117857, B => 
        HIEFFPLA_NET_0_117855, S => \BIT_OS_SEL_3[1]\, Y => 
        HIEFFPLA_NET_0_117867);
    
    HIEFFPLA_INST_0_47073 : MX2
      port map(A => \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[0]_net_1\, 
        B => \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\, S => 
        \BIT_OS_SEL_4[2]\, Y => HIEFFPLA_NET_0_118564);
    
    \U50_PATTERNS/ELINK_DINA_16[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119811, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_18, Q => 
        \U50_PATTERNS/ELINK_DINA_16[4]\);
    
    HIEFFPLA_INST_0_59682 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_2[2]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_18[2]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_1[4]_net_1\, Y
         => HIEFFPLA_NET_0_116362);
    
    HIEFFPLA_INST_0_48094 : MX2
      port map(A => 
        \U_ELK16_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]_net_1\, B => 
        \U_ELK16_CH/ELK_TX_DAT[6]\, S => 
        \U_ELK16_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118379);
    
    HIEFFPLA_INST_0_40702 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_15[4]\, B => 
        HIEFFPLA_NET_0_119570, S => HIEFFPLA_NET_0_119297, Y => 
        HIEFFPLA_NET_0_119819);
    
    \U50_PATTERNS/ELINK_DINA_3[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119767, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_11, Q => 
        \U50_PATTERNS/ELINK_DINA_3[0]\);
    
    HIEFFPLA_INST_0_44425 : XO1
      port map(A => \U50_PATTERNS/U4B_REGCROSS/SAMP_TWO[0]_net_1\, 
        B => \TFC_STOP_ADDR[0]\, C => HIEFFPLA_NET_0_119118, Y
         => HIEFFPLA_NET_0_119122);
    
    \U_ELK7_CH/U_ELK1_SERDAT_SOURCE/SERDAT[4]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117919, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_3, Q => 
        \U_ELK7_CH/ELK_TX_DAT[4]\);
    
    HIEFFPLA_INST_0_60153 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_7[0]\, B => 
        HIEFFPLA_NET_0_116680, S => HIEFFPLA_NET_0_117157, Y => 
        HIEFFPLA_NET_0_116303);
    
    HIEFFPLA_INST_0_57324 : XA1C
      port map(A => HIEFFPLA_NET_0_116709, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_3[8]\, C => 
        HIEFFPLA_NET_0_117179, Y => HIEFFPLA_NET_0_116699);
    
    HIEFFPLA_INST_0_42595 : XA1C
      port map(A => HIEFFPLA_NET_0_119521, B => 
        \U50_PATTERNS/REG_ADDR[5]\, C => HIEFFPLA_NET_0_119452, Y
         => HIEFFPLA_NET_0_119504);
    
    \U_ELK3_CH/U_SLAVE_1ELK/Q[11]\ : DFN1C0
      port map(D => \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/Q[11]_net_1\);
    
    \U50_PATTERNS/TFC_STRT_ADDR_T[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119158, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_5, Q => 
        \U50_PATTERNS/TFC_STRT_ADDR_T[6]\);
    
    HIEFFPLA_INST_0_60911 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_1[2]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_17[2]\, S
         => \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_3[4]_net_1\, 
        Y => HIEFFPLA_NET_0_116200);
    
    HIEFFPLA_INST_0_43077 : NAND2B
      port map(A => HIEFFPLA_NET_0_119003, B => 
        HIEFFPLA_NET_0_119420, Y => HIEFFPLA_NET_0_119385);
    
    \U200A_TFC/GP_PG_SM_0[10]\ : DFN1P0
      port map(D => HIEFFPLA_NET_0_120335, CLK => CLK_40M_GL, PRE
         => P_MASTER_POR_B_c_27_1, Q => 
        \U200A_TFC/GP_PG_SM_0[10]_net_1\);
    
    HIEFFPLA_INST_0_49455 : MX2
      port map(A => \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\, B
         => \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[12]_net_1\, S => 
        \BIT_OS_SEL_7[2]\, Y => HIEFFPLA_NET_0_118128);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_5[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_115992, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_15, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_5[3]\);
    
    HIEFFPLA_INST_0_41913 : NAND2B
      port map(A => HIEFFPLA_NET_0_119248, B => 
        HIEFFPLA_NET_0_119268, Y => HIEFFPLA_NET_0_119664);
    
    \U50_PATTERNS/ELINK_RWA[1]/U1\ : DFN1P0
      port map(D => HIEFFPLA_NET_0_119700, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_6, Q => \U50_PATTERNS/ELINK_RWA[1]\);
    
    HIEFFPLA_INST_0_38831 : MX2
      port map(A => HIEFFPLA_NET_0_119518, B => 
        \U50_PATTERNS/ELINK_ADDRA_13[5]\, S => 
        HIEFFPLA_NET_0_119285, Y => HIEFFPLA_NET_0_120058);
    
    \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_SEL_1[1]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_BIT_OS_VAL[1]\, CLK
         => CLK_40M_GL, CLR => P_MASTER_POR_B_c_27_0, Q => 
        \BIT_OS_SEL_1[1]\);
    
    HIEFFPLA_INST_0_37988 : MX2
      port map(A => \U200B_ELINKS/LOC_STRT_ADDR[1]\, B => 
        \ELKS_STRT_ADDR[1]\, S => 
        \U200B_ELINKS/GP_PG_SM_0[10]_net_1\, Y => 
        HIEFFPLA_NET_0_120178);
    
    HIEFFPLA_INST_0_56551 : AND3
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[5]_net_1\, B => 
        HIEFFPLA_NET_0_117426, C => HIEFFPLA_NET_0_117425, Y => 
        HIEFFPLA_NET_0_116840);
    
    \P_OP_MODE2_TE_pad/U0/U0\ : IOPAD_TRI_U
      port map(D => \P_OP_MODE2_TE_pad/U0/NET1\, E => 
        \P_OP_MODE2_TE_pad/U0/NET2\, PAD => P_OP_MODE2_TE);
    
    HIEFFPLA_INST_0_58419 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_14[0]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_30[0]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_3[4]_net_1\, Y
         => HIEFFPLA_NET_0_116524);
    
    HIEFFPLA_INST_0_37537 : NAND3B
      port map(A => HIEFFPLA_NET_0_120291, B => 
        \U200A_TFC/GP_PG_SM[1]_net_1\, C => \OP_MODE_c[2]\, Y => 
        HIEFFPLA_NET_0_120265);
    
    \U_ELK3_CH/U_SLAVE_1ELK/Q[4]\ : DFN1C0
      port map(D => \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/Q[4]_net_1\);
    
    HIEFFPLA_INST_0_54768 : NAND3
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[1]_net_1\, B => 
        HIEFFPLA_NET_0_117244, C => HIEFFPLA_NET_0_117251, Y => 
        HIEFFPLA_NET_0_117205);
    
    HIEFFPLA_INST_0_40163 : AOI1C
      port map(A => \U50_PATTERNS/ELINK_BLKA[7]\, B => 
        HIEFFPLA_NET_0_119640, C => HIEFFPLA_NET_0_119883, Y => 
        HIEFFPLA_NET_0_119884);
    
    HIEFFPLA_INST_0_40110 : AOI1D
      port map(A => HIEFFPLA_NET_0_119389, B => 
        HIEFFPLA_NET_0_119464, C => \U50_PATTERNS/SM_BANK_SEL[4]\, 
        Y => HIEFFPLA_NET_0_119903);
    
    \U_EXEC_MASTER/MPOR_B_11\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117787, CLK => CLK_40M_GL, CLR
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_1\, Q => 
        P_MASTER_POR_B_c_11);
    
    \U_ELK19_CH/U_ELK1_CMD_TX/SER_OUT_RI\ : DFN1C0
      port map(D => 
        \U_ELK19_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_0, Q => 
        \U_ELK19_CH/U_ELK1_CMD_TX/SER_OUT_RI_net_1\);
    
    \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[5]\ : DFN1C0
      port map(D => \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\);
    
    \U_ELK14_CH/U_SLAVE_1ELK/Q[11]\ : DFN1C0
      port map(D => \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/Q[11]_net_1\);
    
    HIEFFPLA_INST_0_44678 : MX2
      port map(A => \U50_PATTERNS/U4E_REGCROSS/LOCAL_REG_VAL[3]\, 
        B => \U50_PATTERNS/U4E_REGCROSS/SAMP_TWO[3]_net_1\, S => 
        HIEFFPLA_NET_0_119072, Y => HIEFFPLA_NET_0_119067);
    
    \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117041, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_17, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[4]\);
    
    HIEFFPLA_INST_0_37059 : AO1A
      port map(A => HIEFFPLA_NET_0_120337, B => 
        HIEFFPLA_NET_0_120325, C => HIEFFPLA_NET_0_120342, Y => 
        HIEFFPLA_NET_0_120355);
    
    HIEFFPLA_INST_0_38705 : MX2
      port map(A => HIEFFPLA_NET_0_119516, B => 
        \U50_PATTERNS/ELINK_ADDRA_11[7]\, S => 
        HIEFFPLA_NET_0_119280, Y => HIEFFPLA_NET_0_120072);
    
    \U_ELK2_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]\ : DFN1C0
      port map(D => \U_ELK2_CH/U_SLAVE_1ELK/Q[11]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]_net_1\);
    
    \U50_PATTERNS/U4B_REGCROSS/LOCAL_REG_VAL[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119132, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_19, Q => \TFC_STOP_ADDR[1]\);
    
    \U_TFC_CMD_TX/SER_CMD_WORD_F[1]\ : DFN1C0
      port map(D => \U_TFC_CMD_TX/N_SER_CMD_WORD_F[1]\, CLK => 
        CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_TFC_CMD_TX/SER_CMD_WORD_F[1]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_25[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116420, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_20, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_25[0]\);
    
    HIEFFPLA_INST_0_57258 : NAND3A
      port map(A => HIEFFPLA_NET_0_116713, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_3[0]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_3[4]\, Y => 
        HIEFFPLA_NET_0_116716);
    
    HIEFFPLA_INST_0_41656 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_9[6]\, B => 
        HIEFFPLA_NET_0_119566, S => HIEFFPLA_NET_0_119292, Y => 
        HIEFFPLA_NET_0_119713);
    
    \U_ELK13_CH/U_ELK1_SERDAT_SOURCE/SERDAT[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118505, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_4, Q => 
        \U_ELK13_CH/ELK_TX_DAT[3]\);
    
    HIEFFPLA_INST_0_49648 : MX2
      port map(A => \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\, B
         => \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\, S => 
        \BIT_OS_SEL_7[2]\, Y => HIEFFPLA_NET_0_118091);
    
    HIEFFPLA_INST_0_41350 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_5[4]\, B => 
        HIEFFPLA_NET_0_119570, S => HIEFFPLA_NET_0_119251, Y => 
        HIEFFPLA_NET_0_119747);
    
    \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[6]\ : DFN1C0
      port map(D => 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\);
    
    \U50_PATTERNS/U4A_REGCROSS/DELCNT[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119136, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_32, Q => 
        \U50_PATTERNS/U4A_REGCROSS/DELCNT[1]_net_1\);
    
    HIEFFPLA_INST_0_56754 : NAND3A
      port map(A => HIEFFPLA_NET_0_116805, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_0[5]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_0[6]\, Y => 
        HIEFFPLA_NET_0_116807);
    
    HIEFFPLA_INST_0_63131 : AX1A
      port map(A => HIEFFPLA_NET_0_115907, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[7]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[8]\, Y => 
        HIEFFPLA_NET_0_115880);
    
    HIEFFPLA_INST_0_46852 : AND2
      port map(A => \U_ELK11_CH/ELK_TX_DAT[1]\, B => 
        \U_ELK11_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118603);
    
    \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_2S_10\ : DFN1C0
      port map(D => 
        \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_1S_net_1\, CLK
         => CLK60MHZ, CLR => \U_EXEC_MASTER/P_MASTER_POR_B_c_0\, 
        Q => P_USB_MASTER_EN_c_10);
    
    \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[8]\ : DFN1C0
      port map(D => 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\);
    
    \U_ELK4_CH/U_ELK1_SERDAT_SOURCE/SERDAT[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118057, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_16, Q => 
        \U_ELK4_CH/ELK_TX_DAT[1]\);
    
    HIEFFPLA_INST_0_51832 : NAND2
      port map(A => \U_MASTER_DES/U13A_ADJ_160M/BITCNT[0]\, B => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[2]\, Y => 
        HIEFFPLA_NET_0_117682);
    
    \U_ELK2_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0\ : DFN1C0
      port map(D => CLK_40M_GL, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_8, Q => 
        \U_ELK2_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0_net_1\);
    
    HIEFFPLA_INST_0_60348 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_9[2]\, B => 
        HIEFFPLA_NET_0_116687, S => HIEFFPLA_NET_0_117393, Y => 
        HIEFFPLA_NET_0_116277);
    
    HIEFFPLA_INST_0_56818 : AND3
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_0[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_0[2]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_0[0]\, Y => 
        HIEFFPLA_NET_0_116790);
    
    HIEFFPLA_INST_0_46824 : MX2
      port map(A => \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[0]_net_1\, 
        B => \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\, S => 
        \BIT_OS_SEL_5[2]\, Y => HIEFFPLA_NET_0_118609);
    
    HIEFFPLA_INST_0_42989 : NAND3C
      port map(A => HIEFFPLA_NET_0_119418, B => 
        HIEFFPLA_NET_0_119489, C => HIEFFPLA_NET_0_119407, Y => 
        HIEFFPLA_NET_0_119408);
    
    HIEFFPLA_INST_0_51825 : NAND3C
      port map(A => \U_MASTER_DES/U13A_ADJ_160M/BITCNT[5]\, B => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[7]\, C => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[6]\, Y => 
        HIEFFPLA_NET_0_117685);
    
    HIEFFPLA_INST_0_40441 : MX2
      port map(A => HIEFFPLA_NET_0_119560, B => 
        \U50_PATTERNS/ELINK_DINA_11[7]\, S => 
        HIEFFPLA_NET_0_119280, Y => HIEFFPLA_NET_0_119848);
    
    \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[5]\ : DFN1C0
      port map(D => 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\);
    
    HIEFFPLA_INST_0_42606 : XA1C
      port map(A => HIEFFPLA_NET_0_119509, B => 
        \U50_PATTERNS/REG_ADDR[7]\, C => HIEFFPLA_NET_0_119452, Y
         => HIEFFPLA_NET_0_119502);
    
    \U_ELK11_CH/U_SLAVE_1ELK/Q[4]\ : DFN1C0
      port map(D => \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/Q[4]_net_1\);
    
    \U50_PATTERNS/CHKSUM[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120140, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_3, Q => \U50_PATTERNS/CHKSUM[3]\);
    
    HIEFFPLA_INST_0_42773 : AND3A
      port map(A => \U50_PATTERNS/REG_STATE_0[1]_net_1\, B => 
        HIEFFPLA_NET_0_119586, C => HIEFFPLA_NET_0_119430, Y => 
        HIEFFPLA_NET_0_119465);
    
    HIEFFPLA_INST_0_42300 : AOI1B
      port map(A => HIEFFPLA_NET_0_119559, B => 
        \U50_PATTERNS/RD_USB_ADBUS[4]\, C => 
        \U50_PATTERNS/RD_USB_ADBUS[5]\, Y => 
        HIEFFPLA_NET_0_119579);
    
    HIEFFPLA_INST_0_111646 : AO13
      port map(A => HIEFFPLA_NET_0_115835, B => 
        HIEFFPLA_NET_0_116982, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_SEQCNT[4]\, Y => 
        HIEFFPLA_NET_0_115951);
    
    HIEFFPLA_INST_0_56966 : XA1C
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_1[4]\, B => 
        HIEFFPLA_NET_0_116775, C => HIEFFPLA_NET_0_117179, Y => 
        HIEFFPLA_NET_0_116763);
    
    HIEFFPLA_INST_0_46269 : AND2
      port map(A => HIEFFPLA_NET_0_119476, B => 
        \U50_PATTERNS/CHKSUM[5]\, Y => HIEFFPLA_NET_0_118728);
    
    \U_ELK8_CH/U_SLAVE_1ELK/RECD_SER_WORD[5]\ : DFN1C0
      port map(D => \U_ELK8_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[5]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_8[5]\);
    
    \U_ELK14_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]\ : DFN1C0
      port map(D => \U_ELK14_CH/U_SLAVE_1ELK/Q[11]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]_net_1\);
    
    \U50_PATTERNS/U4B_REGCROSS/SAMP_ONE[1]\ : DFN1C0
      port map(D => \U50_PATTERNS/TFC_STOP_ADDR[1]\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_24_0, Q => 
        \U50_PATTERNS/U4B_REGCROSS/SAMP_ONE[1]_net_1\);
    
    HIEFFPLA_INST_0_38216 : MX2
      port map(A => \U50_PATTERNS/CHKSUM[7]\, B => 
        HIEFFPLA_NET_0_120128, S => HIEFFPLA_NET_0_119470, Y => 
        HIEFFPLA_NET_0_120136);
    
    HIEFFPLA_INST_0_38140 : AND3
      port map(A => HIEFFPLA_NET_0_120146, B => \ELKS_ADDRB[5]\, 
        C => \ELKS_ADDRB[4]\, Y => HIEFFPLA_NET_0_120144);
    
    \U_EXEC_MASTER/USB_MASTER_EN/TERMCNT_FG40M1S\ : DFN1C0
      port map(D => 
        \U_EXEC_MASTER/USB_MASTER_EN/TERMCNT_FG40M0S_net_1\, CLK
         => CLK_40M_GL, CLR => P_MASTER_POR_B_c_32_0, Q => 
        \U_EXEC_MASTER/USB_MASTER_EN/TERMCNT_FG40M1S_net_1\);
    
    \U_ELK8_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]\ : DFN1C0
      port map(D => \U_ELK8_CH/U_SLAVE_1ELK/Q[13]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]_net_1\);
    
    \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[7]\ : DFN1C0
      port map(D => 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\);
    
    \U50_PATTERNS/ELINKS_STOP_ADDR[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120125, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_14, Q => 
        \U50_PATTERNS/ELINKS_STOP_ADDR[2]\);
    
    HIEFFPLA_INST_0_45643 : NAND3C
      port map(A => HIEFFPLA_NET_0_118727, B => 
        HIEFFPLA_NET_0_118899, C => HIEFFPLA_NET_0_118873, Y => 
        HIEFFPLA_NET_0_118874);
    
    HIEFFPLA_INST_0_49668 : MX2
      port map(A => \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\, B
         => \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\, S => 
        \BIT_OS_SEL_7[2]\, Y => HIEFFPLA_NET_0_118088);
    
    HIEFFPLA_INST_0_58303 : MX2
      port map(A => HIEFFPLA_NET_0_116533, B => 
        HIEFFPLA_NET_0_116531, S => HIEFFPLA_NET_0_117367, Y => 
        HIEFFPLA_NET_0_116538);
    
    \U_ELK11_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL\ : DFN1C0
      port map(D => \U_ELK11_CH/ELK_IN_F_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL_net_1\);
    
    \U50_PATTERNS/ELINK_BLKA[4]/U1\ : DFN1P0
      port map(D => HIEFFPLA_NET_0_119921, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_19, Q => 
        \U50_PATTERNS/ELINK_BLKA[4]\);
    
    HIEFFPLA_INST_0_57231 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_3[6]\, B => 
        HIEFFPLA_NET_0_116701, S => HIEFFPLA_NET_0_117120, Y => 
        HIEFFPLA_NET_0_116719);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_3[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116007, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_11, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_3[3]\);
    
    HIEFFPLA_INST_0_37755 : NAND3C
      port map(A => \U200B_ELINKS/GP_PG_SM[0]_net_1\, B => 
        \U200B_ELINKS/GP_PG_SM[1]_net_1\, C => 
        HIEFFPLA_NET_0_120220, Y => HIEFFPLA_NET_0_120215);
    
    \U_EXEC_MASTER/MPOR_SALT_B_5\ : DFI1P0
      port map(D => HIEFFPLA_NET_0_117781, CLK => CLK_40M_GL, PRE
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_2\, QN => 
        MASTER_SALT_POR_B_i_0_i_5);
    
    \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[4]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[2]_net_1\, CLK => 
        CCC_160M_ADJ, CLR => P_MASTER_POR_B_c_34_0, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[4]_net_1\);
    
    HIEFFPLA_INST_0_40918 : MX2
      port map(A => HIEFFPLA_NET_0_119570, B => 
        \U50_PATTERNS/ELINK_DINA_18[4]\, S => 
        HIEFFPLA_NET_0_119264, Y => HIEFFPLA_NET_0_119795);
    
    HIEFFPLA_INST_0_52944 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_31[3]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_0[3]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_3[0]\, Y => 
        HIEFFPLA_NET_0_117485);
    
    \U_ELK11_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118606, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_11, Q => 
        \U_ELK11_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]_net_1\);
    
    HIEFFPLA_INST_0_43789 : AND3
      port map(A => HIEFFPLA_NET_0_119591, B => 
        \U50_PATTERNS/RD_USB_ADBUS[2]\, C => 
        \U50_PATTERNS/RD_USB_ADBUS[3]\, Y => 
        HIEFFPLA_NET_0_119214);
    
    HIEFFPLA_INST_0_38552 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_0[6]\, B => 
        HIEFFPLA_NET_0_119517, S => HIEFFPLA_NET_0_119272, Y => 
        HIEFFPLA_NET_0_120089);
    
    \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_2[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_115937, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_24_0, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_2[3]_net_1\);
    
    HIEFFPLA_INST_0_60336 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_9[2]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_25[2]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[4]_net_1\, Y
         => HIEFFPLA_NET_0_116279);
    
    HIEFFPLA_INST_0_52159 : AOI1D
      port map(A => \U_MASTER_DES/U13A_ADJ_160M/BITCNT[7]\, B => 
        HIEFFPLA_NET_0_117687, C => 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM[2]_net_1\, Y => 
        HIEFFPLA_NET_0_117620);
    
    HIEFFPLA_INST_0_51220 : MX2
      port map(A => \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\, B
         => \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[12]_net_1\, S => 
        \BIT_OS_SEL_3[2]\, Y => HIEFFPLA_NET_0_117810);
    
    \U_ELK10_CH/U_SLAVE_1ELK/Q[7]\ : DFN1C0
      port map(D => \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/Q[7]_net_1\);
    
    HIEFFPLA_INST_0_111821 : AX1E
      port map(A => HIEFFPLA_NET_0_117748, B => 
        \U_EXEC_MASTER/USB_MASTER_EN/T_CNT60M[6]_net_1\, C => 
        \U_EXEC_MASTER/USB_MASTER_EN/T_CNT60M[7]_net_1\, Y => 
        HIEFFPLA_NET_0_115829);
    
    HIEFFPLA_INST_0_45492 : AND3A
      port map(A => HIEFFPLA_NET_0_119437, B => 
        \U50_PATTERNS/WR_XFER_TYPE[2]_net_1\, C => 
        HIEFFPLA_NET_0_119367, Y => HIEFFPLA_NET_0_118903);
    
    HIEFFPLA_INST_0_45402 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_4[3]\, C => 
        \U50_PATTERNS/SM_BANK_SEL[15]\, Y => 
        HIEFFPLA_NET_0_118920);
    
    HIEFFPLA_INST_0_61574 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_7[1]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_23[1]\, S
         => \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[4]_net_1\, 
        Y => HIEFFPLA_NET_0_116107);
    
    HIEFFPLA_INST_0_43681 : NAND2B
      port map(A => \U50_PATTERNS/SM_BANK_SEL_0[21]\, B => 
        \U50_PATTERNS/SM_BANK_SEL[18]\, Y => 
        HIEFFPLA_NET_0_119243);
    
    \U_ELK1_CH/ELK_IN_R\ : DFN1C0
      port map(D => \AFLSDF_INV_63\, CLK => CCC_160M_ADJ, CLR => 
        DEV_RST_B_c, Q => \U_ELK1_CH/ELK_IN_R_net_1\);
    
    HIEFFPLA_INST_0_62574 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_7[3]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_8[3]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[0]\, Y => 
        HIEFFPLA_NET_0_115972);
    
    HIEFFPLA_INST_0_56148 : NAND3C
      port map(A => HIEFFPLA_NET_0_116939, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/MAX_CNT[4]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/MAX_CNT[5]\, Y => 
        HIEFFPLA_NET_0_116943);
    
    HIEFFPLA_INST_0_52486 : MX2
      port map(A => HIEFFPLA_NET_0_117505, B => 
        HIEFFPLA_NET_0_117501, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[3]\, Y => 
        HIEFFPLA_NET_0_117557);
    
    \U_ELK2_CH/U_SLAVE_1ELK/RECD_SER_WORD[1]\ : DFN1C0
      port map(D => \U_ELK2_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[1]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_2[1]\);
    
    \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[3]\ : DFN1C0
      port map(D => \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\);
    
    HIEFFPLA_INST_0_57750 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_6[5]\, B => 
        HIEFFPLA_NET_0_116610, S => HIEFFPLA_NET_0_117599, Y => 
        HIEFFPLA_NET_0_116627);
    
    HIEFFPLA_INST_0_51033 : MX2
      port map(A => HIEFFPLA_NET_0_117867, B => 
        HIEFFPLA_NET_0_117845, S => \BIT_OS_SEL_5[0]\, Y => 
        \U_ELK8_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[7]\);
    
    HIEFFPLA_INST_0_38786 : MX2
      port map(A => HIEFFPLA_NET_0_119524, B => 
        \U50_PATTERNS/ELINK_ADDRA_13[0]\, S => 
        HIEFFPLA_NET_0_119285, Y => HIEFFPLA_NET_0_120063);
    
    HIEFFPLA_INST_0_50965 : MX2
      port map(A => \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\, B
         => \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[12]_net_1\, S => 
        \BIT_OS_SEL_4[2]\, Y => HIEFFPLA_NET_0_117856);
    
    HIEFFPLA_INST_0_50358 : AND2A
      port map(A => \OP_MODE_c_0[1]\, B => \PATT_ELK_DAT_6[0]\, Y
         => HIEFFPLA_NET_0_117968);
    
    HIEFFPLA_INST_0_62448 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_5[0]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_6[0]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_2[0]\, Y => 
        HIEFFPLA_NET_0_115988);
    
    \U50_PATTERNS/ELINK_ADDRA_2[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119998, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_21, Q => 
        \U50_PATTERNS/ELINK_ADDRA_2[1]\);
    
    HIEFFPLA_INST_0_45677 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_15[5]\, C => 
        \U50_PATTERNS/SM_BANK_SEL[4]\, Y => HIEFFPLA_NET_0_118866);
    
    HIEFFPLA_INST_0_55628 : MX2
      port map(A => HIEFFPLA_NET_0_115988, B => 
        HIEFFPLA_NET_0_116240, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_1[3]\, Y => 
        HIEFFPLA_NET_0_117012);
    
    \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[3]\ : DFN1C0
      port map(D => 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[3]_net_1\);
    
    \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[1]\ : DFN1C0
      port map(D => 
        \U_ELK11_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\);
    
    HIEFFPLA_INST_0_43404 : MX2
      port map(A => \U50_PATTERNS/SM_BANK_SEL[16]\, B => 
        HIEFFPLA_NET_0_119221, S => HIEFFPLA_NET_0_118691, Y => 
        HIEFFPLA_NET_0_119315);
    
    HIEFFPLA_INST_0_54735 : AND3B
      port map(A => HIEFFPLA_NET_0_117247, B => 
        HIEFFPLA_NET_0_117252, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[1]_net_1\, Y => 
        HIEFFPLA_NET_0_117213);
    
    \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_2S_9\ : DFN1C0
      port map(D => 
        \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_1S_net_1\, CLK
         => CLK60MHZ, CLR => P_MASTER_POR_B_c_0_0, Q => 
        P_USB_MASTER_EN_c_9);
    
    HIEFFPLA_INST_0_50086 : MX2
      port map(A => 
        \U_ELK5_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]_net_1\, B => 
        \U_ELK5_CH/ELK_TX_DAT[6]\, S => 
        \U_ELK5_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118019);
    
    HIEFFPLA_INST_0_37692 : XO1
      port map(A => HIEFFPLA_NET_0_120146, B => \ELKS_ADDRB[4]\, 
        C => \U200B_ELINKS/GP_PG_SM[10]_net_1\, Y => 
        HIEFFPLA_NET_0_120229);
    
    \U_EXEC_MASTER/SYNC_BRD_RST_BI_0\ : DFI1P0
      port map(D => \U_EXEC_MASTER/DEV_RST_1B_i\, CLK => 
        CCC_160M_FXD, PRE => DEV_RST_B_c, QN => 
        \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_0\);
    
    HIEFFPLA_INST_0_55508 : MX2
      port map(A => HIEFFPLA_NET_0_116114, B => 
        HIEFFPLA_NET_0_116011, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[3]\, Y => 
        HIEFFPLA_NET_0_117028);
    
    HIEFFPLA_INST_0_38588 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_10[2]\, B => 
        HIEFFPLA_NET_0_119522, S => HIEFFPLA_NET_0_119239, Y => 
        HIEFFPLA_NET_0_120085);
    
    HIEFFPLA_INST_0_59353 : MX2
      port map(A => HIEFFPLA_NET_0_116398, B => 
        HIEFFPLA_NET_0_116396, S => HIEFFPLA_NET_0_117404, Y => 
        HIEFFPLA_NET_0_116402);
    
    \U_ELK0_CMD_TX/SER_CMD_WORD_R[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118663, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_14, Q => 
        \U_ELK0_CMD_TX/SER_CMD_WORD_R[2]_net_1\);
    
    \U_ELK4_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL\ : DFN1C0
      port map(D => \U_ELK4_CH/ELK_IN_F_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL_net_1\);
    
    HIEFFPLA_INST_0_59154 : AO1C
      port map(A => HIEFFPLA_NET_0_117208, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_24[2]\, C => 
        HIEFFPLA_NET_0_117249, Y => HIEFFPLA_NET_0_116428);
    
    \U_ELK19_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U0\ : IOPADP_BI
      port map(N2PIN => 
        \U_ELK19_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2_N2P\, D => 
        \U_ELK19_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, E => 
        \U_ELK19_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET2\, PAD => 
        ELK19_DAT_P, Y => 
        \U_ELK19_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\);
    
    \U_ELK10_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]\ : DFN1C0
      port map(D => \U_ELK10_CH/U_SLAVE_1ELK/Q[1]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]_net_1\);
    
    HIEFFPLA_INST_0_63169 : AND3
      port map(A => HIEFFPLA_NET_0_117226, B => 
        HIEFFPLA_NET_0_117222, C => HIEFFPLA_NET_0_117338, Y => 
        HIEFFPLA_NET_0_115869);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_7[5]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116598, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_14, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_7[5]\);
    
    \U_ELK14_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118467, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_2, Q => 
        \U_ELK14_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]_net_1\);
    
    HIEFFPLA_INST_0_63092 : AND2B
      port map(A => HIEFFPLA_NET_0_117078, B => 
        HIEFFPLA_NET_0_115882, Y => HIEFFPLA_NET_0_115890);
    
    HIEFFPLA_INST_0_60780 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_31[2]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_15[2]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[4]_net_1\, Y
         => HIEFFPLA_NET_0_116221);
    
    \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[0]\ : DFN1C0
      port map(D => 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[0]_net_1\);
    
    \U_ELK4_CH/U_ELK1_SERDAT_SOURCE/SERDAT[4]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118054, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_16, Q => 
        \U_ELK4_CH/ELK_TX_DAT[4]\);
    
    \U50_PATTERNS/U4B_REGCROSS/SAMP_ONE[7]\ : DFN1C0
      port map(D => \U50_PATTERNS/TFC_STOP_ADDR[7]\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_25, Q => 
        \U50_PATTERNS/U4B_REGCROSS/SAMP_ONE[7]_net_1\);
    
    HIEFFPLA_INST_0_45198 : NAND3C
      port map(A => HIEFFPLA_NET_0_118872, B => 
        HIEFFPLA_NET_0_118726, C => HIEFFPLA_NET_0_118796, Y => 
        HIEFFPLA_NET_0_118967);
    
    HIEFFPLA_INST_0_40184 : AOI1D
      port map(A => HIEFFPLA_NET_0_119389, B => 
        HIEFFPLA_NET_0_119464, C => \U50_PATTERNS/SM_BANK_SEL[8]\, 
        Y => HIEFFPLA_NET_0_119878);
    
    HIEFFPLA_INST_0_37680 : XO1
      port map(A => HIEFFPLA_NET_0_120145, B => \ELKS_ADDRB[2]\, 
        C => \U200B_ELINKS/GP_PG_SM[10]_net_1\, Y => 
        HIEFFPLA_NET_0_120232);
    
    \U_ELK12_CH/U_ELK1_SERDAT_SOURCE/SERDAT[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118550, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_2, Q => 
        \U_ELK12_CH/ELK_TX_DAT[3]\);
    
    HIEFFPLA_INST_0_49421 : MX2
      port map(A => \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\, B
         => \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\, S => 
        \BIT_OS_SEL_7[2]\, Y => HIEFFPLA_NET_0_118133);
    
    HIEFFPLA_INST_0_43337 : AND2
      port map(A => \U50_PATTERNS/SI_CNT[1]\, B => 
        \U50_PATTERNS/SI_CNT[0]\, Y => HIEFFPLA_NET_0_119323);
    
    HIEFFPLA_INST_0_52902 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_23[0]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_24[0]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_2[0]\, Y => 
        HIEFFPLA_NET_0_117492);
    
    HIEFFPLA_INST_0_46438 : AND3A
      port map(A => HIEFFPLA_NET_0_118693, B => 
        HIEFFPLA_NET_0_119392, C => 
        \U50_PATTERNS/WR_XFER_TYPE[1]_net_1\, Y => 
        HIEFFPLA_NET_0_118690);
    
    HIEFFPLA_INST_0_63190 : AND3
      port map(A => HIEFFPLA_NET_0_117226, B => 
        HIEFFPLA_NET_0_117222, C => HIEFFPLA_NET_0_117338, Y => 
        HIEFFPLA_NET_0_115866);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_13[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116540, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_12, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_13[2]\);
    
    \U_ELK5_CH/ELK_IN_F\ : DFN1C0
      port map(D => \U_ELK5_CH/ELK_IN_DDR_F\, CLK => CCC_160M_ADJ, 
        CLR => DEV_RST_B_c, Q => \U_ELK5_CH/ELK_IN_F_net_1\);
    
    \U_ELK10_CH/U_SLAVE_1ELK/Q[10]\ : DFN1C0
      port map(D => \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/Q[10]_net_1\);
    
    \U_ELK3_CH/U_ELK1_CMD_TX/SER_OUT_FI\ : DFI1C0
      port map(D => 
        \U_ELK3_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_14, QN
         => \U_ELK3_CH/U_ELK1_CMD_TX/SER_OUT_FI_i\);
    
    \U_ELK17_CH/ELK_IN_F\ : DFN1C0
      port map(D => \U_ELK17_CH/ELK_IN_DDR_F\, CLK => 
        CCC_160M_ADJ, CLR => DEV_RST_B_c, Q => 
        \U_ELK17_CH/ELK_IN_F_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_23[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116442, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_17_0, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_23[0]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_4[4]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116692, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_9, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_4[4]\);
    
    HIEFFPLA_INST_0_39470 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_3[4]\, B => 
        HIEFFPLA_NET_0_119519, S => HIEFFPLA_NET_0_119247, Y => 
        HIEFFPLA_NET_0_119987);
    
    HIEFFPLA_INST_0_39299 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_1[1]\, B => 
        HIEFFPLA_NET_0_119523, S => HIEFFPLA_NET_0_119243, Y => 
        HIEFFPLA_NET_0_120006);
    
    \U_ELK15_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL\ : DFN1C0
      port map(D => \U_ELK15_CH/ELK_IN_F_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL_net_1\);
    
    HIEFFPLA_INST_0_42271 : AND3
      port map(A => HIEFFPLA_NET_0_119424, B => 
        HIEFFPLA_NET_0_119595, C => HIEFFPLA_NET_0_119600, Y => 
        HIEFFPLA_NET_0_119584);
    
    HIEFFPLA_INST_0_60561 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_13[0]\, B => 
        HIEFFPLA_NET_0_117190, S => HIEFFPLA_NET_0_117137, Y => 
        HIEFFPLA_NET_0_116250);
    
    HIEFFPLA_INST_0_60492 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_11[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_12[1]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_4[0]\, Y => 
        HIEFFPLA_NET_0_116259);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_20[4]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116156, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_2, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_20[4]\);
    
    HIEFFPLA_INST_0_46120 : AO1
      port map(A => HIEFFPLA_NET_0_119244, B => 
        \U50_PATTERNS/ELINK_DOUTA_2[1]\, C => 
        HIEFFPLA_NET_0_118936, Y => HIEFFPLA_NET_0_118761);
    
    HIEFFPLA_INST_0_38233 : AND2A
      port map(A => HIEFFPLA_NET_0_119452, B => 
        \U50_PATTERNS/RD_USB_ADBUS[5]\, Y => 
        HIEFFPLA_NET_0_120130);
    
    \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[10]\ : DFN1C0
      port map(D => \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\);
    
    \U50_PATTERNS/OP_MODE_T[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119606, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_17, Q => 
        \U50_PATTERNS/OP_MODE_T[3]\);
    
    HIEFFPLA_INST_0_54773 : OR3B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[4]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[2]_net_1\, C => 
        HIEFFPLA_NET_0_117241, Y => HIEFFPLA_NET_0_117203);
    
    HIEFFPLA_INST_0_45473 : AO1
      port map(A => HIEFFPLA_NET_0_119276, B => 
        \U50_PATTERNS/ELINK_DOUTA_10[6]\, C => 
        HIEFFPLA_NET_0_118814, Y => HIEFFPLA_NET_0_118907);
    
    \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[7]\ : DFN1C0
      port map(D => 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\);
    
    \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[11]\ : DFN1C0
      port map(D => 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]_net_1\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[11]_net_1\);
    
    HIEFFPLA_INST_0_54784 : MX2
      port map(A => HIEFFPLA_NET_0_117261, B => 
        HIEFFPLA_NET_0_117353, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[1]_net_1\, Y => 
        HIEFFPLA_NET_0_117200);
    
    HIEFFPLA_INST_0_43659 : NAND2B
      port map(A => \U50_PATTERNS/SM_BANK_SEL[6]\, B => 
        \U50_PATTERNS/SM_BANK_SEL[10]\, Y => 
        HIEFFPLA_NET_0_119252);
    
    \U_ELK9_CH/U_ELK1_CMD_TX/SER_OUT_RI\ : DFN1C0
      port map(D => 
        \U_ELK9_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_13, Q
         => \U_ELK9_CH/U_ELK1_CMD_TX/SER_OUT_RI_net_1\);
    
    \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[3]\ : DFN1C0
      port map(D => \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\);
    
    \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[13]\ : DFN1C0
      port map(D => 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]_net_1\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[13]_net_1\);
    
    HIEFFPLA_INST_0_47421 : MX2
      port map(A => HIEFFPLA_NET_0_118485, B => 
        HIEFFPLA_NET_0_118499, S => \BIT_OS_SEL_3[1]\, Y => 
        HIEFFPLA_NET_0_118494);
    
    HIEFFPLA_INST_0_46784 : MX2
      port map(A => HIEFFPLA_NET_0_118634, B => 
        HIEFFPLA_NET_0_118630, S => \BIT_OS_SEL_0[0]\, Y => 
        \U_ELK10_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[5]\);
    
    HIEFFPLA_INST_0_44882 : AND3
      port map(A => HIEFFPLA_NET_0_119556, B => 
        HIEFFPLA_NET_0_119586, C => 
        \U50_PATTERNS/REG_STATE[2]_net_1\, Y => 
        HIEFFPLA_NET_0_119028);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_3[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116338, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_19, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_3[1]\);
    
    \U50_PATTERNS/ELINK_ADDRA_16[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120035, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_8, Q => 
        \U50_PATTERNS/ELINK_ADDRA_16[4]\);
    
    HIEFFPLA_INST_0_37816 : NAND3C
      port map(A => \U200B_ELINKS/GP_PG_SM[6]_net_1\, B => 
        \U200B_ELINKS/GP_PG_SM[7]_net_1\, C => \OP_MODE[4]\, Y
         => HIEFFPLA_NET_0_120201);
    
    \U_ELK9_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL\ : DFN1C0
      port map(D => 
        \U_ELK9_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL_net_1\);
    
    HIEFFPLA_INST_0_44560 : MX2
      port map(A => \ELKS_STOP_ADDR[1]\, B => 
        \U50_PATTERNS/U4D_REGCROSS/SAMP_TWO[1]_net_1\, S => 
        HIEFFPLA_NET_0_119093, Y => HIEFFPLA_NET_0_119090);
    
    HIEFFPLA_INST_0_46216 : AO1
      port map(A => HIEFFPLA_NET_0_119246, B => 
        \U50_PATTERNS/ELINK_DOUTA_3[3]\, C => 
        HIEFFPLA_NET_0_118910, Y => HIEFFPLA_NET_0_118741);
    
    HIEFFPLA_INST_0_45811 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/SM_BANK_SEL[3]\, C => 
        \U50_PATTERNS/ELINK_DOUTA_16[2]\, Y => 
        HIEFFPLA_NET_0_118835);
    
    \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_115929, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_9, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[1]\);
    
    HIEFFPLA_INST_0_61214 : MX2
      port map(A => HIEFFPLA_NET_0_117181, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_20[2]\, S => 
        HIEFFPLA_NET_0_117141, Y => HIEFFPLA_NET_0_116158);
    
    HIEFFPLA_INST_0_52081 : MX2C
      port map(A => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[10]_net_1\, B => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[11]_net_1\, S => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[0]\, Y => 
        HIEFFPLA_NET_0_117640);
    
    \U_ELK3_CH/U_SLAVE_1ELK/RECD_SER_WORD[3]\ : DFN1C0
      port map(D => \U_ELK3_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[3]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_3[3]\);
    
    HIEFFPLA_INST_0_37146 : XO1
      port map(A => \TFC_ADDRB[3]\, B => HIEFFPLA_NET_0_120261, C
         => \U200A_TFC/GP_PG_SM[10]_net_1\, Y => 
        HIEFFPLA_NET_0_120340);
    
    \U50_PATTERNS/U109_PATT_ELINK_BLK/DPRT_512X9_SRAM_R0C0\ : 
        RAM4K9
      generic map(MEMORYFILE => "DPRT_512X9_SRAM_R0C0.mem")

      port map(ADDRA11 => AFLSDF_GND, ADDRA10 => AFLSDF_GND, 
        ADDRA9 => AFLSDF_GND, ADDRA8 => \GND\, ADDRA7 => 
        \U50_PATTERNS/ELINK_ADDRA_9[7]\, ADDRA6 => 
        \U50_PATTERNS/ELINK_ADDRA_9[6]\, ADDRA5 => 
        \U50_PATTERNS/ELINK_ADDRA_9[5]\, ADDRA4 => 
        \U50_PATTERNS/ELINK_ADDRA_9[4]\, ADDRA3 => 
        \U50_PATTERNS/ELINK_ADDRA_9[3]\, ADDRA2 => 
        \U50_PATTERNS/ELINK_ADDRA_9[2]\, ADDRA1 => 
        \U50_PATTERNS/ELINK_ADDRA_9[1]\, ADDRA0 => 
        \U50_PATTERNS/ELINK_ADDRA_9[0]\, ADDRB11 => AFLSDF_GND, 
        ADDRB10 => AFLSDF_GND, ADDRB9 => AFLSDF_GND, ADDRB8 => 
        \GND\, ADDRB7 => \ELKS_ADDRB[7]\, ADDRB6 => 
        \ELKS_ADDRB[6]\, ADDRB5 => \ELKS_ADDRB[5]\, ADDRB4 => 
        \ELKS_ADDRB[4]\, ADDRB3 => \ELKS_ADDRB[3]\, ADDRB2 => 
        \ELKS_ADDRB[2]\, ADDRB1 => \ELKS_ADDRB[1]\, ADDRB0 => 
        \ELKS_ADDRB[0]\, DINA8 => \GND\, DINA7 => 
        \U50_PATTERNS/ELINK_DINA_9[7]\, DINA6 => 
        \U50_PATTERNS/ELINK_DINA_9[6]\, DINA5 => 
        \U50_PATTERNS/ELINK_DINA_9[5]\, DINA4 => 
        \U50_PATTERNS/ELINK_DINA_9[4]\, DINA3 => 
        \U50_PATTERNS/ELINK_DINA_9[3]\, DINA2 => 
        \U50_PATTERNS/ELINK_DINA_9[2]\, DINA1 => 
        \U50_PATTERNS/ELINK_DINA_9[1]\, DINA0 => 
        \U50_PATTERNS/ELINK_DINA_9[0]\, DINB8 => \GND\, DINB7 => 
        \ELK_RX_SER_WORD_9[7]\, DINB6 => \ELK_RX_SER_WORD_9[6]\, 
        DINB5 => \ELK_RX_SER_WORD_9[5]\, DINB4 => 
        \ELK_RX_SER_WORD_9[4]\, DINB3 => \ELK_RX_SER_WORD_9[3]\, 
        DINB2 => \ELK_RX_SER_WORD_9[2]\, DINB1 => 
        \ELK_RX_SER_WORD_9[1]\, DINB0 => \ELK_RX_SER_WORD_9[0]\, 
        WIDTHA0 => \VCC\, WIDTHA1 => \VCC\, WIDTHB0 => \VCC\, 
        WIDTHB1 => \VCC\, PIPEA => \VCC\, PIPEB => \VCC\, WMODEA
         => \GND\, WMODEB => \GND\, BLKA => 
        \U50_PATTERNS/ELINK_BLKA[9]\, BLKB => ELKS_RAM_BLKB_EN, 
        WENA => \U50_PATTERNS/ELINK_RWA[9]\, WENB => ELKS_RWB, 
        CLKA => CLK60MHZ, CLKB => CLK_40M_GL, RESET => 
        P_USB_MASTER_EN_c_0, DOUTA8 => OPEN, DOUTA7 => 
        \U50_PATTERNS/ELINK_DOUTA_9[7]\, DOUTA6 => 
        \U50_PATTERNS/ELINK_DOUTA_9[6]\, DOUTA5 => 
        \U50_PATTERNS/ELINK_DOUTA_9[5]\, DOUTA4 => 
        \U50_PATTERNS/ELINK_DOUTA_9[4]\, DOUTA3 => 
        \U50_PATTERNS/ELINK_DOUTA_9[3]\, DOUTA2 => 
        \U50_PATTERNS/ELINK_DOUTA_9[2]\, DOUTA1 => 
        \U50_PATTERNS/ELINK_DOUTA_9[1]\, DOUTA0 => 
        \U50_PATTERNS/ELINK_DOUTA_9[0]\, DOUTB8 => OPEN, DOUTB7
         => \PATT_ELK_DAT_9[7]\, DOUTB6 => \PATT_ELK_DAT_9[6]\, 
        DOUTB5 => \PATT_ELK_DAT_9[5]\, DOUTB4 => 
        \PATT_ELK_DAT_9[4]\, DOUTB3 => \PATT_ELK_DAT_9[3]\, 
        DOUTB2 => \PATT_ELK_DAT_9[2]\, DOUTB1 => 
        \PATT_ELK_DAT_9[1]\, DOUTB0 => \PATT_ELK_DAT_9[0]\);
    
    \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[4]\ : DFN1C0
      port map(D => 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\);
    
    HIEFFPLA_INST_0_61946 : MX2
      port map(A => HIEFFPLA_NET_0_117096, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_28[0]\, S => 
        HIEFFPLA_NET_0_117146, Y => HIEFFPLA_NET_0_116055);
    
    \U_ELK18_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]\ : DFN1C0
      port map(D => \U_ELK18_CH/U_SLAVE_1ELK/Q[1]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]_net_1\);
    
    \U_ELK6_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117970, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_6, Q => 
        \U_ELK6_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]_net_1\);
    
    \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[11]\ : DFN1C0
      port map(D => 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]_net_1\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[11]_net_1\);
    
    HIEFFPLA_INST_0_62878 : MX2
      port map(A => HIEFFPLA_NET_0_115898, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[10]\, S => 
        HIEFFPLA_NET_0_117073, Y => HIEFFPLA_NET_0_115933);
    
    HIEFFPLA_INST_0_62391 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_5[0]\, 
        B => HIEFFPLA_NET_0_117096, S => HIEFFPLA_NET_0_117172, Y
         => HIEFFPLA_NET_0_115995);
    
    \U_ELK8_CH/U_SLAVE_1ELK/Q[9]\ : DFN1C0
      port map(D => \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/Q[9]_net_1\);
    
    HIEFFPLA_INST_0_38110 : OA1A
      port map(A => HIEFFPLA_NET_0_120226, B => 
        \U200B_ELINKS/GP_PG_SM[10]_net_1\, C => \ELKS_ADDRB[0]\, 
        Y => HIEFFPLA_NET_0_120150);
    
    \U50_PATTERNS/REG_STATE[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119364, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_22_0, Q => 
        \U50_PATTERNS/REG_STATE[0]_net_1\);
    
    HIEFFPLA_INST_0_46383 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/SM_BANK_SEL[11]\, C => 
        \U50_PATTERNS/ELINK_DOUTA_8[1]\, Y => 
        HIEFFPLA_NET_0_118702);
    
    \U50_PATTERNS/OP_MODE_T[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119607, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_17, Q => 
        \U50_PATTERNS/OP_MODE_T[2]\);
    
    \U50_PATTERNS/ELINK_RWA[0]/U1\ : DFN1P0
      port map(D => HIEFFPLA_NET_0_119711, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_6, Q => \U50_PATTERNS/ELINK_RWA[0]\);
    
    HIEFFPLA_INST_0_42233 : NAND2A
      port map(A => \U50_PATTERNS/RD_USB_ADBUS[4]\, B => 
        \U50_PATTERNS/RD_USB_ADBUS[5]\, Y => 
        HIEFFPLA_NET_0_119596);
    
    \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_4[4]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_115935, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_24_0, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_4[4]_net_1\);
    
    \U50_PATTERNS/ELINK_ADDRA_18[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120016, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_12, Q => 
        \U50_PATTERNS/ELINK_ADDRA_18[7]\);
    
    HIEFFPLA_INST_0_63202 : MX2
      port map(A => \U_TFC_CMD_TX/SER_CMD_WORD_F[0]_net_1\, B => 
        \TFC_TX_DAT[2]\, S => \U_TFC_CMD_TX/START_RISE_net_1\, Y
         => \U_TFC_CMD_TX/N_SER_CMD_WORD_F[1]\);
    
    \U_ELK2_CH/U_ELK1_CMD_TX/SER_OUT_FI\ : DFN1C0
      port map(D => 
        \U_ELK2_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_5, Q => 
        \U_ELK2_CH/U_ELK1_CMD_TX/SER_OUT_FI_net_1\);
    
    HIEFFPLA_INST_0_51557 : AND2
      port map(A => 
        \U_EXEC_MASTER/USB_MASTER_EN/T_CNT60M[6]_net_1\, B => 
        \U_EXEC_MASTER/USB_MASTER_EN/T_CNT60M[5]_net_1\, Y => 
        HIEFFPLA_NET_0_117744);
    
    \U_ELK15_CH/U_ELK1_SERDAT_SOURCE/SERDAT[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118415, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_8, Q => 
        \U_ELK15_CH/ELK_TX_DAT[3]\);
    
    \U50_PATTERNS/U4B_REGCROSS/SAMP_ONE[6]\ : DFN1C0
      port map(D => \U50_PATTERNS/TFC_STOP_ADDR[6]\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_25, Q => 
        \U50_PATTERNS/U4B_REGCROSS/SAMP_ONE[6]_net_1\);
    
    HIEFFPLA_INST_0_50093 : MX2
      port map(A => 
        \U_ELK5_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]_net_1\, B => 
        \U_ELK5_CH/ELK_TX_DAT[3]\, S => 
        \U_ELK5_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118017);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_18[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116495, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_19, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_18[0]\);
    
    \U50_PATTERNS/U4C_REGCROSS/SAMP_TWO[1]\ : DFN1C0
      port map(D => \U50_PATTERNS/U4C_REGCROSS/SAMP_ONE[1]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_22_0, Q => 
        \U50_PATTERNS/U4C_REGCROSS/SAMP_TWO[1]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_17[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116501, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_18, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_17[0]\);
    
    \U50_PATTERNS/U4A_REGCROSS/SAMP_ONE[3]\ : DFN1C0
      port map(D => \U50_PATTERNS/TFC_STRT_ADDR[3]\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_32, Q => 
        \U50_PATTERNS/U4A_REGCROSS/SAMP_ONE[3]_net_1\);
    
    \U50_PATTERNS/ELINK_ADDRA_19[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120008, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_13, Q => 
        \U50_PATTERNS/ELINK_ADDRA_19[7]\);
    
    HIEFFPLA_INST_0_45322 : AO1
      port map(A => HIEFFPLA_NET_0_119277, B => 
        \U50_PATTERNS/ELINK_DOUTA_11[5]\, C => 
        HIEFFPLA_NET_0_118823, Y => HIEFFPLA_NET_0_118941);
    
    \U_ELK2_CH/U_ELK1_SERDAT_SOURCE/SERDAT[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118147, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_13, Q => 
        \U_ELK2_CH/ELK_TX_DAT[1]\);
    
    HIEFFPLA_INST_0_58133 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_10[2]\, B => 
        HIEFFPLA_NET_0_116687, S => HIEFFPLA_NET_0_117165, Y => 
        HIEFFPLA_NET_0_116560);
    
    \U_ELK5_CH/U_SLAVE_1ELK/RECD_SER_WORD[0]\ : DFN1C0
      port map(D => \U_ELK5_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[0]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_5[0]\);
    
    HIEFFPLA_INST_0_52319 : NAND3A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[1]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[0]_net_1\, C => 
        HIEFFPLA_NET_0_117594, Y => HIEFFPLA_NET_0_117582);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_18[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116494, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_19, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_18[1]\);
    
    AFLSDF_INV_42 : INV
      port map(A => DCB_SALT_SEL_c, Y => \AFLSDF_INV_42\);
    
    HIEFFPLA_INST_0_46580 : AND2A
      port map(A => \OP_MODE_c_4[1]\, B => \PATT_ELK_DAT_0[4]\, Y
         => HIEFFPLA_NET_0_118656);
    
    \U50_PATTERNS/SM_BANK_SEL[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119304, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_7, Q => 
        \U50_PATTERNS/SM_BANK_SEL[6]\);
    
    HIEFFPLA_INST_0_50688 : MX2
      port map(A => HIEFFPLA_NET_0_117907, B => 
        HIEFFPLA_NET_0_117903, S => \BIT_OS_SEL_4[1]\, Y => 
        HIEFFPLA_NET_0_117905);
    
    \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[10]\ : DFN1C0
      port map(D => 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\);
    
    HIEFFPLA_INST_0_52258 : AO1
      port map(A => HIEFFPLA_NET_0_117587, B => 
        HIEFFPLA_NET_0_117604, C => HIEFFPLA_NET_0_117179, Y => 
        HIEFFPLA_NET_0_117599);
    
    HIEFFPLA_INST_0_49114 : NAND2B
      port map(A => \OP_MODE_c_5[1]\, B => \PATT_ELK_DAT_1[1]\, Y
         => HIEFFPLA_NET_0_118192);
    
    \U_ELK9_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U0\ : IOPADP_BI
      port map(N2PIN => 
        \U_ELK9_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2_N2P\, D => 
        \U_ELK9_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, E => 
        \U_ELK9_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET2\, PAD => 
        ELK9_DAT_P, Y => 
        \U_ELK9_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\);
    
    HIEFFPLA_INST_0_60035 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_5[3]\, B => 
        HIEFFPLA_NET_0_116315, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_0[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116319);
    
    HIEFFPLA_INST_0_55160 : AND3
      port map(A => HIEFFPLA_NET_0_115918, B => 
        HIEFFPLA_NET_0_117065, C => HIEFFPLA_NET_0_115910, Y => 
        HIEFFPLA_NET_0_117108);
    
    HIEFFPLA_INST_0_47236 : MX2
      port map(A => \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[2]_net_1\, 
        B => \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\, S => 
        \BIT_OS_SEL_3[2]\, Y => HIEFFPLA_NET_0_118530);
    
    HIEFFPLA_INST_0_45076 : AND3A
      port map(A => \U50_PATTERNS/REG_STATE_0[2]_net_1\, B => 
        HIEFFPLA_NET_0_119378, C => 
        \U50_PATTERNS/REG_STATE_0[4]_net_1\, Y => 
        HIEFFPLA_NET_0_118986);
    
    HIEFFPLA_INST_0_38442 : MX2
      port map(A => \U50_PATTERNS/ELINKS_STRT_ADDR_T[1]\, B => 
        \U50_PATTERNS/RD_USB_ADBUS[1]\, S => 
        HIEFFPLA_NET_0_119493, Y => HIEFFPLA_NET_0_120102);
    
    \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[4]\ : DFN1C0
      port map(D => 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\);
    
    \P_CCC_160M_FXD_pad/U0/U1\ : IOTRI_OB_EB
      port map(D => CCC_160M_FXD, E => \VCC\, DOUT => 
        \P_CCC_160M_FXD_pad/U0/NET1\, EOUT => 
        \P_CCC_160M_FXD_pad/U0/NET2\);
    
    HIEFFPLA_INST_0_58685 : AO1B
      port map(A => HIEFFPLA_NET_0_117204, B => 
        HIEFFPLA_NET_0_116345, C => HIEFFPLA_NET_0_117231, Y => 
        HIEFFPLA_NET_0_116487);
    
    \U_ELK6_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0\ : DFN1C0
      port map(D => CLK_40M_GL, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_10, Q => 
        \U_ELK6_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0_net_1\);
    
    HIEFFPLA_INST_0_60241 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_8[1]\, B => 
        HIEFFPLA_NET_0_116677, S => HIEFFPLA_NET_0_117160, Y => 
        HIEFFPLA_NET_0_116292);
    
    HIEFFPLA_INST_0_39173 : MX2
      port map(A => HIEFFPLA_NET_0_119520, B => 
        \U50_PATTERNS/ELINK_ADDRA_18[3]\, S => 
        HIEFFPLA_NET_0_119264, Y => HIEFFPLA_NET_0_120020);
    
    \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[14]\ : DFN1C0
      port map(D => 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[14]_net_1\);
    
    HIEFFPLA_INST_0_42972 : AND3B
      port map(A => \U50_PATTERNS/REG_STATE[4]_net_1\, B => 
        HIEFFPLA_NET_0_119017, C => HIEFFPLA_NET_0_119375, Y => 
        HIEFFPLA_NET_0_119413);
    
    HIEFFPLA_INST_0_52982 : MX2
      port map(A => HIEFFPLA_NET_0_117464, B => 
        HIEFFPLA_NET_0_117460, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[2]\, Y => 
        HIEFFPLA_NET_0_117480);
    
    \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[12]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[10]_net_1\, CLK => 
        CCC_160M_ADJ, CLR => P_MASTER_POR_B_c_26, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[12]_net_1\);
    
    \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[7]\ : DFN1C0
      port map(D => \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\);
    
    \U_ELK12_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U0\ : IOPADP_BI
      port map(N2PIN => 
        \U_ELK12_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2_N2P\, D => 
        \U_ELK12_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, E => 
        \U_ELK12_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET2\, PAD => 
        ELK12_DAT_P, Y => 
        \U_ELK12_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\);
    
    HIEFFPLA_INST_0_43213 : AO1
      port map(A => HIEFFPLA_NET_0_119465, B => 
        HIEFFPLA_NET_0_119336, C => HIEFFPLA_NET_0_119335, Y => 
        HIEFFPLA_NET_0_119346);
    
    HIEFFPLA_INST_0_39929 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_9[7]\, B => 
        HIEFFPLA_NET_0_119516, S => HIEFFPLA_NET_0_119292, Y => 
        HIEFFPLA_NET_0_119936);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_5[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116319, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_1, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_5[3]\);
    
    \U50_PATTERNS/ELINK_ADDRA_18[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120017, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_12, Q => 
        \U50_PATTERNS/ELINK_ADDRA_18[6]\);
    
    HIEFFPLA_INST_0_40146 : AOI1D
      port map(A => HIEFFPLA_NET_0_119389, B => 
        HIEFFPLA_NET_0_119464, C => 
        \U50_PATTERNS/SM_BANK_SEL[16]\, Y => 
        HIEFFPLA_NET_0_119891);
    
    HIEFFPLA_INST_0_44670 : MX2
      port map(A => \OP_MODE_c[2]\, B => 
        \U50_PATTERNS/U4E_REGCROSS/SAMP_TWO[2]_net_1\, S => 
        HIEFFPLA_NET_0_119072, Y => HIEFFPLA_NET_0_119068);
    
    HIEFFPLA_INST_0_58754 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_19[1]\, B => 
        HIEFFPLA_NET_0_116677, S => HIEFFPLA_NET_0_117092, Y => 
        HIEFFPLA_NET_0_116480);
    
    \U_ELK17_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL\ : DFN1C0
      port map(D => 
        \U_ELK17_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL_net_1\);
    
    \U_ELK12_CH/U_ELK1_CMD_TX/SER_OUT_RI\ : DFN1C0
      port map(D => 
        \U_ELK12_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_10, Q
         => \U_ELK12_CH/U_ELK1_CMD_TX/SER_OUT_RI_net_1\);
    
    HIEFFPLA_INST_0_43117 : AND2B
      port map(A => \U50_PATTERNS/REG_STATE[2]_net_1\, B => 
        \U50_PATTERNS/REG_STATE[0]_net_1\, Y => 
        HIEFFPLA_NET_0_119370);
    
    \U_ELK15_CH/U_SLAVE_1ELK/RECD_SER_WORD[0]\ : DFN1C0
      port map(D => \U_ELK15_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[0]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_15[0]\);
    
    \U50_PATTERNS/ELINK_DINA_1[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119780, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_7, Q => 
        \U50_PATTERNS/ELINK_DINA_1[3]\);
    
    \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[12]\ : DFN1C0
      port map(D => 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[12]_net_1\);
    
    \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[13]\ : DFN1C0
      port map(D => \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\, 
        CLK => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[13]_net_1\);
    
    \U63_TS_SIWU_BUF/_TRIBUFF_F_24U[0]_/U0/U1\ : IOTRI_OB_EB
      port map(D => USB_SIWU_BI, E => P_USB_MASTER_EN_c, DOUT => 
        \U63_TS_SIWU_BUF/\\\\TRIBUFF_F_24U[0]\\\\/U0/NET1\, EOUT
         => \U63_TS_SIWU_BUF/\\\\TRIBUFF_F_24U[0]\\\\/U0/NET2\);
    
    \U_ELK18_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]\ : DFN1C0
      port map(D => \U_ELK18_CH/U_SLAVE_1ELK/Q[2]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]_net_1\);
    
    \U_ELK18_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL\ : DFN1C0
      port map(D => \U_ELK18_CH/ELK_IN_F_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL_net_1\);
    
    \U_ELK16_CH/U_SLAVE_1ELK/Q[1]\ : DFN1C0
      port map(D => \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/Q[1]_net_1\);
    
    \U_ELK13_CH/U_SLAVE_1ELK/Q[13]\ : DFN1C0
      port map(D => \U_ELK13_CH/U_SLAVE_1ELK/ADJ_Q[13]_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/Q[13]_net_1\);
    
    \U_ELK4_CH/ELK_IN_F\ : DFN1C0
      port map(D => \AFLSDF_INV_64\, CLK => CCC_160M_ADJ, CLR => 
        DEV_RST_B_c, Q => \U_ELK4_CH/ELK_IN_F_net_1\);
    
    \U_ELK11_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118607, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_11, Q => 
        \U_ELK11_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]_net_1\);
    
    HIEFFPLA_INST_0_47469 : MX2
      port map(A => HIEFFPLA_NET_0_118491, B => 
        HIEFFPLA_NET_0_118488, S => \BIT_OS_SEL_3[1]\, Y => 
        HIEFFPLA_NET_0_118487);
    
    \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[9]\ : DFN1C0
      port map(D => \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\);
    
    HIEFFPLA_INST_0_62813 : XA1B
      port map(A => HIEFFPLA_NET_0_115876, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[2]_net_1\, C => 
        HIEFFPLA_NET_0_117102, Y => HIEFFPLA_NET_0_115943);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_21[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116143, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_3, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_21[2]\);
    
    HIEFFPLA_INST_0_46929 : MX2
      port map(A => HIEFFPLA_NET_0_118585, B => 
        HIEFFPLA_NET_0_118581, S => \BIT_OS_SEL_5[1]\, Y => 
        HIEFFPLA_NET_0_118583);
    
    HIEFFPLA_INST_0_41897 : AOI1C
      port map(A => \U50_PATTERNS/ELINK_RWA[7]\, B => 
        HIEFFPLA_NET_0_119640, C => HIEFFPLA_NET_0_119669, Y => 
        HIEFFPLA_NET_0_119670);
    
    HIEFFPLA_INST_0_41744 : MX2
      port map(A => HIEFFPLA_NET_0_119680, B => 
        \U50_PATTERNS/ELINK_RWA[19]\, S => 
        \U50_PATTERNS/SM_BANK_SEL_0[20]\, Y => 
        HIEFFPLA_NET_0_119701);
    
    HIEFFPLA_INST_0_51482 : MX2
      port map(A => HIEFFPLA_NET_0_117759, B => 
        \U_EXEC_MASTER/PRESCALE[2]\, S => HIEFFPLA_NET_0_117787, 
        Y => HIEFFPLA_NET_0_117766);
    
    HIEFFPLA_INST_0_55786 : MX2
      port map(A => HIEFFPLA_NET_0_116996, B => 
        HIEFFPLA_NET_0_116981, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[4]\, Y => 
        HIEFFPLA_NET_0_116990);
    
    \U_ELK9_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]\ : DFN1C0
      port map(D => \U_ELK9_CH/U_SLAVE_1ELK/Q[5]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]_net_1\);
    
    \U_ELK8_CH/U_SLAVE_1ELK/Q[13]\ : DFN1C0
      port map(D => \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[13]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/Q[13]_net_1\);
    
    \U200A_TFC/LOC_STRT_ADDR[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120276, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_5, Q => \U200A_TFC/LOC_STRT_ADDR[6]\);
    
    HIEFFPLA_INST_0_37929 : AO1C
      port map(A => \U200B_ELINKS/N_232_li\, B => ALIGN_ACTIVE, C
         => P_USB_MASTER_EN_c, Y => HIEFFPLA_NET_0_120188);
    
    \U_ELK5_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118022, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_5, Q => 
        \U_ELK5_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]_net_1\);
    
    HIEFFPLA_INST_0_61073 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_19[3]\, B => 
        HIEFFPLA_NET_0_117075, S => HIEFFPLA_NET_0_117170, Y => 
        HIEFFPLA_NET_0_116177);
    
    HIEFFPLA_INST_0_60630 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_13[3]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_29[3]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_2[4]_net_1\, Y
         => HIEFFPLA_NET_0_116241);
    
    HIEFFPLA_INST_0_60375 : MX2
      port map(A => HIEFFPLA_NET_0_117114, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_10[1]\, S => 
        HIEFFPLA_NET_0_117154, Y => HIEFFPLA_NET_0_116274);
    
    HIEFFPLA_INST_0_62073 : MX2
      port map(A => HIEFFPLA_NET_0_116135, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_29[2]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_2[3]\, Y => 
        HIEFFPLA_NET_0_116039);
    
    HIEFFPLA_INST_0_39380 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_2[2]\, B => 
        HIEFFPLA_NET_0_119522, S => HIEFFPLA_NET_0_119278, Y => 
        HIEFFPLA_NET_0_119997);
    
    \U_ELK6_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]\ : DFN1C0
      port map(D => \U_ELK6_CH/U_SLAVE_1ELK/Q[4]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]_net_1\);
    
    HIEFFPLA_INST_0_53807 : NAND3C
      port map(A => HIEFFPLA_NET_0_116773, B => 
        HIEFFPLA_NET_0_117310, C => HIEFFPLA_NET_0_117407, Y => 
        HIEFFPLA_NET_0_117349);
    
    \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[0]\ : DFN1C0
      port map(D => 
        \U_ELK18_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\);
    
    HIEFFPLA_INST_0_61424 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_22[2]\, B => 
        HIEFFPLA_NET_0_117181, S => HIEFFPLA_NET_0_117080, Y => 
        HIEFFPLA_NET_0_116128);
    
    \U_ELK13_CH/U_ELK1_SERDAT_SOURCE/SERDAT[6]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118502, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_4, Q => 
        \U_ELK13_CH/ELK_TX_DAT[6]\);
    
    HIEFFPLA_INST_0_59574 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_29[2]\, B => 
        HIEFFPLA_NET_0_116369, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_0[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116376);
    
    HIEFFPLA_INST_0_60902 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_17[4]\, B => 
        HIEFFPLA_NET_0_117166, S => HIEFFPLA_NET_0_117169, Y => 
        HIEFFPLA_NET_0_116201);
    
    HIEFFPLA_INST_0_46222 : AO1
      port map(A => HIEFFPLA_NET_0_119276, B => 
        \U50_PATTERNS/ELINK_DOUTA_10[4]\, C => 
        HIEFFPLA_NET_0_118909, Y => HIEFFPLA_NET_0_118739);
    
    HIEFFPLA_INST_0_38225 : AND2A
      port map(A => HIEFFPLA_NET_0_119452, B => 
        \U50_PATTERNS/RD_USB_ADBUS[1]\, Y => 
        HIEFFPLA_NET_0_120134);
    
    HIEFFPLA_INST_0_51409 : NAND2A
      port map(A => HIEFFPLA_NET_0_117778, B => 
        \U_EXEC_MASTER/DEL_CNT[3]\, Y => HIEFFPLA_NET_0_117782);
    
    HIEFFPLA_INST_0_44317 : XO1
      port map(A => \U50_PATTERNS/U4A_REGCROSS/SAMP_TWO[1]_net_1\, 
        B => \TFC_STRT_ADDR[1]\, C => HIEFFPLA_NET_0_119140, Y
         => HIEFFPLA_NET_0_119144);
    
    \U_ELK8_CH/U_SLAVE_1ELK/RECD_SER_WORD[0]\ : DFN1C0
      port map(D => \U_ELK8_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[0]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_8[0]\);
    
    \U_ELK9_CH/U_SLAVE_1ELK/Q[10]\ : DFN1C0
      port map(D => \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/Q[10]_net_1\);
    
    HIEFFPLA_INST_0_52353 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_BIT_OS_VAL[3]\, B
         => HIEFFPLA_NET_0_117573, S => HIEFFPLA_NET_0_117111, Y
         => HIEFFPLA_NET_0_117577);
    
    \U_ELK2_CH/U_ELK1_SERDAT_SOURCE/SERDAT[4]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118144, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_13, Q => 
        \U_ELK2_CH/ELK_TX_DAT[4]\);
    
    AFLSDF_INV_31 : INV
      port map(A => DCB_SALT_SEL_c, Y => \AFLSDF_INV_31\);
    
    \U_ELK19_CH/U_SLAVE_1ELK/Q[5]\ : DFN1C0
      port map(D => \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/Q[5]_net_1\);
    
    HIEFFPLA_INST_0_52154 : AND2
      port map(A => 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM[5]_net_1\, B => 
        HIEFFPLA_NET_0_117689, Y => HIEFFPLA_NET_0_117622);
    
    HIEFFPLA_INST_0_60280 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_8[2]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_24[2]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_1[4]_net_1\, Y
         => HIEFFPLA_NET_0_116287);
    
    HIEFFPLA_INST_0_45995 : AND3B
      port map(A => HIEFFPLA_NET_0_119426, B => 
        HIEFFPLA_NET_0_119379, C => \U50_PATTERNS/OP_MODE[0]\, Y
         => HIEFFPLA_NET_0_118794);
    
    HIEFFPLA_INST_0_49499 : MX2
      port map(A => HIEFFPLA_NET_0_118137, B => 
        HIEFFPLA_NET_0_118134, S => \BIT_OS_SEL_1[0]\, Y => 
        \U_ELK2_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[2]\);
    
    HIEFFPLA_INST_0_45905 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/SM_BANK_SEL[13]\, C => 
        \U50_PATTERNS/ELINK_DOUTA_6[5]\, Y => 
        HIEFFPLA_NET_0_118815);
    
    \U_ELK5_CH/U_ELK1_CMD_TX/SER_OUT_FDEL\ : DFN1C0
      port map(D => \U_ELK5_CH/U_ELK1_CMD_TX/SER_OUT_FI_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_8, Q
         => \U_ELK5_CH/ELK_OUT_F\);
    
    HIEFFPLA_INST_0_55500 : MX2
      port map(A => HIEFFPLA_NET_0_116991, B => 
        HIEFFPLA_NET_0_117034, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[2]\, Y => 
        HIEFFPLA_NET_0_117029);
    
    HIEFFPLA_INST_0_46185 : AO1
      port map(A => HIEFFPLA_NET_0_119288, B => 
        \U50_PATTERNS/ELINK_DOUTA_16[6]\, C => 
        HIEFFPLA_NET_0_118924, Y => HIEFFPLA_NET_0_118747);
    
    HIEFFPLA_INST_0_50899 : MX2
      port map(A => \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[1]_net_1\, B
         => \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\, S => 
        \BIT_OS_SEL_3[2]\, Y => HIEFFPLA_NET_0_117866);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_4[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_115998, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_13, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_4[2]\);
    
    \U_ELK14_CH/U_ELK1_CMD_TX/START_RISE\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118464, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_0, Q => 
        \U_ELK14_CH/U_ELK1_CMD_TX/START_RISE_net_1\);
    
    \U50_PATTERNS/ELINK_ADDRA_9[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119940, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_10, Q => 
        \U50_PATTERNS/ELINK_ADDRA_9[3]\);
    
    HIEFFPLA_INST_0_57561 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_5[3]\, B => 
        HIEFFPLA_NET_0_116642, S => HIEFFPLA_NET_0_117121, Y => 
        HIEFFPLA_NET_0_116658);
    
    HIEFFPLA_INST_0_52896 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_27[3]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_28[3]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_1[0]\, Y => 
        HIEFFPLA_NET_0_117493);
    
    \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[12]\ : DFN1C0
      port map(D => 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]_net_1\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[12]_net_1\);
    
    HIEFFPLA_INST_0_55906 : MX2
      port map(A => HIEFFPLA_NET_0_116001, B => 
        HIEFFPLA_NET_0_116257, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[3]\, Y => 
        HIEFFPLA_NET_0_116975);
    
    HIEFFPLA_INST_0_55366 : NAND3
      port map(A => HIEFFPLA_NET_0_115902, B => 
        HIEFFPLA_NET_0_115900, C => HIEFFPLA_NET_0_115915, Y => 
        HIEFFPLA_NET_0_117049);
    
    HIEFFPLA_INST_0_61064 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_19[2]\, B => 
        HIEFFPLA_NET_0_117131, S => HIEFFPLA_NET_0_117170, Y => 
        HIEFFPLA_NET_0_116178);
    
    HIEFFPLA_INST_0_58073 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_0[3]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_16[3]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_1[4]_net_1\, Y
         => HIEFFPLA_NET_0_116568);
    
    \U_ELK15_CH/U_SLAVE_1ELK/Q[3]\ : DFN1C0
      port map(D => \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/Q[3]_net_1\);
    
    HIEFFPLA_INST_0_58604 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_17[2]\, B => 
        HIEFFPLA_NET_0_116687, S => HIEFFPLA_NET_0_117161, Y => 
        HIEFFPLA_NET_0_116499);
    
    HIEFFPLA_INST_0_40396 : MX2
      port map(A => HIEFFPLA_NET_0_119575, B => 
        \U50_PATTERNS/ELINK_DINA_11[2]\, S => 
        HIEFFPLA_NET_0_119280, Y => HIEFFPLA_NET_0_119853);
    
    \U_ELK9_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]\ : DFN1C0
      port map(D => \U_ELK9_CH/U_SLAVE_1ELK/Q[4]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]_net_1\);
    
    \U_ELK13_CH/U_SLAVE_1ELK/RECD_SER_WORD[5]\ : DFN1C0
      port map(D => \U_ELK13_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[5]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_13[5]\);
    
    \U50_PATTERNS/REG_ADDR[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119530, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_10, Q => \U50_PATTERNS/REG_ADDR[3]\);
    
    HIEFFPLA_INST_0_60998 : MX2
      port map(A => HIEFFPLA_NET_0_117186, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_18[3]\, S => 
        HIEFFPLA_NET_0_117134, Y => HIEFFPLA_NET_0_116187);
    
    \U_ELK0_SERDAT_SOURCE/SERDAT[6]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118654, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_10, Q => \ELK0_TX_DAT[6]\);
    
    \U50_PATTERNS/U4E_REGCROSS/SAMP_TWO[2]\ : DFN1C0
      port map(D => \U50_PATTERNS/U4E_REGCROSS/SAMP_ONE[2]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_23, Q => 
        \U50_PATTERNS/U4E_REGCROSS/SAMP_TWO[2]_net_1\);
    
    HIEFFPLA_INST_0_53471 : AOI1D
      port map(A => HIEFFPLA_NET_0_116686, B => 
        HIEFFPLA_NET_0_116649, C => HIEFFPLA_NET_0_117337, Y => 
        HIEFFPLA_NET_0_117403);
    
    \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[2]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[0]_net_1\, CLK => 
        CCC_160M_ADJ, CLR => P_MASTER_POR_B_c_34_0, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[2]_net_1\);
    
    \U_ELK4_CH/U_SLAVE_1ELK/Q[10]\ : DFN1C0
      port map(D => \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/Q[10]_net_1\);
    
    HIEFFPLA_INST_0_62057 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_29[4]\, B => 
        HIEFFPLA_NET_0_117100, S => HIEFFPLA_NET_0_117072, Y => 
        HIEFFPLA_NET_0_116041);
    
    HIEFFPLA_INST_0_38031 : AO1A
      port map(A => HIEFFPLA_NET_0_120221, B => 
        HIEFFPLA_NET_0_120220, C => HIEFFPLA_NET_0_120165, Y => 
        HIEFFPLA_NET_0_120170);
    
    HIEFFPLA_INST_0_62328 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_3[1]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_4[1]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_4[0]\, Y => 
        HIEFFPLA_NET_0_116003);
    
    \U_MASTER_DES/U13A_ADJ_160M/CCC1_MODE\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117671, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_25, Q => \U_MASTER_DES/AUX_MODE\);
    
    \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[10]\ : DFN1C0
      port map(D => 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\);
    
    \U50_PATTERNS/ELINK_ADDRA_4[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119979, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_2_0, Q => 
        \U50_PATTERNS/ELINK_ADDRA_4[4]\);
    
    HIEFFPLA_INST_0_62146 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_30[0]\, B => 
        HIEFFPLA_NET_0_117190, S => HIEFFPLA_NET_0_117330, Y => 
        HIEFFPLA_NET_0_116030);
    
    HIEFFPLA_INST_0_49688 : MX2
      port map(A => \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\, B
         => \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[12]_net_1\, S => 
        \BIT_OS_SEL_7[2]\, Y => HIEFFPLA_NET_0_118085);
    
    \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[6]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117099, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_27, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[6]_net_1\);
    
    \U_ELK19_CH/U_SLAVE_1ELK/Q[10]\ : DFN1C0
      port map(D => \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/Q[10]_net_1\);
    
    \U_ELK18_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]\ : DFN1C0
      port map(D => \U_ELK18_CH/U_SLAVE_1ELK/Q[0]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]_net_1\);
    
    HIEFFPLA_INST_0_52534 : MX2
      port map(A => HIEFFPLA_NET_0_117491, B => 
        HIEFFPLA_NET_0_117487, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_2[3]\, Y => 
        HIEFFPLA_NET_0_117551);
    
    HIEFFPLA_INST_0_41927 : AND3C
      port map(A => HIEFFPLA_NET_0_119245, B => 
        HIEFFPLA_NET_0_119262, C => \U50_PATTERNS/SM_BANK_SEL[3]\, 
        Y => HIEFFPLA_NET_0_119659);
    
    HIEFFPLA_INST_0_49373 : MX2
      port map(A => HIEFFPLA_NET_0_118131, B => 
        HIEFFPLA_NET_0_118128, S => \BIT_OS_SEL[1]\, Y => 
        HIEFFPLA_NET_0_118140);
    
    HIEFFPLA_INST_0_51713 : NAND2B
      port map(A => 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM[4]_net_1\, B => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[39]_net_1\, Y => 
        HIEFFPLA_NET_0_117713);
    
    HIEFFPLA_INST_0_42064 : NAND3C
      port map(A => HIEFFPLA_NET_0_119438, B => 
        HIEFFPLA_NET_0_119366, C => HIEFFPLA_NET_0_119437, Y => 
        HIEFFPLA_NET_0_119622);
    
    \U50_PATTERNS/U4A_REGCROSS/SAMP_TWO[6]\ : DFN1C0
      port map(D => \U50_PATTERNS/U4A_REGCROSS/SAMP_ONE[6]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_22, Q => 
        \U50_PATTERNS/U4A_REGCROSS/SAMP_TWO[6]_net_1\);
    
    \U50_PATTERNS/TFC_ADDRA[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119207, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_9, Q => \U50_PATTERNS/TFC_ADDRA[0]\);
    
    HIEFFPLA_INST_0_49531 : MX2
      port map(A => HIEFFPLA_NET_0_118140, B => 
        HIEFFPLA_NET_0_118132, S => \BIT_OS_SEL_1[0]\, Y => 
        \U_ELK2_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[6]\);
    
    HIEFFPLA_INST_0_49200 : MX2
      port map(A => \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\, B
         => \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[11]_net_1\, S => 
        \BIT_OS_SEL[2]\, Y => HIEFFPLA_NET_0_118174);
    
    HIEFFPLA_INST_0_48816 : MX2
      port map(A => \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[0]_net_1\, 
        B => \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\, S => 
        \BIT_OS_SEL_0[2]\, Y => HIEFFPLA_NET_0_118249);
    
    \U50_PATTERNS/U4C_REGCROSS/SAMP_TWO[3]\ : DFN1C0
      port map(D => \U50_PATTERNS/U4C_REGCROSS/SAMP_ONE[3]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_22_0, Q => 
        \U50_PATTERNS/U4C_REGCROSS/SAMP_TWO[3]_net_1\);
    
    HIEFFPLA_INST_0_51423 : NAND3
      port map(A => \U_EXEC_MASTER/DEL_CNT[0]\, B => 
        \U_EXEC_MASTER/DEL_CNT[1]\, C => 
        \U_EXEC_MASTER/DEL_CNT[2]\, Y => HIEFFPLA_NET_0_117778);
    
    HIEFFPLA_INST_0_41934 : NAND2B
      port map(A => \U50_PATTERNS/ELINK_RWA[15]\, B => 
        HIEFFPLA_NET_0_119654, Y => HIEFFPLA_NET_0_119655);
    
    HIEFFPLA_INST_0_39560 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_4[6]\, B => 
        HIEFFPLA_NET_0_119517, S => HIEFFPLA_NET_0_119284, Y => 
        HIEFFPLA_NET_0_119977);
    
    \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[3]\\\\/U0/U0\ : 
        IOPAD_BI_U
      port map(D => 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[3]\\\\/U0/NET1\, 
        E => 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[3]\\\\/U0/NET2\, 
        Y => 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[3]\\\\/U0/NET3\, 
        PAD => BIDIR_USB_ADBUS(3));
    
    HIEFFPLA_INST_0_57202 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_3[3]\, B => 
        HIEFFPLA_NET_0_116705, S => HIEFFPLA_NET_0_117120, Y => 
        HIEFFPLA_NET_0_116722);
    
    HIEFFPLA_INST_0_47126 : AND2A
      port map(A => \OP_MODE_c_3[1]\, B => \PATT_ELK_DAT_12[5]\, 
        Y => HIEFFPLA_NET_0_118548);
    
    HIEFFPLA_INST_0_41035 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_1[1]\, B => 
        HIEFFPLA_NET_0_119576, S => HIEFFPLA_NET_0_119243, Y => 
        HIEFFPLA_NET_0_119782);
    
    \U_ELK8_CH/U_SLAVE_1ELK/Q[0]\ : DFN1C0
      port map(D => \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/Q[0]_net_1\);
    
    HIEFFPLA_INST_0_56953 : AND3B
      port map(A => HIEFFPLA_NET_0_117179, B => 
        HIEFFPLA_NET_0_116758, C => HIEFFPLA_NET_0_116769, Y => 
        HIEFFPLA_NET_0_116766);
    
    HIEFFPLA_INST_0_39704 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_6[6]\, B => 
        HIEFFPLA_NET_0_119517, S => HIEFFPLA_NET_0_119258, Y => 
        HIEFFPLA_NET_0_119961);
    
    \U50_PATTERNS/U4C_REGCROSS/LOCAL_REG_VAL[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119110, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_21, Q => \ELKS_STRT_ADDR[2]\);
    
    \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[6]\ : DFN1C0
      port map(D => 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\);
    
    \U200B_ELINKS/LOC_STRT_ADDR[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120172, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_12, Q => 
        \U200B_ELINKS/LOC_STRT_ADDR[7]\);
    
    HIEFFPLA_INST_0_61910 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_11[3]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_27[3]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_2[4]_net_1\, Y
         => HIEFFPLA_NET_0_116061);
    
    \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[4]\ : DFN1C0
      port map(D => \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\);
    
    HIEFFPLA_INST_0_56751 : NAND3C
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_0[6]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_0[5]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_0[4]\, Y => 
        HIEFFPLA_NET_0_116808);
    
    \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[1]\ : DFN1C0
      port map(D => 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[1]_net_1\);
    
    HIEFFPLA_INST_0_37082 : XO1
      port map(A => HIEFFPLA_NET_0_120257, B => \TFC_ADDRB[2]\, C
         => \U200A_TFC/GP_PG_SM[10]_net_1\, Y => 
        HIEFFPLA_NET_0_120351);
    
    \U_ELK12_CH/U_ELK1_CMD_TX/SER_OUT_FDEL\ : DFN1C0
      port map(D => \U_ELK12_CH/U_ELK1_CMD_TX/SER_OUT_FI_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_12, Q
         => \U_ELK12_CH/ELK_OUT_F\);
    
    HIEFFPLA_INST_0_46626 : NAND2B
      port map(A => \OP_MODE_c_3[1]\, B => \PATT_ELK_DAT_10[3]\, 
        Y => HIEFFPLA_NET_0_118640);
    
    \U_ELK9_CH/U_SLAVE_1ELK/Q[7]\ : DFN1C0
      port map(D => \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/Q[7]_net_1\);
    
    HIEFFPLA_INST_0_54944 : AND2A
      port map(A => HIEFFPLA_NET_0_117329, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_3[6]_net_1\, Y => 
        HIEFFPLA_NET_0_117163);
    
    HIEFFPLA_INST_0_49973 : MX2
      port map(A => HIEFFPLA_NET_0_118047, B => 
        HIEFFPLA_NET_0_118045, S => \BIT_OS_SEL_6[1]\, Y => 
        HIEFFPLA_NET_0_118035);
    
    \U_ELK12_CH/U_ELK1_SERDAT_SOURCE/SERDAT[6]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118547, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_2, Q => 
        \U_ELK12_CH/ELK_TX_DAT[6]\);
    
    \U50_PATTERNS/ELINK_ADDRA_6[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119961, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_4, Q => 
        \U50_PATTERNS/ELINK_ADDRA_6[6]\);
    
    HIEFFPLA_INST_0_63053 : AND3B
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[13]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[11]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[0]_net_1\, Y => 
        HIEFFPLA_NET_0_115903);
    
    \U50_PATTERNS/ELINK_DINA_16[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119808, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_18, Q => 
        \U50_PATTERNS/ELINK_DINA_16[7]\);
    
    \U50_PATTERNS/ELINK_DINA_9[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119718, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_19, Q => 
        \U50_PATTERNS/ELINK_DINA_9[1]\);
    
    \U_ELK16_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]\ : DFN1C0
      port map(D => \U_ELK16_CH/U_SLAVE_1ELK/Q[9]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]_net_1\);
    
    \U_ELK0_CMD_TX/SER_OUT_FI\ : DFI1C0
      port map(D => \U_ELK0_CMD_TX/SER_CMD_WORD_F[3]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_13, QN
         => \U_ELK0_CMD_TX/SER_OUT_FI_i\);
    
    HIEFFPLA_INST_0_38426 : MX2
      port map(A => \U50_PATTERNS/ELINKS_STRT_ADDR[7]\, B => 
        \U50_PATTERNS/ELINKS_STRT_ADDR_T[7]\, S => 
        HIEFFPLA_NET_0_119472, Y => HIEFFPLA_NET_0_120104);
    
    HIEFFPLA_INST_0_39542 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_4[4]\, B => 
        HIEFFPLA_NET_0_119519, S => HIEFFPLA_NET_0_119284, Y => 
        HIEFFPLA_NET_0_119979);
    
    \U50_PATTERNS/ELINK_ADDRA_5[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119969, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_3, Q => 
        \U50_PATTERNS/ELINK_ADDRA_5[6]\);
    
    \U_ELK19_CH/U_SLAVE_1ELK/Q[8]\ : DFN1C0
      port map(D => \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/Q[8]_net_1\);
    
    \P_USB_RXF_B_pad/U0/U1\ : IOIN_IRP
      port map(PRE => \AFLSDF_INV_0\, ICLK => CLK60MHZ, YIN => 
        \P_USB_RXF_B_pad/U0/NET1\, Y => \U50_PATTERNS/USB_RXF_B\);
    
    HIEFFPLA_INST_0_56021 : MX2
      port map(A => HIEFFPLA_NET_0_117013, B => 
        HIEFFPLA_NET_0_116037, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[2]\, Y => 
        HIEFFPLA_NET_0_116960);
    
    HIEFFPLA_INST_0_55213 : AND3B
      port map(A => HIEFFPLA_NET_0_117245, B => 
        HIEFFPLA_NET_0_117241, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[6]_net_1\, Y => 
        HIEFFPLA_NET_0_117088);
    
    \U_EXEC_MASTER/MPOR_SALT_B_0\ : DFI1P0
      port map(D => HIEFFPLA_NET_0_117781, CLK => CLK_40M_GL, PRE
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i\, QN => 
        MASTER_SALT_POR_B_i_0_i_0);
    
    HIEFFPLA_INST_0_53250 : XA1B
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[1]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[0]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[8]_net_1\, Y => 
        HIEFFPLA_NET_0_117446);
    
    HIEFFPLA_INST_0_61388 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_21[3]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_22[3]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_3[0]\, Y => 
        HIEFFPLA_NET_0_116133);
    
    \U50_PATTERNS/U4B_REGCROSS/LOCAL_REG_VAL[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119133, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_19, Q => \TFC_STOP_ADDR[0]\);
    
    HIEFFPLA_INST_0_57101 : AND2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_2[3]\, B => 
        HIEFFPLA_NET_0_116746, Y => HIEFFPLA_NET_0_116743);
    
    HIEFFPLA_INST_0_48082 : MX2
      port map(A => 
        \U_ELK16_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]_net_1\, B => 
        \U_ELK16_CH/ELK_TX_DAT[2]\, S => 
        \U_ELK16_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118381);
    
    \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117037, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_17_0, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[3]\);
    
    HIEFFPLA_INST_0_44584 : MX2
      port map(A => \ELKS_STOP_ADDR[4]\, B => 
        \U50_PATTERNS/U4D_REGCROSS/SAMP_TWO[4]_net_1\, S => 
        HIEFFPLA_NET_0_119093, Y => HIEFFPLA_NET_0_119087);
    
    HIEFFPLA_INST_0_53700 : AND3
      port map(A => HIEFFPLA_NET_0_117415, B => 
        HIEFFPLA_NET_0_116589, C => HIEFFPLA_NET_0_117361, Y => 
        HIEFFPLA_NET_0_117370);
    
    HIEFFPLA_INST_0_46830 : MX2
      port map(A => \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\, 
        B => \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[14]_net_1\, S => 
        \BIT_OS_SEL_7[2]\, Y => HIEFFPLA_NET_0_118608);
    
    \U50_PATTERNS/U4D_REGCROSS/SAMP_ONE[4]\ : DFN1C0
      port map(D => \U50_PATTERNS/ELINKS_STOP_ADDR[4]\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_25, Q => 
        \U50_PATTERNS/U4D_REGCROSS/SAMP_ONE[4]_net_1\);
    
    HIEFFPLA_INST_0_60001 : MX2
      port map(A => HIEFFPLA_NET_0_116815, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_4[3]\, S => 
        HIEFFPLA_NET_0_117202, Y => HIEFFPLA_NET_0_116323);
    
    HIEFFPLA_INST_0_39335 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_1[5]\, B => 
        HIEFFPLA_NET_0_119518, S => HIEFFPLA_NET_0_119243, Y => 
        HIEFFPLA_NET_0_120002);
    
    \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[1]\ : DFN1C0
      port map(D => 
        \U_ELK16_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\);
    
    \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[1]\ : DFN1C0
      port map(D => 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[1]_net_1\);
    
    HIEFFPLA_INST_0_40100 : AOI1D
      port map(A => HIEFFPLA_NET_0_119389, B => 
        HIEFFPLA_NET_0_119464, C => \U50_PATTERNS/SM_BANK_SEL[6]\, 
        Y => HIEFFPLA_NET_0_119906);
    
    \U_ELK15_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U1\ : IOBI_ID_OD_EB
      port map(DR => \U_ELK15_CH/ELK_OUT_R\, DF => 
        \U_ELK15_CH/ELK_OUT_F\, CLR => \GND\, E => 
        \AFLSDF_INV_24\, ICLK => CCC_160M_ADJ, OCLK => 
        CCC_160M_FXD, YIN => 
        \U_ELK15_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\, DOUT => 
        \U_ELK15_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, EOUT => 
        \U_ELK15_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET2\, YR => 
        \U_ELK15_CH/ELK_IN_DDR_R\, YF => 
        \U_ELK15_CH/ELK_IN_DDR_F\);
    
    HIEFFPLA_INST_0_55802 : MX2
      port map(A => HIEFFPLA_NET_0_116972, B => 
        HIEFFPLA_NET_0_117026, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[4]\, Y => 
        HIEFFPLA_NET_0_116988);
    
    HIEFFPLA_INST_0_62266 : AND2A
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[0]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_31[3]\, Y
         => HIEFFPLA_NET_0_116012);
    
    HIEFFPLA_INST_0_59394 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_26[1]\, B => 
        HIEFFPLA_NET_0_116742, S => HIEFFPLA_NET_0_117337, Y => 
        HIEFFPLA_NET_0_116397);
    
    HIEFFPLA_INST_0_55874 : MX2
      port map(A => HIEFFPLA_NET_0_116154, B => 
        HIEFFPLA_NET_0_116058, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[3]\, Y => 
        HIEFFPLA_NET_0_116979);
    
    HIEFFPLA_INST_0_57462 : AO1A
      port map(A => HIEFFPLA_NET_0_116678, B => 
        HIEFFPLA_NET_0_116742, C => HIEFFPLA_NET_0_116593, Y => 
        HIEFFPLA_NET_0_116677);
    
    HIEFFPLA_INST_0_44893 : AND3A
      port map(A => \U50_PATTERNS/REG_STATE_0[5]_net_1\, B => 
        HIEFFPLA_NET_0_119456, C => \U50_PATTERNS/USB_RXF_B\, Y
         => HIEFFPLA_NET_0_119026);
    
    HIEFFPLA_INST_0_58688 : AO1
      port map(A => HIEFFPLA_NET_0_116589, B => 
        HIEFFPLA_NET_0_117204, C => HIEFFPLA_NET_0_116483, Y => 
        HIEFFPLA_NET_0_116486);
    
    \U200A_TFC/RX_SER_WORD_2DEL[5]\ : DFN1C0
      port map(D => \U200A_TFC/RX_SER_WORD_1DEL[5]_net_1\, CLK
         => CLK_40M_GL, CLR => P_MASTER_POR_B_c, Q => 
        \U200A_TFC/RX_SER_WORD_2DEL[5]_net_1\);
    
    \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[5]\ : DFN1C0
      port map(D => 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\);
    
    HIEFFPLA_INST_0_48961 : MX2
      port map(A => \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\, 
        B => \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[12]_net_1\, S => 
        \BIT_OS_SEL_0[2]\, Y => HIEFFPLA_NET_0_118218);
    
    HIEFFPLA_INST_0_46603 : AND2
      port map(A => \U_ELK10_CH/ELK_TX_DAT[1]\, B => 
        \U_ELK10_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118648);
    
    HIEFFPLA_INST_0_37053 : AO1A
      port map(A => HIEFFPLA_NET_0_120338, B => 
        HIEFFPLA_NET_0_120325, C => HIEFFPLA_NET_0_120343, Y => 
        HIEFFPLA_NET_0_120357);
    
    \U_ELK0_CMD_TX/CLK40M_GEN_DEL0\ : DFN1C0
      port map(D => CLK_40M_GL, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_5, Q => 
        \U_ELK0_CMD_TX/CLK40M_GEN_DEL0_net_1\);
    
    \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[1]\ : DFN1C0
      port map(D => 
        \U_ELK4_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\);
    
    \U_ELK11_CH/U_ELK1_SERDAT_SOURCE/SERDAT[7]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118591, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_0, Q => 
        \U_ELK11_CH/ELK_TX_DAT[7]\);
    
    HIEFFPLA_INST_0_58367 : AND3A
      port map(A => HIEFFPLA_NET_0_117396, B => 
        HIEFFPLA_NET_0_116620, C => HIEFFPLA_NET_0_116649, Y => 
        HIEFFPLA_NET_0_116529);
    
    \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[13]\ : DFN1C0
      port map(D => 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[13]_net_1\);
    
    \U_ELK15_CH/U_ELK1_CMD_TX/SER_OUT_RDEL\ : DFN1C0
      port map(D => \U_ELK15_CH/U_ELK1_CMD_TX/SER_OUT_RI_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_5, Q
         => \U_ELK15_CH/ELK_OUT_R\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_8[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_115967, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_19, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_8[3]\);
    
    \U50_PATTERNS/REG_STATE[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119363, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_22_0, Q => 
        \U50_PATTERNS/REG_STATE[3]_net_1\);
    
    HIEFFPLA_INST_0_50262 : MX2
      port map(A => HIEFFPLA_NET_0_117997, B => 
        HIEFFPLA_NET_0_117996, S => \BIT_OS_SEL_0[0]\, Y => 
        \U_ELK5_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[4]\);
    
    HIEFFPLA_INST_0_43889 : MX2
      port map(A => HIEFFPLA_NET_0_119198, B => 
        \U50_PATTERNS/TFC_BLKA\, S => HIEFFPLA_NET_0_119294, Y
         => HIEFFPLA_NET_0_119199);
    
    HIEFFPLA_INST_0_43714 : NAND2B
      port map(A => \U50_PATTERNS/SM_BANK_SEL[5]\, B => 
        HIEFFPLA_NET_0_119242, Y => HIEFFPLA_NET_0_119234);
    
    HIEFFPLA_INST_0_63065 : AND2A
      port map(A => HIEFFPLA_NET_0_117078, B => 
        HIEFFPLA_NET_0_115896, Y => HIEFFPLA_NET_0_115897);
    
    \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[0]\ : DFN1C0
      port map(D => 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[0]_net_1\);
    
    HIEFFPLA_INST_0_44408 : MX2B
      port map(A => HIEFFPLA_NET_0_119124, B => 
        HIEFFPLA_NET_0_119135, S => 
        \U50_PATTERNS/U4B_REGCROSS/SYNC_SM[0]_net_1\, Y => 
        HIEFFPLA_NET_0_119125);
    
    \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[8]\ : DFN1C0
      port map(D => \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\);
    
    \U50_PATTERNS/USB_RD_BI/U1\ : DFN1P0
      port map(D => HIEFFPLA_NET_0_119036, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_13, Q => USB_RD_BI);
    
    HIEFFPLA_INST_0_41584 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_8[6]\, B => 
        HIEFFPLA_NET_0_119566, S => HIEFFPLA_NET_0_119291, Y => 
        HIEFFPLA_NET_0_119721);
    
    HIEFFPLA_INST_0_37774 : AO1A
      port map(A => HIEFFPLA_NET_0_120193, B => 
        HIEFFPLA_NET_0_120190, C => HIEFFPLA_NET_0_120210, Y => 
        HIEFFPLA_NET_0_120211);
    
    HIEFFPLA_INST_0_58543 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_16[1]\, B => 
        HIEFFPLA_NET_0_116677, S => HIEFFPLA_NET_0_117215, Y => 
        HIEFFPLA_NET_0_116507);
    
    \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[12]\ : DFN1C0
      port map(D => \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\, 
        CLK => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\);
    
    HIEFFPLA_INST_0_61352 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_21[0]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_22[0]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_3[0]\, Y => 
        HIEFFPLA_NET_0_116139);
    
    \U_ELK15_CH/U_ELK1_SERDAT_SOURCE/SERDAT[6]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118412, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_8, Q => 
        \U_ELK15_CH/ELK_TX_DAT[6]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_11[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116553, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_8, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_11[1]\);
    
    HIEFFPLA_INST_0_59492 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_11[3]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_27[3]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_5[4]_net_1\, Y
         => HIEFFPLA_NET_0_116387);
    
    HIEFFPLA_INST_0_52010 : AND2A
      port map(A => \U_MASTER_DES/U13A_ADJ_160M/BITCNT[0]\, B => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[50]\, Y => 
        HIEFFPLA_NET_0_117653);
    
    HIEFFPLA_INST_0_56922 : NAND3B
      port map(A => HIEFFPLA_NET_0_116771, B => 
        HIEFFPLA_NET_0_116772, C => HIEFFPLA_NET_0_116779, Y => 
        HIEFFPLA_NET_0_116774);
    
    HIEFFPLA_INST_0_43928 : MX2
      port map(A => HIEFFPLA_NET_0_119574, B => 
        \U50_PATTERNS/TFC_DINA[3]\, S => HIEFFPLA_NET_0_119294, Y
         => HIEFFPLA_NET_0_119194);
    
    \U_ELK8_CH/U_SLAVE_1ELK/Q[7]\ : DFN1C0
      port map(D => \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/Q[7]_net_1\);
    
    \U_ELK1_CH/U_SLAVE_1ELK/RECD_SER_WORD[6]\ : DFN1C0
      port map(D => \U_ELK1_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[6]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_1[6]\);
    
    HIEFFPLA_INST_0_37964 : MX2
      port map(A => \U200B_ELINKS/LOC_STOP_ADDR[5]\, B => 
        \ELKS_STOP_ADDR[5]\, S => 
        \U200B_ELINKS/GP_PG_SM_0[10]_net_1\, Y => 
        HIEFFPLA_NET_0_120182);
    
    \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[0]\ : DFN1C0
      port map(D => 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[0]_net_1\);
    
    HIEFFPLA_INST_0_48451 : MX2
      port map(A => \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\, 
        B => \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[12]_net_1\, S => 
        \BIT_OS_SEL_0[2]\, Y => HIEFFPLA_NET_0_118309);
    
    HIEFFPLA_INST_0_44629 : XO1
      port map(A => \U50_PATTERNS/U4D_REGCROSS/SAMP_TWO[2]_net_1\, 
        B => \ELKS_STOP_ADDR[2]\, C => HIEFFPLA_NET_0_119077, Y
         => HIEFFPLA_NET_0_119081);
    
    HIEFFPLA_INST_0_49634 : MX2
      port map(A => HIEFFPLA_NET_0_118088, B => 
        HIEFFPLA_NET_0_118085, S => \BIT_OS_SEL[1]\, Y => 
        HIEFFPLA_NET_0_118093);
    
    HIEFFPLA_INST_0_43009 : NOR3B
      port map(A => HIEFFPLA_NET_0_119430, B => 
        HIEFFPLA_NET_0_119016, C => HIEFFPLA_NET_0_119380, Y => 
        HIEFFPLA_NET_0_119404);
    
    \U_ELK5_CH/U_SLAVE_1ELK/Q[2]\ : DFN1C0
      port map(D => \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/Q[2]_net_1\);
    
    HIEFFPLA_INST_0_63007 : NAND3A
      port map(A => HIEFFPLA_NET_0_115907, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[8]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[7]\, Y => 
        HIEFFPLA_NET_0_115916);
    
    HIEFFPLA_INST_0_44118 : MX2
      port map(A => \U50_PATTERNS/TFC_STRT_ADDR[1]\, B => 
        \U50_PATTERNS/TFC_STRT_ADDR_T[1]\, S => 
        HIEFFPLA_NET_0_119472, Y => HIEFFPLA_NET_0_119171);
    
    HIEFFPLA_INST_0_55003 : OA1A
      port map(A => HIEFFPLA_NET_0_117240, B => 
        HIEFFPLA_NET_0_117247, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_3[6]_net_1\, Y => 
        HIEFFPLA_NET_0_117143);
    
    HIEFFPLA_INST_0_40095 : AOI1D
      port map(A => HIEFFPLA_NET_0_119389, B => 
        HIEFFPLA_NET_0_119464, C => \U50_PATTERNS/SM_BANK_SEL[7]\, 
        Y => HIEFFPLA_NET_0_119908);
    
    HIEFFPLA_INST_0_42647 : AND3B
      port map(A => HIEFFPLA_NET_0_119379, B => 
        \U50_PATTERNS/REG_STATE_0[2]_net_1\, C => 
        HIEFFPLA_NET_0_119400, Y => HIEFFPLA_NET_0_119492);
    
    \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[10]\ : DFN1C0
      port map(D => 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\);
    
    \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[5]\ : DFN1C0
      port map(D => 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\);
    
    HIEFFPLA_INST_0_44920 : NAND3B
      port map(A => \U50_PATTERNS/REG_STATE[4]_net_1\, B => 
        HIEFFPLA_NET_0_119449, C => 
        \U50_PATTERNS/REG_STATE[0]_net_1\, Y => 
        HIEFFPLA_NET_0_119019);
    
    \U_ELK14_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]\ : DFN1C0
      port map(D => \U_ELK14_CH/U_SLAVE_1ELK/Q[5]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]_net_1\);
    
    HIEFFPLA_INST_0_60393 : MX2
      port map(A => HIEFFPLA_NET_0_117075, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_10[3]\, S => 
        HIEFFPLA_NET_0_117154, Y => HIEFFPLA_NET_0_116272);
    
    HIEFFPLA_INST_0_48121 : AND2A
      port map(A => \OP_MODE_c_2[1]\, B => \PATT_ELK_DAT_16[4]\, 
        Y => HIEFFPLA_NET_0_118369);
    
    HIEFFPLA_INST_0_47375 : AND2A
      port map(A => \OP_MODE_c[1]\, B => \PATT_ELK_DAT_13[5]\, Y
         => HIEFFPLA_NET_0_118503);
    
    HIEFFPLA_INST_0_45807 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_12[1]\, C => 
        \U50_PATTERNS/SM_BANK_SEL[7]\, Y => HIEFFPLA_NET_0_118836);
    
    \U_ELK6_CH/U_ELK1_SERDAT_SOURCE/SERDAT[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117966, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_1, Q => 
        \U_ELK6_CH/ELK_TX_DAT[2]\);
    
    \U_ELK15_CH/U_SLAVE_1ELK/Q[0]\ : DFN1C0
      port map(D => \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/Q[0]_net_1\);
    
    HIEFFPLA_INST_0_53600 : MX2
      port map(A => HIEFFPLA_NET_0_117195, B => 
        HIEFFPLA_NET_0_117327, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[2]_net_1\, Y
         => HIEFFPLA_NET_0_117384);
    
    HIEFFPLA_INST_0_49449 : MX2
      port map(A => \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\, B
         => \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[11]_net_1\, S => 
        \BIT_OS_SEL_7[2]\, Y => HIEFFPLA_NET_0_118129);
    
    \U_ELK16_CH/U_SLAVE_1ELK/Q[6]\ : DFN1C0
      port map(D => \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/Q[6]_net_1\);
    
    HIEFFPLA_INST_0_56514 : AND3A
      port map(A => HIEFFPLA_NET_0_117430, B => \BIT_OS_SEL_1[2]\, 
        C => \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[6]_net_1\, 
        Y => HIEFFPLA_NET_0_116848);
    
    HIEFFPLA_INST_0_39695 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_6[5]\, B => 
        HIEFFPLA_NET_0_119518, S => HIEFFPLA_NET_0_119258, Y => 
        HIEFFPLA_NET_0_119962);
    
    HIEFFPLA_INST_0_57632 : NAND2A
      port map(A => HIEFFPLA_NET_0_116648, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_5[0]\, Y => 
        HIEFFPLA_NET_0_116647);
    
    HIEFFPLA_INST_0_39994 : MX2
      port map(A => HIEFFPLA_NET_0_119900, B => 
        \U50_PATTERNS/ELINK_BLKA[17]\, S => 
        \U50_PATTERNS/SM_BANK_SEL[20]\, Y => 
        HIEFFPLA_NET_0_119927);
    
    \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[7]\ : DFN1C0
      port map(D => 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\);
    
    \U_ELK15_CH/U_SLAVE_1ELK/Q[6]\ : DFN1C0
      port map(D => \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/Q[6]_net_1\);
    
    HIEFFPLA_INST_0_45438 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_18[7]\, C => 
        \U50_PATTERNS/SM_BANK_SEL[1]\, Y => HIEFFPLA_NET_0_118914);
    
    HIEFFPLA_INST_0_59332 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_26[1]\, B => 
        HIEFFPLA_NET_0_116401, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_2[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116405);
    
    \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_SEL_3[2]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_BIT_OS_VAL[2]\, CLK
         => CLK_40M_GL, CLR => P_MASTER_POR_B_c_27_1, Q => 
        \BIT_OS_SEL_3[2]\);
    
    HIEFFPLA_INST_0_57300 : AO1A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_3[3]\, B => 
        HIEFFPLA_NET_0_116714, C => HIEFFPLA_NET_0_117179, Y => 
        HIEFFPLA_NET_0_116704);
    
    HIEFFPLA_INST_0_50099 : MX2
      port map(A => 
        \U_ELK5_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]_net_1\, B => 
        \U_ELK5_CH/ELK_TX_DAT[5]\, S => 
        \U_ELK5_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118016);
    
    \U50_PATTERNS/U4A_REGCROSS/DELCNT[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119155, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_32, Q => 
        \U50_PATTERNS/U4A_REGCROSS/DELCNT[0]_net_1\);
    
    \U50_PATTERNS/ELINK_ADDRA_13[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120057, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_3, Q => 
        \U50_PATTERNS/ELINK_ADDRA_13[6]\);
    
    \U200B_ELINKS/LOC_STRT_ADDR[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120179, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_11, Q => 
        \U200B_ELINKS/LOC_STRT_ADDR[0]\);
    
    HIEFFPLA_INST_0_43239 : NAND3C
      port map(A => HIEFFPLA_NET_0_119358, B => 
        HIEFFPLA_NET_0_118995, C => HIEFFPLA_NET_0_119365, Y => 
        HIEFFPLA_NET_0_119341);
    
    \U200A_TFC/RX_SER_WORD_3DEL[1]\ : DFN1P0
      port map(D => \AFLSDF_INV_65\, CLK => CLK_40M_GL, PRE => 
        P_MASTER_POR_B_c_24, Q => 
        \U200A_TFC/RX_SER_WORD_3DEL_i_0[1]\);
    
    \U200A_TFC/LOC_STRT_ADDR[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120279, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_4, Q => \U200A_TFC/LOC_STRT_ADDR[3]\);
    
    HIEFFPLA_INST_0_42537 : OA1A
      port map(A => HIEFFPLA_NET_0_119433, B => 
        HIEFFPLA_NET_0_119010, C => \U50_PATTERNS/REG_ADDR[7]\, Y
         => HIEFFPLA_NET_0_119516);
    
    HIEFFPLA_INST_0_60098 : NAND3B
      port map(A => HIEFFPLA_NET_0_116304, B => 
        HIEFFPLA_NET_0_116305, C => HIEFFPLA_NET_0_116306, Y => 
        HIEFFPLA_NET_0_116310);
    
    HIEFFPLA_INST_0_54457 : AO1C
      port map(A => HIEFFPLA_NET_0_116589, B => 
        HIEFFPLA_NET_0_116620, C => HIEFFPLA_NET_0_117208, Y => 
        HIEFFPLA_NET_0_117263);
    
    \U200A_TFC/GP_PG_SM[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120319, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_28, Q => 
        \U200A_TFC/GP_PG_SM[2]_net_1\);
    
    HIEFFPLA_INST_0_49469 : MX2
      port map(A => HIEFFPLA_NET_0_118125, B => 
        HIEFFPLA_NET_0_118136, S => \BIT_OS_SEL[1]\, Y => 
        HIEFFPLA_NET_0_118126);
    
    HIEFFPLA_INST_0_38166 : MX2
      port map(A => \U50_PATTERNS/CHKSUM[2]\, B => 
        HIEFFPLA_NET_0_120133, S => HIEFFPLA_NET_0_119470, Y => 
        HIEFFPLA_NET_0_120141);
    
    \U_EXEC_MASTER/MPOR_SALT_B_11\ : DFI1P0
      port map(D => HIEFFPLA_NET_0_117781, CLK => CLK_40M_GL, PRE
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_2\, QN => 
        MASTER_SALT_POR_B_i_0_i_11);
    
    \U_ELK6_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U1\ : IOBI_ID_OD_EB
      port map(DR => \U_ELK6_CH/ELK_OUT_R\, DF => 
        \U_ELK6_CH/ELK_OUT_F\, CLR => \GND\, E => \AFLSDF_INV_44\, 
        ICLK => CCC_160M_ADJ, OCLK => CCC_160M_FXD, YIN => 
        \U_ELK6_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\, DOUT => 
        \U_ELK6_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, EOUT => 
        \U_ELK6_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET2\, YR => 
        \U_ELK6_CH/ELK_IN_DDR_R\, YF => \U_ELK6_CH/ELK_IN_DDR_F\);
    
    HIEFFPLA_INST_0_50377 : MX2
      port map(A => HIEFFPLA_NET_0_117955, B => 
        HIEFFPLA_NET_0_117953, S => \BIT_OS_SEL_5[1]\, Y => 
        HIEFFPLA_NET_0_117959);
    
    \U50_PATTERNS/U4B_REGCROSS/SAMP_ONE[4]\ : DFN1C0
      port map(D => \U50_PATTERNS/TFC_STOP_ADDR[4]\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_25, Q => 
        \U50_PATTERNS/U4B_REGCROSS/SAMP_ONE[4]_net_1\);
    
    \U_EXEC_MASTER/MPOR_B_27_0\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117787, CLK => CLK_40M_GL, CLR
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_0\, Q => 
        P_MASTER_POR_B_c_27_0);
    
    HIEFFPLA_INST_0_41071 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_1[5]\, B => 
        HIEFFPLA_NET_0_119567, S => HIEFFPLA_NET_0_119243, Y => 
        HIEFFPLA_NET_0_119778);
    
    \P_CLK_40M_GL_pad/U0/U0\ : IOPAD_TRI_U
      port map(D => \P_CLK_40M_GL_pad/U0/NET1\, E => 
        \P_CLK_40M_GL_pad/U0/NET2\, PAD => P_CLK_40M_GL);
    
    \U_ELK1_CH/U_SLAVE_1ELK/Q[11]\ : DFN1C0
      port map(D => \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/Q[11]_net_1\);
    
    HIEFFPLA_INST_0_42071 : AO1A
      port map(A => HIEFFPLA_NET_0_119622, B => 
        \U50_PATTERNS/TFC_STOP_ADDR[1]\, C => 
        HIEFFPLA_NET_0_118670, Y => HIEFFPLA_NET_0_119621);
    
    HIEFFPLA_INST_0_40909 : MX2
      port map(A => HIEFFPLA_NET_0_119574, B => 
        \U50_PATTERNS/ELINK_DINA_18[3]\, S => 
        HIEFFPLA_NET_0_119264, Y => HIEFFPLA_NET_0_119796);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_0[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116824, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_2, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_0[0]\);
    
    HIEFFPLA_INST_0_62221 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_31[0]\, B => 
        HIEFFPLA_NET_0_117190, S => HIEFFPLA_NET_0_117319, Y => 
        HIEFFPLA_NET_0_116020);
    
    HIEFFPLA_INST_0_46140 : AO1
      port map(A => HIEFFPLA_NET_0_119244, B => 
        \U50_PATTERNS/ELINK_DOUTA_2[5]\, C => 
        HIEFFPLA_NET_0_118932, Y => HIEFFPLA_NET_0_118757);
    
    \U_ELK6_CH/U_ELK1_CMD_TX/SER_OUT_FI\ : DFN1C0
      port map(D => 
        \U_ELK6_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_3, Q => 
        \U_ELK6_CH/U_ELK1_CMD_TX/SER_OUT_FI_net_1\);
    
    HIEFFPLA_INST_0_37097 : AND3B
      port map(A => \U200A_TFC/LOC_STRT_ADDR[0]\, B => 
        HIEFFPLA_NET_0_120293, C => HIEFFPLA_NET_0_120328, Y => 
        HIEFFPLA_NET_0_120348);
    
    \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[3]\ : DFN1C0
      port map(D => \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[6]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[4]_net_1\, CLK => 
        CCC_160M_ADJ, CLR => P_MASTER_POR_B_c_34_0, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[6]_net_1\);
    
    HIEFFPLA_INST_0_51856 : XA1
      port map(A => \U_MASTER_DES/U13A_ADJ_160M/BITCNT[6]\, B => 
        HIEFFPLA_NET_0_117690, C => HIEFFPLA_NET_0_117674, Y => 
        HIEFFPLA_NET_0_117676);
    
    \U_ELK1_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL\ : DFN1C0
      port map(D => 
        \U_ELK1_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL_net_1\);
    
    \U_ELK11_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]\ : DFN1C0
      port map(D => \U_ELK11_CH/U_SLAVE_1ELK/Q[3]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]_net_1\);
    
    HIEFFPLA_INST_0_52764 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_3[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_4[1]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[0]\, Y => 
        HIEFFPLA_NET_0_117515);
    
    HIEFFPLA_INST_0_46416 : NAND3C
      port map(A => \U50_PATTERNS/WR_XFER_TYPE[4]_net_1\, B => 
        \U50_PATTERNS/WR_XFER_TYPE[5]_net_1\, C => 
        \U50_PATTERNS/WR_XFER_TYPE[2]_net_1\, Y => 
        HIEFFPLA_NET_0_118695);
    
    HIEFFPLA_INST_0_43589 : AND2A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/SM_BANK_SEL[9]\, Y => HIEFFPLA_NET_0_119276);
    
    HIEFFPLA_INST_0_43222 : AO1A
      port map(A => HIEFFPLA_NET_0_119359, B => 
        HIEFFPLA_NET_0_119429, C => HIEFFPLA_NET_0_119343, Y => 
        HIEFFPLA_NET_0_119344);
    
    \U_ELK9_CH/ELK_IN_R\ : DFN1C0
      port map(D => \U_ELK9_CH/ELK_IN_DDR_R\, CLK => CCC_160M_ADJ, 
        CLR => DEV_RST_B_c, Q => \U_ELK9_CH/ELK_IN_R_net_1\);
    
    HIEFFPLA_INST_0_38885 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_14[3]\, B => 
        HIEFFPLA_NET_0_119520, S => HIEFFPLA_NET_0_119249, Y => 
        HIEFFPLA_NET_0_120052);
    
    \U_ELK18_CH/U_SLAVE_1ELK/Q[14]\ : DFN1C0
      port map(D => \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[14]_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/Q[14]_net_1\);
    
    HIEFFPLA_INST_0_40202 : AOI1D
      port map(A => HIEFFPLA_NET_0_119389, B => 
        HIEFFPLA_NET_0_119464, C => \U50_PATTERNS/SM_BANK_SEL[0]\, 
        Y => HIEFFPLA_NET_0_119874);
    
    \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[2]\ : DFN1C0
      port map(D => 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[2]_net_1\);
    
    \U50_PATTERNS/ELINK_DINA_18[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119796, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_21, Q => 
        \U50_PATTERNS/ELINK_DINA_18[3]\);
    
    HIEFFPLA_INST_0_56398 : NAND3C
      port map(A => HIEFFPLA_NET_0_116829, B => 
        HIEFFPLA_NET_0_116845, C => HIEFFPLA_NET_0_116853, Y => 
        HIEFFPLA_NET_0_116877);
    
    \U_ELK16_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]\ : DFN1C0
      port map(D => \U_ELK16_CH/U_SLAVE_1ELK/Q[11]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]_net_1\);
    
    \U_ELK8_CH/U_ELK1_SERDAT_SOURCE/SERDAT[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117877, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_5, Q => 
        \U_ELK8_CH/ELK_TX_DAT[1]\);
    
    HIEFFPLA_INST_0_61730 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_9[1]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_25[1]\, S
         => \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_3[4]_net_1\, 
        Y => HIEFFPLA_NET_0_116086);
    
    HIEFFPLA_INST_0_52806 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_7[0]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_8[0]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_2[0]\, Y => 
        HIEFFPLA_NET_0_117508);
    
    HIEFFPLA_INST_0_45563 : NAND3B
      port map(A => HIEFFPLA_NET_0_118781, B => 
        HIEFFPLA_NET_0_118787, C => HIEFFPLA_NET_0_119427, Y => 
        HIEFFPLA_NET_0_118889);
    
    \U_MASTER_DES/U13A_ADJ_160M/BITCNT[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117694, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_14, Q => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[4]\);
    
    \U200A_TFC/LOC_STRT_ADDR[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120278, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_4, Q => \U200A_TFC/LOC_STRT_ADDR[4]\);
    
    HIEFFPLA_INST_0_41134 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_2[4]\, B => 
        HIEFFPLA_NET_0_119570, S => HIEFFPLA_NET_0_119278, Y => 
        HIEFFPLA_NET_0_119771);
    
    HIEFFPLA_INST_0_55154 : AND3
      port map(A => HIEFFPLA_NET_0_117354, B => 
        HIEFFPLA_NET_0_117085, C => HIEFFPLA_NET_0_116813, Y => 
        HIEFFPLA_NET_0_117110);
    
    HIEFFPLA_INST_0_52654 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_17[0]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_18[0]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_3[0]\, Y => 
        HIEFFPLA_NET_0_117532);
    
    HIEFFPLA_INST_0_37423 : MX2
      port map(A => \U200A_TFC/LOC_STOP_ADDR[3]\, B => 
        \TFC_STOP_ADDR[3]\, S => \U200A_TFC/GP_PG_SM_0[10]_net_1\, 
        Y => HIEFFPLA_NET_0_120287);
    
    HIEFFPLA_INST_0_60486 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_11[0]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_12[0]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_4[0]\, Y => 
        HIEFFPLA_NET_0_116260);
    
    HIEFFPLA_INST_0_37306 : AND3
      port map(A => \U200A_TFC/GP_PG_SM[4]_net_1\, B => 
        HIEFFPLA_NET_0_120326, C => HIEFFPLA_NET_0_120293, Y => 
        HIEFFPLA_NET_0_120298);
    
    \U50_PATTERNS/U4E_REGCROSS/SAMP_TWO[3]\ : DFN1C0
      port map(D => \U50_PATTERNS/U4E_REGCROSS/SAMP_ONE[3]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_23, Q => 
        \U50_PATTERNS/U4E_REGCROSS/SAMP_TWO[3]_net_1\);
    
    HIEFFPLA_INST_0_59744 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_30[2]\, B => 
        HIEFFPLA_NET_0_116348, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_1[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116354);
    
    \U_ELK4_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118066, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_1, Q => 
        \U_ELK4_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]_net_1\);
    
    HIEFFPLA_INST_0_41977 : AND3C
      port map(A => HIEFFPLA_NET_0_119238, B => 
        HIEFFPLA_NET_0_119270, C => 
        \U50_PATTERNS/SM_BANK_SEL[13]\, Y => 
        HIEFFPLA_NET_0_119640);
    
    HIEFFPLA_INST_0_62382 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_4[4]\, 
        B => HIEFFPLA_NET_0_117100, S => HIEFFPLA_NET_0_117148, Y
         => HIEFFPLA_NET_0_115996);
    
    HIEFFPLA_INST_0_56783 : XA1B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_0[2]\, B => 
        HIEFFPLA_NET_0_116791, C => HIEFFPLA_NET_0_117085, Y => 
        HIEFFPLA_NET_0_116798);
    
    HIEFFPLA_INST_0_52818 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_7[2]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_8[2]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_2[0]\, Y => 
        HIEFFPLA_NET_0_117506);
    
    HIEFFPLA_INST_0_45244 : NAND2B
      port map(A => HIEFFPLA_NET_0_118734, B => 
        HIEFFPLA_NET_0_118746, Y => HIEFFPLA_NET_0_118959);
    
    HIEFFPLA_INST_0_60366 : MX2
      port map(A => HIEFFPLA_NET_0_117096, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_10[0]\, S => 
        HIEFFPLA_NET_0_117154, Y => HIEFFPLA_NET_0_116275);
    
    HIEFFPLA_INST_0_60804 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_15[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_16[1]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[0]\, Y => 
        HIEFFPLA_NET_0_116217);
    
    \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[13]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[11]_net_1\, CLK => 
        CCC_160M_ADJ, CLR => P_MASTER_POR_B_c_26, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[13]_net_1\);
    
    HIEFFPLA_INST_0_57155 : XA1B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_2[6]\, B => 
        HIEFFPLA_NET_0_116744, C => HIEFFPLA_NET_0_117179, Y => 
        HIEFFPLA_NET_0_116729);
    
    HIEFFPLA_INST_0_56259 : AND2B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/RECD_SER_WORD[6]_net_1\, 
        B => 
        \U_MASTER_DES/U13C_MASTER_DESER/RECD_SER_WORD[5]_net_1\, 
        Y => HIEFFPLA_NET_0_116905);
    
    HIEFFPLA_INST_0_51473 : MX2
      port map(A => HIEFFPLA_NET_0_117761, B => 
        \U_EXEC_MASTER/PRESCALE[1]\, S => HIEFFPLA_NET_0_117787, 
        Y => HIEFFPLA_NET_0_117767);
    
    \U50_PATTERNS/ELINK_ADDRA_12[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120067, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_2_0, Q => 
        \U50_PATTERNS/ELINK_ADDRA_12[4]\);
    
    HIEFFPLA_INST_0_50360 : NAND2B
      port map(A => \OP_MODE_c_0[1]\, B => \PATT_ELK_DAT_6[2]\, Y
         => HIEFFPLA_NET_0_117966);
    
    HIEFFPLA_INST_0_49680 : MX2
      port map(A => HIEFFPLA_NET_0_118091, B => 
        HIEFFPLA_NET_0_118088, S => \BIT_OS_SEL[1]\, Y => 
        HIEFFPLA_NET_0_118086);
    
    HIEFFPLA_INST_0_40288 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_0[6]\, B => 
        HIEFFPLA_NET_0_119566, S => HIEFFPLA_NET_0_119272, Y => 
        HIEFFPLA_NET_0_119865);
    
    HIEFFPLA_INST_0_54125 : MX2
      port map(A => HIEFFPLA_NET_0_116360, B => 
        HIEFFPLA_NET_0_116558, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_1[3]_net_1\, Y
         => HIEFFPLA_NET_0_117305);
    
    HIEFFPLA_INST_0_51401 : NAND2
      port map(A => \U_EXEC_MASTER/DEL_CNT[0]\, B => 
        \U_EXEC_MASTER/DEL_CNT[1]\, Y => HIEFFPLA_NET_0_117786);
    
    HIEFFPLA_INST_0_37262 : AND3
      port map(A => HIEFFPLA_NET_0_120327, B => 
        HIEFFPLA_NET_0_120303, C => HIEFFPLA_NET_0_120333, Y => 
        HIEFFPLA_NET_0_120311);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_10[4]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116271, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_18, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_10[4]\);
    
    HIEFFPLA_INST_0_43115 : NAND2
      port map(A => \U50_PATTERNS/REG_STATE[2]_net_1\, B => 
        \U50_PATTERNS/REG_STATE[0]_net_1\, Y => 
        HIEFFPLA_NET_0_119372);
    
    \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[1]\ : DFN1C0
      port map(D => 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[1]_net_1\);
    
    \U50_PATTERNS/U4E_REGCROSS/LOCAL_REG_VAL[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119063, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_6, Q => 
        \U50_PATTERNS/U4E_REGCROSS/LOCAL_REG_VAL[7]\);
    
    \U_ELK18_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]\ : DFN1C0
      port map(D => \U_ELK18_CH/U_SLAVE_1ELK/Q[3]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]_net_1\);
    
    HIEFFPLA_INST_0_42749 : AND3C
      port map(A => HIEFFPLA_NET_0_119017, B => 
        \U50_PATTERNS/REG_STATE_0[1]_net_1\, C => 
        \U50_PATTERNS/REG_STATE_0[2]_net_1\, Y => 
        HIEFFPLA_NET_0_119469);
    
    HIEFFPLA_INST_0_49491 : MX2
      port map(A => HIEFFPLA_NET_0_118126, B => 
        HIEFFPLA_NET_0_118137, S => \BIT_OS_SEL_1[0]\, Y => 
        \U_ELK2_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[1]\);
    
    \U_ELK15_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]\ : DFN1C0
      port map(D => \U_ELK15_CH/U_SLAVE_1ELK/Q[7]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]_net_1\);
    
    HIEFFPLA_INST_0_51779 : MX2
      port map(A => \U_MASTER_DES/U13A_ADJ_160M/BITCNT[5]\, B => 
        HIEFFPLA_NET_0_117677, S => HIEFFPLA_NET_0_117630, Y => 
        HIEFFPLA_NET_0_117693);
    
    HIEFFPLA_INST_0_50439 : MX2
      port map(A => HIEFFPLA_NET_0_117952, B => 
        HIEFFPLA_NET_0_117948, S => \BIT_OS_SEL_5[1]\, Y => 
        HIEFFPLA_NET_0_117950);
    
    \U50_PATTERNS/TFC_STOP_ADDR_T[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119173, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_15, Q => 
        \U50_PATTERNS/TFC_STOP_ADDR_T[7]\);
    
    HIEFFPLA_INST_0_57509 : XA1B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_4[5]\, B => 
        HIEFFPLA_NET_0_116684, C => HIEFFPLA_NET_0_117179, Y => 
        HIEFFPLA_NET_0_116666);
    
    HIEFFPLA_INST_0_41730 : MX2
      port map(A => HIEFFPLA_NET_0_119682, B => 
        \U50_PATTERNS/ELINK_RWA[17]\, S => 
        \U50_PATTERNS/SM_BANK_SEL_0[20]\, Y => 
        HIEFFPLA_NET_0_119703);
    
    HIEFFPLA_INST_0_48075 : MX2
      port map(A => \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\, 
        B => \U_ELK15_CH/U_SLAVE_1ELK/ARB_BYTE[14]_net_1\, S => 
        \BIT_OS_SEL_4[2]\, Y => HIEFFPLA_NET_0_118383);
    
    \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[3]\ : DFN1C0
      port map(D => \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\);
    
    HIEFFPLA_INST_0_50357 : AND2
      port map(A => CLK_40M_GL, B => 
        \U_ELK6_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0_net_1\, Y => 
        HIEFFPLA_NET_0_117969);
    
    HIEFFPLA_INST_0_42046 : AND3
      port map(A => \U50_PATTERNS/TFC_DOUTA[5]\, B => 
        HIEFFPLA_NET_0_118997, C => HIEFFPLA_NET_0_119365, Y => 
        HIEFFPLA_NET_0_119624);
    
    \U200A_TFC/LOC_STOP_ADDR[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120284, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_1, Q => \U200A_TFC/LOC_STOP_ADDR[6]\);
    
    HIEFFPLA_INST_0_59764 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_14[3]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_30[3]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_3[4]_net_1\, Y
         => HIEFFPLA_NET_0_116351);
    
    \U_TFC_CMD_TX/SER_CMD_WORD_R[2]\ : DFN1C0
      port map(D => \U_TFC_CMD_TX/N_SER_CMD_WORD_R[2]\, CLK => 
        CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_TFC_CMD_TX/SER_CMD_WORD_R[2]_net_1\);
    
    HIEFFPLA_INST_0_53150 : MX2
      port map(A => HIEFFPLA_NET_0_117539, B => 
        HIEFFPLA_NET_0_117535, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_1[3]\, Y => 
        HIEFFPLA_NET_0_117459);
    
    HIEFFPLA_INST_0_49862 : NAND2B
      port map(A => \OP_MODE_c_1[1]\, B => \PATT_ELK_DAT_4[2]\, Y
         => HIEFFPLA_NET_0_118056);
    
    HIEFFPLA_INST_0_60947 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_17[3]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_18[3]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_4[0]\, Y => 
        HIEFFPLA_NET_0_116194);
    
    HIEFFPLA_INST_0_38035 : AOI1A
      port map(A => HIEFFPLA_NET_0_120232, B => 
        HIEFFPLA_NET_0_120220, C => HIEFFPLA_NET_0_120168, Y => 
        HIEFFPLA_NET_0_120169);
    
    \U50_PATTERNS/ELINK_ADDRA_3[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119986, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_1, Q => 
        \U50_PATTERNS/ELINK_ADDRA_3[5]\);
    
    \U200A_TFC/LOC_STOP_ADDR[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120285, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_1, Q => \U200A_TFC/LOC_STOP_ADDR[5]\);
    
    HIEFFPLA_INST_0_37940 : MX2
      port map(A => \U200B_ELINKS/LOC_STOP_ADDR[1]\, B => 
        \ELKS_STOP_ADDR[1]\, S => 
        \U200B_ELINKS/GP_PG_SM_0[10]_net_1\, Y => 
        HIEFFPLA_NET_0_120186);
    
    \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[10]\ : DFN1C0
      port map(D => 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]_net_1\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\);
    
    HIEFFPLA_INST_0_52462 : MX2
      port map(A => HIEFFPLA_NET_0_117508, B => 
        HIEFFPLA_NET_0_117504, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[3]\, Y => 
        HIEFFPLA_NET_0_117560);
    
    HIEFFPLA_INST_0_111347 : NAND3C
      port map(A => HIEFFPLA_NET_0_116806, B => 
        HIEFFPLA_NET_0_116742, C => HIEFFPLA_NET_0_116687, Y => 
        HIEFFPLA_NET_0_115841);
    
    HIEFFPLA_INST_0_60852 : MX2
      port map(A => HIEFFPLA_NET_0_117166, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_16[4]\, S => 
        HIEFFPLA_NET_0_117142, Y => HIEFFPLA_NET_0_116211);
    
    HIEFFPLA_INST_0_48200 : MX2
      port map(A => HIEFFPLA_NET_0_118358, B => 
        HIEFFPLA_NET_0_118355, S => \BIT_OS_SEL_2[1]\, Y => 
        HIEFFPLA_NET_0_118354);
    
    \U_ELK12_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]\ : DFN1C0
      port map(D => \U_ELK12_CH/U_SLAVE_1ELK/Q[7]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]_net_1\);
    
    HIEFFPLA_INST_0_57827 : AO1A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_6[3]\, B => 
        HIEFFPLA_NET_0_116623, C => HIEFFPLA_NET_0_117179, Y => 
        HIEFFPLA_NET_0_116612);
    
    HIEFFPLA_INST_0_61310 : MX2
      port map(A => HIEFFPLA_NET_0_117167, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_21[1]\, S => 
        HIEFFPLA_NET_0_117144, Y => HIEFFPLA_NET_0_116144);
    
    \U50_PATTERNS/ELINK_DINA_19[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119790, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_0, Q => 
        \U50_PATTERNS/ELINK_DINA_19[1]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_6[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116314, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_2, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_6[0]\);
    
    \U_ELK8_CH/U_SLAVE_1ELK/Q[12]\ : DFN1C0
      port map(D => \U_ELK8_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/Q[12]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_5[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116658, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_11, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_5[3]\);
    
    \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[12]\ : DFN1C0
      port map(D => \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\);
    
    HIEFFPLA_INST_0_60786 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_31[3]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_15[3]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[4]_net_1\, Y
         => HIEFFPLA_NET_0_116220);
    
    HIEFFPLA_INST_0_43626 : AND2B
      port map(A => \U50_PATTERNS/SM_BANK_SEL[21]\, B => 
        \U50_PATTERNS/SM_BANK_SEL[1]\, Y => HIEFFPLA_NET_0_119264);
    
    HIEFFPLA_INST_0_41287 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_4[5]\, B => 
        HIEFFPLA_NET_0_119567, S => HIEFFPLA_NET_0_119284, Y => 
        HIEFFPLA_NET_0_119754);
    
    HIEFFPLA_INST_0_58079 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_0[0]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_16[0]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_1[4]_net_1\, Y
         => HIEFFPLA_NET_0_116567);
    
    HIEFFPLA_INST_0_54472 : MX2
      port map(A => HIEFFPLA_NET_0_117271, B => 
        HIEFFPLA_NET_0_117288, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[2]_net_1\, Y => 
        HIEFFPLA_NET_0_117261);
    
    HIEFFPLA_INST_0_42424 : AND2
      port map(A => HIEFFPLA_NET_0_119473, B => 
        \U50_PATTERNS/RD_XFER_TYPE[2]_net_1\, Y => 
        HIEFFPLA_NET_0_119539);
    
    HIEFFPLA_INST_0_49001 : MX2
      port map(A => HIEFFPLA_NET_0_118228, B => 
        HIEFFPLA_NET_0_118227, S => \BIT_OS_SEL_2[0]\, Y => 
        \U_ELK19_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[2]\);
    
    \U_ELK2_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2\ : IOPADN_BI
      port map(DB => \U_ELK2_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, 
        E => \U_ELK2_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET3\, PAD => 
        ELK2_DAT_N, N2POUT => 
        \U_ELK2_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2_N2P\);
    
    \U50_PATTERNS/TFC_STOP_ADDR[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119184, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_8, Q => 
        \U50_PATTERNS/TFC_STOP_ADDR[4]\);
    
    HIEFFPLA_INST_0_59364 : MX2A
      port map(A => HIEFFPLA_NET_0_117397, B => 
        HIEFFPLA_NET_0_116397, S => HIEFFPLA_NET_0_117404, Y => 
        HIEFFPLA_NET_0_116401);
    
    HIEFFPLA_INST_0_44915 : AND2A
      port map(A => \U50_PATTERNS/USB_RXF_B\, B => 
        \U50_PATTERNS/REG_STATE[2]_net_1\, Y => 
        HIEFFPLA_NET_0_119021);
    
    \U_ELK8_CH/U_ELK1_SERDAT_SOURCE/SERDAT[4]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117874, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_5, Q => 
        \U_ELK8_CH/ELK_TX_DAT[4]\);
    
    \U_ELK15_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]\ : DFN1C0
      port map(D => \U_ELK15_CH/U_SLAVE_1ELK/Q[3]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]_net_1\);
    
    HIEFFPLA_INST_0_61877 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_27[4]\, B => 
        HIEFFPLA_NET_0_117100, S => HIEFFPLA_NET_0_117196, Y => 
        HIEFFPLA_NET_0_116066);
    
    HIEFFPLA_INST_0_60929 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_17[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_18[1]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_4[0]\, Y => 
        HIEFFPLA_NET_0_116197);
    
    HIEFFPLA_INST_0_46517 : AOI1C
      port map(A => HIEFFPLA_NET_0_119596, B => 
        HIEFFPLA_NET_0_119571, C => 
        \U50_PATTERNS/WR_XFER_TYPE[2]_net_1\, Y => 
        HIEFFPLA_NET_0_118674);
    
    HIEFFPLA_INST_0_39029 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_16[3]\, B => 
        HIEFFPLA_NET_0_119520, S => HIEFFPLA_NET_0_119257, Y => 
        HIEFFPLA_NET_0_120036);
    
    \U_ELK6_CH/U_SLAVE_1ELK/RECD_SER_WORD[2]\ : DFN1C0
      port map(D => \U_ELK6_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[2]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_6[2]\);
    
    \U_ELK2_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U3\ : IOBI_ID_OD_EB
      port map(DR => \U_ELK2_CH/ELK_OUT_R\, DF => 
        \U_ELK2_CH/ELK_OUT_F\, CLR => \GND\, E => \AFLSDF_INV_37\, 
        ICLK => CCC_160M_ADJ, OCLK => CCC_160M_FXD, YIN => 
        \U_ELK2_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\, DOUT => OPEN, 
        EOUT => \U_ELK2_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET3\, YR
         => OPEN, YF => OPEN);
    
    HIEFFPLA_INST_0_37515 : NAND2B
      port map(A => \U200A_TFC/RX_SER_WORD_3DEL_i_0[7]\, B => 
        \U200A_TFC/RX_SER_WORD_3DEL[6]_net_1\, Y => 
        HIEFFPLA_NET_0_120270);
    
    \U_ELK7_CH/U_ELK1_CMD_TX/SER_OUT_FI\ : DFN1C0
      port map(D => 
        \U_ELK7_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_13, Q
         => \U_ELK7_CH/U_ELK1_CMD_TX/SER_OUT_FI_net_1\);
    
    \U50_PATTERNS/ELINK_ADDRA_5[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119970, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_3, Q => 
        \U50_PATTERNS/ELINK_ADDRA_5[5]\);
    
    HIEFFPLA_INST_0_59228 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_25[2]\, B => 
        HIEFFPLA_NET_0_116414, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_2[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116418);
    
    HIEFFPLA_INST_0_47250 : MX2
      port map(A => HIEFFPLA_NET_0_118540, B => 
        HIEFFPLA_NET_0_118538, S => \BIT_OS_SEL_5[0]\, Y => 
        \U_ELK12_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[1]\);
    
    HIEFFPLA_INST_0_58318 : AO1B
      port map(A => HIEFFPLA_NET_0_117396, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_13[2]\, C => 
        HIEFFPLA_NET_0_117367, Y => HIEFFPLA_NET_0_116535);
    
    \U_ELK5_CH/U_SLAVE_1ELK/RECD_SER_WORD[5]\ : DFN1C0
      port map(D => \U_ELK5_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[5]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_5[5]\);
    
    HIEFFPLA_INST_0_58200 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_11[3]\, B => 
        HIEFFPLA_NET_0_116549, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_0[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116551);
    
    HIEFFPLA_INST_0_61130 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_1[1]\, 
        B => HIEFFPLA_NET_0_117167, S => HIEFFPLA_NET_0_117149, Y
         => HIEFFPLA_NET_0_116169);
    
    HIEFFPLA_INST_0_58981 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_5[3]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_21[3]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_5[4]_net_1\, Y
         => HIEFFPLA_NET_0_116451);
    
    HIEFFPLA_INST_0_42512 : MX2
      port map(A => \U50_PATTERNS/REG_ADDR[8]\, B => 
        HIEFFPLA_NET_0_119501, S => HIEFFPLA_NET_0_119007, Y => 
        HIEFFPLA_NET_0_119525);
    
    HIEFFPLA_INST_0_54598 : AND3B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[4]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[2]_net_1\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[1]_net_1\, Y => 
        HIEFFPLA_NET_0_117235);
    
    HIEFFPLA_INST_0_49250 : MX2
      port map(A => HIEFFPLA_NET_0_118185, B => 
        HIEFFPLA_NET_0_118183, S => \BIT_OS_SEL_2[0]\, Y => 
        \U_ELK1_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[2]\);
    
    \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[8]\ : DFN1C0
      port map(D => \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\);
    
    \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[2]\ : DFN1C0
      port map(D => 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_BYTE[2]_net_1\);
    
    HIEFFPLA_INST_0_56477 : AO1
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[5]_net_1\, B => 
        HIEFFPLA_NET_0_117428, C => HIEFFPLA_NET_0_116839, Y => 
        HIEFFPLA_NET_0_116855);
    
    HIEFFPLA_INST_0_37029 : AO1A
      port map(A => \TFC_STRT_ADDR[1]\, B => 
        HIEFFPLA_NET_0_120349, C => HIEFFPLA_NET_0_120347, Y => 
        HIEFFPLA_NET_0_120365);
    
    HIEFFPLA_INST_0_57855 : AOI1
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_6[0]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_6[1]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_6[2]\, Y => 
        HIEFFPLA_NET_0_116606);
    
    HIEFFPLA_INST_0_46115 : AO1
      port map(A => HIEFFPLA_NET_0_119276, B => 
        \U50_PATTERNS/ELINK_DOUTA_10[0]\, C => 
        HIEFFPLA_NET_0_118937, Y => HIEFFPLA_NET_0_118762);
    
    AFLSDF_INV_52 : INV
      port map(A => CLK_40M_GL, Y => \AFLSDF_INV_52\);
    
    HIEFFPLA_INST_0_63214 : MX2
      port map(A => \U_TFC_CMD_TX/SER_CMD_WORD_F[2]_net_1\, B => 
        \TFC_TX_DAT[6]\, S => \U_TFC_CMD_TX/START_RISE_net_1\, Y
         => \U_TFC_CMD_TX/N_SER_CMD_WORD_F[3]\);
    
    HIEFFPLA_INST_0_37517 : NAND3C
      port map(A => HIEFFPLA_NET_0_120270, B => 
        \U200A_TFC/RX_SER_WORD_3DEL[4]_net_1\, C => 
        \U200A_TFC/RX_SER_WORD_3DEL[5]_net_1\, Y => 
        HIEFFPLA_NET_0_120269);
    
    \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[3]\ : DFN1C0
      port map(D => 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[3]_net_1\);
    
    HIEFFPLA_INST_0_49112 : AND2
      port map(A => CLK_40M_GL, B => 
        \U_ELK1_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0_net_1\, Y => 
        HIEFFPLA_NET_0_118194);
    
    \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[14]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[12]_net_1\, CLK => 
        CCC_160M_ADJ, CLR => P_MASTER_POR_B_c_26, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[14]_net_1\);
    
    HIEFFPLA_INST_0_46071 : AND3A
      port map(A => HIEFFPLA_NET_0_119376, B => 
        \U50_PATTERNS/TFC_STRT_ADDR[0]\, C => 
        HIEFFPLA_NET_0_119431, Y => HIEFFPLA_NET_0_118773);
    
    HIEFFPLA_INST_0_44198 : MX2
      port map(A => \U50_PATTERNS/TFC_STRT_ADDR_T[3]\, B => 
        \U50_PATTERNS/RD_USB_ADBUS[3]\, S => 
        HIEFFPLA_NET_0_119491, Y => HIEFFPLA_NET_0_119161);
    
    HIEFFPLA_INST_0_56725 : NAND3C
      port map(A => HIEFFPLA_NET_0_116773, B => 
        HIEFFPLA_NET_0_117343, C => HIEFFPLA_NET_0_116803, Y => 
        HIEFFPLA_NET_0_116814);
    
    \U50_PATTERNS/TFC_STOP_ADDR[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119186, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_8, Q => 
        \U50_PATTERNS/TFC_STOP_ADDR[2]\);
    
    HIEFFPLA_INST_0_113943 : AO18
      port map(A => HIEFFPLA_NET_0_115821, B => \ELKS_ADDRB[4]\, 
        C => \U200B_ELINKS/LOC_STOP_ADDR[4]\, Y => 
        HIEFFPLA_NET_0_115808);
    
    HIEFFPLA_INST_0_37781 : NOR3B
      port map(A => HIEFFPLA_NET_0_120158, B => 
        HIEFFPLA_NET_0_120160, C => HIEFFPLA_NET_0_120208, Y => 
        HIEFFPLA_NET_0_120209);
    
    HIEFFPLA_INST_0_48642 : MX2
      port map(A => \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[1]_net_1\, 
        B => \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\, S => 
        \BIT_OS_SEL_0[2]\, Y => HIEFFPLA_NET_0_118273);
    
    AFLSDF_INV_15 : INV
      port map(A => DCB_SALT_SEL_c, Y => \AFLSDF_INV_15\);
    
    \U50_PATTERNS/U4D_REGCROSS/LOCAL_REG_VAL[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119089, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_3, Q => \ELKS_STOP_ADDR[2]\);
    
    HIEFFPLA_INST_0_161268 : DFN1C0
      port map(D => \U_ELK1_CH/U_ELK1_CMD_TX/START_RISE_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_4, Q
         => HIEFFPLA_NET_0_161287);
    
    \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[4]\ : DFN1C0
      port map(D => \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\);
    
    \U_ELK10_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]\ : DFN1C0
      port map(D => \U_ELK10_CH/U_SLAVE_1ELK/Q[7]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]_net_1\);
    
    HIEFFPLA_INST_0_61940 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_27[4]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_28[4]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[0]\, Y => 
        HIEFFPLA_NET_0_116056);
    
    HIEFFPLA_INST_0_46760 : MX2
      port map(A => HIEFFPLA_NET_0_118629, B => 
        HIEFFPLA_NET_0_118625, S => \BIT_OS_SEL_0[0]\, Y => 
        \U_ELK10_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[2]\);
    
    HIEFFPLA_INST_0_57589 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_5[6]\, B => 
        HIEFFPLA_NET_0_116638, S => HIEFFPLA_NET_0_117121, Y => 
        HIEFFPLA_NET_0_116655);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_11[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116263, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_20, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_11[2]\);
    
    \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[11]\ : DFN1C0
      port map(D => \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\);
    
    HIEFFPLA_INST_0_60570 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_13[1]\, B => 
        HIEFFPLA_NET_0_117167, S => HIEFFPLA_NET_0_117137, Y => 
        HIEFFPLA_NET_0_116249);
    
    \U50_PATTERNS/ELINK_DINA_8[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119721, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_18, Q => 
        \U50_PATTERNS/ELINK_DINA_8[6]\);
    
    HIEFFPLA_INST_0_57250 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_3[8]\, B => 
        HIEFFPLA_NET_0_116699, S => HIEFFPLA_NET_0_117120, Y => 
        HIEFFPLA_NET_0_116717);
    
    HIEFFPLA_INST_0_39569 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_4[7]\, B => 
        HIEFFPLA_NET_0_119516, S => HIEFFPLA_NET_0_119284, Y => 
        HIEFFPLA_NET_0_119976);
    
    HIEFFPLA_INST_0_44325 : XO1
      port map(A => \TFC_STRT_ADDR[5]\, B => 
        \U50_PATTERNS/U4A_REGCROSS/SAMP_TWO[5]_net_1\, C => 
        HIEFFPLA_NET_0_119141, Y => HIEFFPLA_NET_0_119142);
    
    \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_115937, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_24_0, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[3]_net_1\);
    
    \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[4]\ : DFN1C0
      port map(D => \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\);
    
    \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[5]\ : DFN1C0
      port map(D => \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\);
    
    HIEFFPLA_INST_0_49084 : MX2
      port map(A => 
        \U_ELK1_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]_net_1\, B => 
        \U_ELK1_CH/ELK_TX_DAT[4]\, S => 
        \U_ELK1_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118200);
    
    HIEFFPLA_INST_0_60860 : AND2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[4]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_16[2]\, Y => 
        HIEFFPLA_NET_0_116208);
    
    HIEFFPLA_INST_0_40103 : AOI1A
      port map(A => \U50_PATTERNS/ELINK_BLKA[14]\, B => 
        HIEFFPLA_NET_0_119235, C => HIEFFPLA_NET_0_119877, Y => 
        HIEFFPLA_NET_0_119905);
    
    HIEFFPLA_INST_0_37396 : MX2
      port map(A => \U200A_TFC/N_232_li\, B => DCB_SALT_SEL_c, S
         => \U200A_TFC/GP_PG_SM[10]_net_1\, Y => 
        HIEFFPLA_NET_0_120292);
    
    HIEFFPLA_INST_0_59669 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_2[3]\, B => 
        HIEFFPLA_NET_0_116358, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_1[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116364);
    
    HIEFFPLA_INST_0_40891 : MX2
      port map(A => HIEFFPLA_NET_0_119576, B => 
        \U50_PATTERNS/ELINK_DINA_18[1]\, S => 
        HIEFFPLA_NET_0_119264, Y => HIEFFPLA_NET_0_119798);
    
    \U_ELK3_CH/ELK_IN_F\ : DFN1C0
      port map(D => \AFLSDF_INV_66\, CLK => CCC_160M_ADJ, CLR => 
        DEV_RST_B_c, Q => \U_ELK3_CH/ELK_IN_F_net_1\);
    
    \U_ELK13_CH/U_SLAVE_1ELK/RECD_SER_WORD[3]\ : DFN1C0
      port map(D => \U_ELK13_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[3]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_13[3]\);
    
    \U_ELK13_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]\ : DFN1C0
      port map(D => \U_ELK13_CH/U_SLAVE_1ELK/Q[7]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]_net_1\);
    
    HIEFFPLA_INST_0_59177 : AOI1D
      port map(A => HIEFFPLA_NET_0_116345, B => 
        HIEFFPLA_NET_0_116740, C => HIEFFPLA_NET_0_117208, Y => 
        HIEFFPLA_NET_0_116424);
    
    \U50_PATTERNS/U4A_REGCROSS/SAMP_TWO[4]\ : DFN1C0
      port map(D => \U50_PATTERNS/U4A_REGCROSS/SAMP_ONE[4]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_22, Q => 
        \U50_PATTERNS/U4A_REGCROSS/SAMP_TWO[4]_net_1\);
    
    HIEFFPLA_INST_0_47101 : AND2
      port map(A => \U_ELK12_CH/ELK_TX_DAT[1]\, B => 
        \U_ELK12_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118558);
    
    \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117060, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_26, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[1]_net_1\);
    
    HIEFFPLA_INST_0_56245 : AND2A
      port map(A => DCB_SALT_SEL_c, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/RECD_SER_WORD[5]_net_1\, 
        Y => \TFC_RX_SER_WORD[5]\);
    
    HIEFFPLA_INST_0_47443 : MX2
      port map(A => \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\, 
        B => \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[11]_net_1\, S => 
        \BIT_OS_SEL_3[2]\, Y => HIEFFPLA_NET_0_118491);
    
    HIEFFPLA_INST_0_41800 : MX2
      port map(A => HIEFFPLA_NET_0_119668, B => 
        \U50_PATTERNS/ELINK_RWA[8]\, S => 
        \U50_PATTERNS/SM_BANK_SEL_0[20]\, Y => 
        HIEFFPLA_NET_0_119693);
    
    \U_ELK9_CH/U_SLAVE_1ELK/Q[0]\ : DFN1C0
      port map(D => \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/Q[0]_net_1\);
    
    \U_ELK19_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]\ : DFN1C0
      port map(D => \U_ELK19_CH/U_SLAVE_1ELK/Q[5]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]_net_1\);
    
    HIEFFPLA_INST_0_46455 : AND3C
      port map(A => HIEFFPLA_NET_0_118674, B => 
        HIEFFPLA_NET_0_119577, C => HIEFFPLA_NET_0_118679, Y => 
        HIEFFPLA_NET_0_118687);
    
    HIEFFPLA_INST_0_44800 : MX2
      port map(A => USB_OE_BI, B => HIEFFPLA_NET_0_119044, S => 
        HIEFFPLA_NET_0_119043, Y => HIEFFPLA_NET_0_119045);
    
    \U_EXEC_MASTER/MPOR_B_22\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117787, CLK => CLK_40M_GL, CLR
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_1\, Q => 
        P_MASTER_POR_B_c_22);
    
    \U_ELK7_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL\ : DFN1C0
      port map(D => 
        \U_ELK7_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL_net_1\);
    
    \U_ELK19_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]\ : DFN1C0
      port map(D => \U_ELK19_CH/U_SLAVE_1ELK/Q[10]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]_net_1\);
    
    HIEFFPLA_INST_0_54545 : NAND2B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[3]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[0]_net_1\, Y => 
        HIEFFPLA_NET_0_117252);
    
    \U50_PATTERNS/ELINK_DINA_15[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119819, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_16, Q => 
        \U50_PATTERNS/ELINK_DINA_15[4]\);
    
    \U200B_ELINKS/GP_PG_SM_0[10]\ : DFN1P0
      port map(D => HIEFFPLA_NET_0_120227, CLK => CLK_40M_GL, PRE
         => P_MASTER_POR_B_c_34_0, Q => 
        \U200B_ELINKS/GP_PG_SM_0[10]_net_1\);
    
    HIEFFPLA_INST_0_52129 : NAND2A
      port map(A => HIEFFPLA_NET_0_117629, B => 
        HIEFFPLA_NET_0_117631, Y => HIEFFPLA_NET_0_117630);
    
    HIEFFPLA_INST_0_46062 : AND3A
      port map(A => HIEFFPLA_NET_0_119376, B => 
        \U50_PATTERNS/TFC_STRT_ADDR[6]\, C => 
        HIEFFPLA_NET_0_119431, Y => HIEFFPLA_NET_0_118775);
    
    HIEFFPLA_INST_0_57211 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_3[4]\, B => 
        HIEFFPLA_NET_0_116703, S => HIEFFPLA_NET_0_117120, Y => 
        HIEFFPLA_NET_0_116721);
    
    HIEFFPLA_INST_0_44304 : MX2B
      port map(A => HIEFFPLA_NET_0_119145, B => 
        HIEFFPLA_NET_0_119156, S => 
        \U50_PATTERNS/U4A_REGCROSS/SYNC_SM[0]_net_1\, Y => 
        HIEFFPLA_NET_0_119146);
    
    \U_ELK10_CH/U_ELK1_SERDAT_SOURCE/SERDAT[4]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118639, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_17, Q => 
        \U_ELK10_CH/ELK_TX_DAT[4]\);
    
    HIEFFPLA_INST_0_37791 : AND3
      port map(A => HIEFFPLA_NET_0_120223, B => 
        HIEFFPLA_NET_0_120199, C => HIEFFPLA_NET_0_120233, Y => 
        HIEFFPLA_NET_0_120206);
    
    \U50_PATTERNS/ELINK_DINA_8[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119725, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_18, Q => 
        \U50_PATTERNS/ELINK_DINA_8[2]\);
    
    HIEFFPLA_INST_0_40092 : AOI1C
      port map(A => \U50_PATTERNS/ELINK_BLKA[12]\, B => 
        HIEFFPLA_NET_0_119659, C => HIEFFPLA_NET_0_119908, Y => 
        HIEFFPLA_NET_0_119909);
    
    \U_TFC_SERDAT_SOURCE/SERDAT[4]\ : DFN1C0
      port map(D => \U_TFC_SERDAT_SOURCE/N_SERDAT[4]\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \TFC_TX_DAT[4]\);
    
    \U_ELK4_CH/U_ELK1_CMD_TX/SER_OUT_RI\ : DFI1C0
      port map(D => 
        \U_ELK4_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_4, QN
         => \U_ELK4_CH/U_ELK1_CMD_TX/SER_OUT_RI_i\);
    
    HIEFFPLA_INST_0_45005 : NAND3C
      port map(A => HIEFFPLA_NET_0_119485, B => 
        HIEFFPLA_NET_0_119460, C => HIEFFPLA_NET_0_118993, Y => 
        HIEFFPLA_NET_0_119002);
    
    HIEFFPLA_INST_0_40043 : MX2
      port map(A => HIEFFPLA_NET_0_119888, B => 
        \U50_PATTERNS/ELINK_BLKA[5]\, S => 
        \U50_PATTERNS/SM_BANK_SEL[20]\, Y => 
        HIEFFPLA_NET_0_119920);
    
    \U_ELK8_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117880, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_15, Q => 
        \U_ELK8_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]_net_1\);
    
    HIEFFPLA_INST_0_57599 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_5[7]\, B => 
        HIEFFPLA_NET_0_116637, S => HIEFFPLA_NET_0_117121, Y => 
        HIEFFPLA_NET_0_116654);
    
    HIEFFPLA_INST_0_39371 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_2[1]\, B => 
        HIEFFPLA_NET_0_119523, S => HIEFFPLA_NET_0_119278, Y => 
        HIEFFPLA_NET_0_119998);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_29[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116043, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_16_0, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_29[2]\);
    
    \U50_PATTERNS/U4E_REGCROSS/LOCAL_REG_VAL_6[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119056, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_0_0, Q => \OP_MODE_c_6[1]\);
    
    HIEFFPLA_INST_0_42251 : OR3B
      port map(A => \U50_PATTERNS/RD_USB_ADBUS[1]\, B => 
        \U50_PATTERNS/RD_USB_ADBUS[0]\, C => 
        HIEFFPLA_NET_0_119585, Y => HIEFFPLA_NET_0_119590);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_2[8]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116747, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_6, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_2[8]\);
    
    \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[6]\ : DFN1C0
      port map(D => \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\);
    
    \U_ELK19_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118246, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_7, Q => 
        \U_ELK19_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]_net_1\);
    
    \U50_PATTERNS/ELINK_DINA_1[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119776, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_7, Q => 
        \U50_PATTERNS/ELINK_DINA_1[7]\);
    
    HIEFFPLA_INST_0_54189 : MX2
      port map(A => HIEFFPLA_NET_0_116362, B => 
        HIEFFPLA_NET_0_116556, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_1[3]_net_1\, Y
         => HIEFFPLA_NET_0_117297);
    
    HIEFFPLA_INST_0_58341 : AOI1A
      port map(A => HIEFFPLA_NET_0_116708, B => 
        HIEFFPLA_NET_0_116804, C => HIEFFPLA_NET_0_117396, Y => 
        HIEFFPLA_NET_0_116532);
    
    HIEFFPLA_INST_0_53997 : MX2
      port map(A => HIEFFPLA_NET_0_117289, B => 
        HIEFFPLA_NET_0_117385, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[2]_net_1\, Y
         => HIEFFPLA_NET_0_117322);
    
    HIEFFPLA_INST_0_48511 : MX2
      port map(A => HIEFFPLA_NET_0_118320, B => 
        HIEFFPLA_NET_0_118315, S => \BIT_OS_SEL_3[0]\, Y => 
        \U_ELK17_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[3]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_115925, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_9, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[5]\);
    
    \U50_PATTERNS/WR_XFER_TYPE[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118686, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c, Q => 
        \U50_PATTERNS/WR_XFER_TYPE[3]_net_1\);
    
    HIEFFPLA_INST_0_56779 : XA1B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_0[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_0[0]\, C => 
        HIEFFPLA_NET_0_117179, Y => HIEFFPLA_NET_0_116799);
    
    HIEFFPLA_INST_0_41332 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_5[2]\, B => 
        HIEFFPLA_NET_0_119575, S => HIEFFPLA_NET_0_119251, Y => 
        HIEFFPLA_NET_0_119749);
    
    \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[13]\ : DFN1C0
      port map(D => \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[13]_net_1\);
    
    HIEFFPLA_INST_0_46340 : AO1
      port map(A => HIEFFPLA_NET_0_119276, B => 
        \U50_PATTERNS/ELINK_DOUTA_10[2]\, C => 
        HIEFFPLA_NET_0_118712, Y => HIEFFPLA_NET_0_118713);
    
    \U_MASTER_DES/U13C_MASTER_DESER/Q[7]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[7]_net_1\, CLK => 
        CCC_160M_FXD, CLR => P_MASTER_POR_B_c_34, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/Q[7]_net_1\);
    
    \U_ELK9_CH/U_ELK1_SERDAT_SOURCE/SERDAT[7]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117826, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_7, Q => 
        \U_ELK9_CH/ELK_TX_DAT[7]\);
    
    HIEFFPLA_INST_0_39479 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_3[5]\, B => 
        HIEFFPLA_NET_0_119518, S => HIEFFPLA_NET_0_119247, Y => 
        HIEFFPLA_NET_0_119986);
    
    HIEFFPLA_INST_0_51714 : NAND2B
      port map(A => 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM[4]_net_1\, B => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[40]_net_1\, Y => 
        HIEFFPLA_NET_0_117712);
    
    HIEFFPLA_INST_0_45956 : NAND3C
      port map(A => HIEFFPLA_NET_0_118948, B => 
        HIEFFPLA_NET_0_118836, C => HIEFFPLA_NET_0_118957, Y => 
        HIEFFPLA_NET_0_118802);
    
    \P_ELK0_SYNC_DET_pad/U0/U1\ : IOTRI_OB_EB
      port map(D => P_ELK0_SYNC_DET_c, E => \VCC\, DOUT => 
        \P_ELK0_SYNC_DET_pad/U0/NET1\, EOUT => 
        \P_ELK0_SYNC_DET_pad/U0/NET2\);
    
    HIEFFPLA_INST_0_51732 : AXOI5
      port map(A => HIEFFPLA_NET_0_117674, B => 
        HIEFFPLA_NET_0_117630, C => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[0]\, Y => 
        HIEFFPLA_NET_0_117698);
    
    HIEFFPLA_INST_0_47166 : MX2
      port map(A => HIEFFPLA_NET_0_118531, B => 
        HIEFFPLA_NET_0_118544, S => \BIT_OS_SEL_4[1]\, Y => 
        HIEFFPLA_NET_0_118540);
    
    HIEFFPLA_INST_0_42347 : AND3A
      port map(A => HIEFFPLA_NET_0_119596, B => 
        HIEFFPLA_NET_0_119586, C => 
        \U50_PATTERNS/RD_USB_ADBUS[7]\, Y => 
        HIEFFPLA_NET_0_119561);
    
    \U_ELK7_CH/U_ELK1_CMD_TX/SER_OUT_FDEL\ : DFN1C0
      port map(D => \U_ELK7_CH/U_ELK1_CMD_TX/SER_OUT_FI_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_12, Q
         => \U_ELK7_CH/ELK_OUT_F\);
    
    HIEFFPLA_INST_0_45279 : AO1
      port map(A => HIEFFPLA_NET_0_119277, B => 
        \U50_PATTERNS/ELINK_DOUTA_11[6]\, C => 
        HIEFFPLA_NET_0_118839, Y => HIEFFPLA_NET_0_118952);
    
    \U_ELK9_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117840, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_4, Q => 
        \U_ELK9_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]_net_1\);
    
    \U_ELK18_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U1\ : IOBI_ID_OD_EB
      port map(DR => \U_ELK18_CH/ELK_OUT_R\, DF => 
        \U_ELK18_CH/ELK_OUT_F\, CLR => \GND\, E => 
        \AFLSDF_INV_30\, ICLK => CCC_160M_ADJ, OCLK => 
        CCC_160M_FXD, YIN => 
        \U_ELK18_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\, DOUT => 
        \U_ELK18_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, EOUT => 
        \U_ELK18_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET2\, YR => 
        \U_ELK18_CH/ELK_IN_DDR_R\, YF => 
        \U_ELK18_CH/ELK_IN_DDR_F\);
    
    \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[9]\ : DFN1C0
      port map(D => 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\);
    
    HIEFFPLA_INST_0_37102 : AND3B
      port map(A => \U200A_TFC/LOC_STRT_ADDR[1]\, B => 
        HIEFFPLA_NET_0_120293, C => HIEFFPLA_NET_0_120328, Y => 
        HIEFFPLA_NET_0_120347);
    
    \U_ELK6_CH/U_SLAVE_1ELK/RECD_SER_WORD[1]\ : DFN1C0
      port map(D => \U_ELK6_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[1]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_6[1]\);
    
    HIEFFPLA_INST_0_57473 : AND3A
      port map(A => HIEFFPLA_NET_0_116686, B => 
        HIEFFPLA_NET_0_116735, C => HIEFFPLA_NET_0_116620, Y => 
        HIEFFPLA_NET_0_116675);
    
    \U_ELK12_CH/U_SLAVE_1ELK/Q[2]\ : DFN1C0
      port map(D => \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/Q[2]_net_1\);
    
    HIEFFPLA_INST_0_45443 : AO1
      port map(A => HIEFFPLA_NET_0_119283, B => 
        \U50_PATTERNS/ELINK_DOUTA_13[0]\, C => 
        HIEFFPLA_NET_0_118812, Y => HIEFFPLA_NET_0_118913);
    
    HIEFFPLA_INST_0_52576 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_1[3]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_2[3]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[0]\, Y => 
        HIEFFPLA_NET_0_117545);
    
    \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[12]\ : DFN1C0
      port map(D => 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[12]_net_1\);
    
    \U50_PATTERNS/U118_PATT_ELINK_BLK/DPRT_512X9_SRAM_R0C0\ : 
        RAM4K9
      generic map(MEMORYFILE => "DPRT_512X9_SRAM_R0C0.mem")

      port map(ADDRA11 => AFLSDF_GND, ADDRA10 => AFLSDF_GND, 
        ADDRA9 => AFLSDF_GND, ADDRA8 => \GND\, ADDRA7 => 
        \U50_PATTERNS/ELINK_ADDRA_18[7]\, ADDRA6 => 
        \U50_PATTERNS/ELINK_ADDRA_18[6]\, ADDRA5 => 
        \U50_PATTERNS/ELINK_ADDRA_18[5]\, ADDRA4 => 
        \U50_PATTERNS/ELINK_ADDRA_18[4]\, ADDRA3 => 
        \U50_PATTERNS/ELINK_ADDRA_18[3]\, ADDRA2 => 
        \U50_PATTERNS/ELINK_ADDRA_18[2]\, ADDRA1 => 
        \U50_PATTERNS/ELINK_ADDRA_18[1]\, ADDRA0 => 
        \U50_PATTERNS/ELINK_ADDRA_18[0]\, ADDRB11 => AFLSDF_GND, 
        ADDRB10 => AFLSDF_GND, ADDRB9 => AFLSDF_GND, ADDRB8 => 
        \GND\, ADDRB7 => \ELKS_ADDRB[7]\, ADDRB6 => 
        \ELKS_ADDRB_0[6]\, ADDRB5 => \ELKS_ADDRB[5]\, ADDRB4 => 
        \ELKS_ADDRB_0[4]\, ADDRB3 => \ELKS_ADDRB[3]\, ADDRB2 => 
        \ELKS_ADDRB_0[2]\, ADDRB1 => \ELKS_ADDRB[1]\, ADDRB0 => 
        \ELKS_ADDRB[0]\, DINA8 => \GND\, DINA7 => 
        \U50_PATTERNS/ELINK_DINA_18[7]\, DINA6 => 
        \U50_PATTERNS/ELINK_DINA_18[6]\, DINA5 => 
        \U50_PATTERNS/ELINK_DINA_18[5]\, DINA4 => 
        \U50_PATTERNS/ELINK_DINA_18[4]\, DINA3 => 
        \U50_PATTERNS/ELINK_DINA_18[3]\, DINA2 => 
        \U50_PATTERNS/ELINK_DINA_18[2]\, DINA1 => 
        \U50_PATTERNS/ELINK_DINA_18[1]\, DINA0 => 
        \U50_PATTERNS/ELINK_DINA_18[0]\, DINB8 => \GND\, DINB7
         => \ELK_RX_SER_WORD_18[7]\, DINB6 => 
        \ELK_RX_SER_WORD_18[6]\, DINB5 => \ELK_RX_SER_WORD_18[5]\, 
        DINB4 => \ELK_RX_SER_WORD_18[4]\, DINB3 => 
        \ELK_RX_SER_WORD_18[3]\, DINB2 => \ELK_RX_SER_WORD_18[2]\, 
        DINB1 => \ELK_RX_SER_WORD_18[1]\, DINB0 => 
        \ELK_RX_SER_WORD_18[0]\, WIDTHA0 => \VCC\, WIDTHA1 => 
        \VCC\, WIDTHB0 => \VCC\, WIDTHB1 => \VCC\, PIPEA => \VCC\, 
        PIPEB => \VCC\, WMODEA => \GND\, WMODEB => \GND\, BLKA
         => \U50_PATTERNS/ELINK_BLKA[18]\, BLKB => 
        ELKS_RAM_BLKB_EN, WENA => \U50_PATTERNS/ELINK_RWA[18]\, 
        WENB => ELKS_RWB, CLKA => CLK60MHZ, CLKB => CLK_40M_GL, 
        RESET => P_USB_MASTER_EN_c_0, DOUTA8 => OPEN, DOUTA7 => 
        \U50_PATTERNS/ELINK_DOUTA_18[7]\, DOUTA6 => 
        \U50_PATTERNS/ELINK_DOUTA_18[6]\, DOUTA5 => 
        \U50_PATTERNS/ELINK_DOUTA_18[5]\, DOUTA4 => 
        \U50_PATTERNS/ELINK_DOUTA_18[4]\, DOUTA3 => 
        \U50_PATTERNS/ELINK_DOUTA_18[3]\, DOUTA2 => 
        \U50_PATTERNS/ELINK_DOUTA_18[2]\, DOUTA1 => 
        \U50_PATTERNS/ELINK_DOUTA_18[1]\, DOUTA0 => 
        \U50_PATTERNS/ELINK_DOUTA_18[0]\, DOUTB8 => OPEN, DOUTB7
         => \PATT_ELK_DAT_18[7]\, DOUTB6 => \PATT_ELK_DAT_18[6]\, 
        DOUTB5 => \PATT_ELK_DAT_18[5]\, DOUTB4 => 
        \PATT_ELK_DAT_18[4]\, DOUTB3 => \PATT_ELK_DAT_18[3]\, 
        DOUTB2 => \PATT_ELK_DAT_18[2]\, DOUTB1 => 
        \PATT_ELK_DAT_18[1]\, DOUTB0 => \PATT_ELK_DAT_18[0]\);
    
    \U_EXEC_MASTER/DEL_CNT[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117795, CLK => CLK_40M_GL, CLR
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i\, Q => 
        \U_EXEC_MASTER/DEL_CNT[0]\);
    
    HIEFFPLA_INST_0_60660 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_13[3]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_14[3]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_3[0]\, Y => 
        HIEFFPLA_NET_0_116236);
    
    HIEFFPLA_INST_0_48586 : MX2
      port map(A => 
        \U_ELK18_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]_net_1\, B => 
        \U_ELK18_CH/ELK_TX_DAT[4]\, S => 
        \U_ELK18_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118290);
    
    HIEFFPLA_INST_0_56392 : NAND3C
      port map(A => HIEFFPLA_NET_0_116831, B => 
        HIEFFPLA_NET_0_116847, C => HIEFFPLA_NET_0_116855, Y => 
        HIEFFPLA_NET_0_116879);
    
    HIEFFPLA_INST_0_54979 : AO1C
      port map(A => HIEFFPLA_NET_0_117216, B => 
        HIEFFPLA_NET_0_117164, C => HIEFFPLA_NET_0_117180, Y => 
        HIEFFPLA_NET_0_117149);
    
    HIEFFPLA_INST_0_50111 : NAND2B
      port map(A => \OP_MODE_c_4[1]\, B => \PATT_ELK_DAT_5[2]\, Y
         => HIEFFPLA_NET_0_118011);
    
    HIEFFPLA_INST_0_49441 : MX2
      port map(A => HIEFFPLA_NET_0_118135, B => 
        HIEFFPLA_NET_0_118131, S => \BIT_OS_SEL[1]\, Y => 
        HIEFFPLA_NET_0_118130);
    
    HIEFFPLA_INST_0_45334 : AO1
      port map(A => HIEFFPLA_NET_0_119244, B => 
        \U50_PATTERNS/ELINK_DOUTA_2[7]\, C => 
        HIEFFPLA_NET_0_118821, Y => HIEFFPLA_NET_0_118938);
    
    \U_ELK15_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0\ : DFN1C0
      port map(D => CLK_40M_GL, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_8, Q => 
        \U_ELK15_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0_net_1\);
    
    HIEFFPLA_INST_0_44647 : XO1
      port map(A => \U50_PATTERNS/U4D_REGCROSS/SAMP_TWO[6]_net_1\, 
        B => \ELKS_STOP_ADDR[6]\, C => HIEFFPLA_NET_0_119074, Y
         => HIEFFPLA_NET_0_119075);
    
    \U_ELK2_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]\ : DFN1C0
      port map(D => \U_ELK2_CH/U_SLAVE_1ELK/Q[10]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]_net_1\);
    
    HIEFFPLA_INST_0_57779 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_6[8]\, B => 
        HIEFFPLA_NET_0_116607, S => HIEFFPLA_NET_0_117599, Y => 
        HIEFFPLA_NET_0_116624);
    
    HIEFFPLA_INST_0_45787 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_7[3]\, C => 
        \U50_PATTERNS/SM_BANK_SEL[12]\, Y => 
        HIEFFPLA_NET_0_118842);
    
    HIEFFPLA_INST_0_161271 : DFN1C0
      port map(D => \U_ELK16_CH/U_ELK1_CMD_TX/START_RISE_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_10, Q
         => HIEFFPLA_NET_0_161284);
    
    HIEFFPLA_INST_0_42564 : AND3A
      port map(A => HIEFFPLA_NET_0_119449, B => 
        HIEFFPLA_NET_0_119494, C => HIEFFPLA_NET_0_119511, Y => 
        HIEFFPLA_NET_0_119510);
    
    \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[13]\ : DFN1C0
      port map(D => 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]_net_1\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[13]_net_1\);
    
    \U_ELK13_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2\ : IOPADN_BI
      port map(DB => \U_ELK13_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, 
        E => \U_ELK13_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET3\, PAD
         => ELK13_DAT_N, N2POUT => 
        \U_ELK13_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2_N2P\);
    
    HIEFFPLA_INST_0_50905 : MX2
      port map(A => HIEFFPLA_NET_0_117863, B => 
        HIEFFPLA_NET_0_117861, S => \BIT_OS_SEL_3[1]\, Y => 
        HIEFFPLA_NET_0_117865);
    
    HIEFFPLA_INST_0_41772 : MX2
      port map(A => HIEFFPLA_NET_0_119675, B => 
        \U50_PATTERNS/ELINK_RWA[4]\, S => 
        \U50_PATTERNS/SM_BANK_SEL_0[20]\, Y => 
        HIEFFPLA_NET_0_119697);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_1[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116787, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_4, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_1[1]\);
    
    HIEFFPLA_INST_0_48174 : MX2
      port map(A => \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\, 
        B => \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\, S => 
        \BIT_OS_SEL_1[2]\, Y => HIEFFPLA_NET_0_118358);
    
    HIEFFPLA_INST_0_40161 : AOI1D
      port map(A => HIEFFPLA_NET_0_119389, B => 
        HIEFFPLA_NET_0_119464, C => 
        \U50_PATTERNS/SM_BANK_SEL[13]\, Y => 
        HIEFFPLA_NET_0_119885);
    
    HIEFFPLA_INST_0_37654 : NAND2B
      port map(A => \U200B_ELINKS/LOC_STRT_ADDR[7]\, B => 
        HIEFFPLA_NET_0_120190, Y => HIEFFPLA_NET_0_120239);
    
    \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[10]\ : DFN1C0
      port map(D => \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\);
    
    \U50_PATTERNS/U4C_REGCROSS/LOCAL_REG_VAL[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119108, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_21, Q => \ELKS_STRT_ADDR[4]\);
    
    HIEFFPLA_INST_0_61850 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_27[1]\, B => 
        HIEFFPLA_NET_0_117114, S => HIEFFPLA_NET_0_117196, Y => 
        HIEFFPLA_NET_0_116069);
    
    \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[12]\ : DFN1C0
      port map(D => 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[12]_net_1\);
    
    HIEFFPLA_INST_0_54891 : NAND2B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_0[6]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_0[8]_net_1\, Y => 
        HIEFFPLA_NET_0_117179);
    
    HIEFFPLA_INST_0_55072 : AND3
      port map(A => HIEFFPLA_NET_0_117101, B => 
        HIEFFPLA_NET_0_117360, C => HIEFFPLA_NET_0_117415, Y => 
        HIEFFPLA_NET_0_117127);
    
    HIEFFPLA_INST_0_48368 : NAND2B
      port map(A => \OP_MODE_c_6[1]\, B => \PATT_ELK_DAT_17[2]\, 
        Y => HIEFFPLA_NET_0_118326);
    
    HIEFFPLA_INST_0_55850 : MX2
      port map(A => HIEFFPLA_NET_0_116994, B => 
        HIEFFPLA_NET_0_116968, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[1]\, Y => 
        HIEFFPLA_NET_0_116982);
    
    HIEFFPLA_INST_0_49461 : MX2
      port map(A => HIEFFPLA_NET_0_118133, B => 
        HIEFFPLA_NET_0_118129, S => \BIT_OS_SEL[1]\, Y => 
        HIEFFPLA_NET_0_118127);
    
    \U_ELK12_CH/U_SLAVE_1ELK/RECD_SER_WORD[3]\ : DFN1C0
      port map(D => \U_ELK12_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[3]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_12[3]\);
    
    \U_ELK5_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL\ : DFN1C0
      port map(D => \U_ELK5_CH/ELK_IN_F_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL_net_1\);
    
    \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[5]\ : DFN1C0
      port map(D => 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\);
    
    HIEFFPLA_INST_0_61055 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_19[1]\, B => 
        HIEFFPLA_NET_0_117114, S => HIEFFPLA_NET_0_117170, Y => 
        HIEFFPLA_NET_0_116179);
    
    HIEFFPLA_INST_0_45528 : AO1A
      port map(A => HIEFFPLA_NET_0_119475, B => 
        \U50_PATTERNS/ELINKS_STOP_ADDR[1]\, C => 
        HIEFFPLA_NET_0_118811, Y => HIEFFPLA_NET_0_118896);
    
    \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[3]\ : DFN1C0
      port map(D => 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[3]_net_1\);
    
    HIEFFPLA_INST_0_45689 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_19[1]\, C => 
        \U50_PATTERNS/SM_BANK_SEL[0]\, Y => HIEFFPLA_NET_0_118864);
    
    HIEFFPLA_INST_0_115745 : NAND2A
      port map(A => \ELKS_ADDRB[0]\, B => 
        \U200B_ELINKS/LOC_STOP_ADDR[0]\, Y => 
        HIEFFPLA_NET_0_115806);
    
    \U200B_ELINKS/ADDR_POINTER[7]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120248, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_32, Q => \ELKS_ADDRB[7]\);
    
    HIEFFPLA_INST_0_61190 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_1[4]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_2[4]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_1[0]\, Y => 
        HIEFFPLA_NET_0_116161);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_8[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116292, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_5, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_8[1]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_22[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116129, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_5, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_22[1]\);
    
    HIEFFPLA_INST_0_46634 : MX2
      port map(A => \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\, 
        B => \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\, S => 
        \BIT_OS_SEL_5[2]\, Y => HIEFFPLA_NET_0_118635);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_30[4]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116026, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_8, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_30[4]\);
    
    HIEFFPLA_INST_0_55319 : AO1A
      port map(A => HIEFFPLA_NET_0_115917, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[0]_net_1\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[1]_net_1\, Y => 
        HIEFFPLA_NET_0_117061);
    
    \U_ELK17_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]\ : DFN1C0
      port map(D => \U_ELK17_CH/U_SLAVE_1ELK/Q[1]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]_net_1\);
    
    HIEFFPLA_INST_0_61103 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_3[3]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_19[3]\, S
         => \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_1[4]_net_1\, 
        Y => HIEFFPLA_NET_0_116173);
    
    \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[14]\ : DFN1C0
      port map(D => 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[14]_net_1\);
    
    \U50_PATTERNS/ELINK_DINA_4[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119757, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_13, Q => 
        \U50_PATTERNS/ELINK_DINA_4[2]\);
    
    HIEFFPLA_INST_0_56942 : NAND3
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_1[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_1[2]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_1[0]\, Y => 
        HIEFFPLA_NET_0_116769);
    
    HIEFFPLA_INST_0_56606 : AND3
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[10]_net_1\, B
         => HIEFFPLA_NET_0_117424, C => HIEFFPLA_NET_0_117427, Y
         => HIEFFPLA_NET_0_116829);
    
    \U_ELK15_CH/U_SLAVE_1ELK/RECD_SER_WORD[7]\ : DFN1C0
      port map(D => \U_ELK15_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[7]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_15[7]\);
    
    HIEFFPLA_INST_0_44443 : AND2
      port map(A => \U50_PATTERNS/U4C_REGCROSS/DELCNT[0]_net_1\, 
        B => \U50_PATTERNS/U4C_REGCROSS/DELCNT[1]_net_1\, Y => 
        HIEFFPLA_NET_0_119114);
    
    HIEFFPLA_INST_0_48871 : NAND2B
      port map(A => \OP_MODE_c_6[1]\, B => \PATT_ELK_DAT_19[7]\, 
        Y => HIEFFPLA_NET_0_118231);
    
    HIEFFPLA_INST_0_38894 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_14[4]\, B => 
        HIEFFPLA_NET_0_119519, S => HIEFFPLA_NET_0_119249, Y => 
        HIEFFPLA_NET_0_120051);
    
    \U_ELK11_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118604, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_11, Q => 
        \U_ELK11_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]_net_1\);
    
    HIEFFPLA_INST_0_48495 : MX2
      port map(A => HIEFFPLA_NET_0_118310, B => 
        HIEFFPLA_NET_0_118306, S => \BIT_OS_SEL_3[0]\, Y => 
        \U_ELK17_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[1]\);
    
    \P_ELK0_SYNC_DET_pad/U0/U0\ : IOPAD_TRI_U
      port map(D => \P_ELK0_SYNC_DET_pad/U0/NET1\, E => 
        \P_ELK0_SYNC_DET_pad/U0/NET2\, PAD => P_ELK0_SYNC_DET);
    
    HIEFFPLA_INST_0_161258 : DFN1C0
      port map(D => \TFC_IN_R\, CLK => CCC_160M_ADJ, CLR => 
        P_MASTER_POR_B_c_26, Q => HIEFFPLA_NET_0_161297);
    
    \U_ELK5_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]\ : DFN1C0
      port map(D => \U_ELK5_CH/U_SLAVE_1ELK/Q[3]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]_net_1\);
    
    HIEFFPLA_INST_0_44995 : OA1A
      port map(A => HIEFFPLA_NET_0_119379, B => 
        HIEFFPLA_NET_0_119371, C => \U50_PATTERNS/USB_TXE_B\, Y
         => HIEFFPLA_NET_0_119004);
    
    \U61_TS_WR_BUF/_TRIBUFF_F_24U[0]_/U0/U1\ : IOTRI_OB_EB
      port map(D => USB_WR_BI, E => P_USB_MASTER_EN_c, DOUT => 
        \U61_TS_WR_BUF/\\\\TRIBUFF_F_24U[0]\\\\/U0/NET1\, EOUT
         => \U61_TS_WR_BUF/\\\\TRIBUFF_F_24U[0]\\\\/U0/NET2\);
    
    \U50_PATTERNS/ELINK_DINA_1[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119782, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_7, Q => 
        \U50_PATTERNS/ELINK_DINA_1[1]\);
    
    HIEFFPLA_INST_0_48614 : AND2
      port map(A => CLK_40M_GL, B => 
        \U_ELK18_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0_net_1\, Y => 
        HIEFFPLA_NET_0_118284);
    
    \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[46]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117726, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_18, Q => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[46]\);
    
    \U50_PATTERNS/ELINK_DINA_2[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119770, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_9, Q => 
        \U50_PATTERNS/ELINK_DINA_2[5]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_3[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116010, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_11, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_3[0]\);
    
    HIEFFPLA_INST_0_51503 : NOR3B
      port map(A => \U_EXEC_MASTER/CCC_1_LOCK_STAT_1D_net_1\, B
         => HIEFFPLA_NET_0_117764, C => 
        \U_EXEC_MASTER/PRESCALE[0]\, Y => HIEFFPLA_NET_0_117762);
    
    HIEFFPLA_INST_0_41080 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_1[6]\, B => 
        HIEFFPLA_NET_0_119566, S => HIEFFPLA_NET_0_119243, Y => 
        HIEFFPLA_NET_0_119777);
    
    HIEFFPLA_INST_0_59581 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_29[3]\, B => 
        HIEFFPLA_NET_0_116368, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_0[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116375);
    
    HIEFFPLA_INST_0_56037 : MX2
      port map(A => HIEFFPLA_NET_0_117020, B => 
        HIEFFPLA_NET_0_116036, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[2]\, Y => 
        HIEFFPLA_NET_0_116958);
    
    HIEFFPLA_INST_0_42213 : MX2
      port map(A => \U50_PATTERNS/OP_MODE_T[7]\, B => 
        \U50_PATTERNS/RD_USB_ADBUS[7]\, S => 
        HIEFFPLA_NET_0_119440, Y => HIEFFPLA_NET_0_119602);
    
    \U_ELK6_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U0\ : IOPADP_BI
      port map(N2PIN => 
        \U_ELK6_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2_N2P\, D => 
        \U_ELK6_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, E => 
        \U_ELK6_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET2\, PAD => 
        ELK6_DAT_P, Y => 
        \U_ELK6_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\);
    
    HIEFFPLA_INST_0_50792 : MX2
      port map(A => HIEFFPLA_NET_0_117889, B => 
        HIEFFPLA_NET_0_117910, S => \BIT_OS_SEL_4[1]\, Y => 
        HIEFFPLA_NET_0_117891);
    
    HIEFFPLA_INST_0_43201 : AND3A
      port map(A => \U50_PATTERNS/REG_STATE_0[4]_net_1\, B => 
        HIEFFPLA_NET_0_119552, C => HIEFFPLA_NET_0_119338, Y => 
        HIEFFPLA_NET_0_119348);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_3[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116009, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_11, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_3[1]\);
    
    \U200B_ELINKS/GP_PG_SM[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120216, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_29, Q => 
        \U200B_ELINKS/GP_PG_SM[1]_net_1\);
    
    \U_ELK9_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117842, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_3, Q => 
        \U_ELK9_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]_net_1\);
    
    HIEFFPLA_INST_0_42117 : MX2
      port map(A => \U50_PATTERNS/OP_MODE[3]\, B => 
        \U50_PATTERNS/OP_MODE_T[3]\, S => HIEFFPLA_NET_0_119472, 
        Y => HIEFFPLA_NET_0_119614);
    
    \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[7]\ : DFN1C0
      port map(D => \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\);
    
    HIEFFPLA_INST_0_61922 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_11[4]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_27[4]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_2[4]_net_1\, Y
         => HIEFFPLA_NET_0_116059);
    
    \U50_PATTERNS/USB_WR_BI/U1\ : DFN1P0
      port map(D => HIEFFPLA_NET_0_118990, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_19, Q => USB_WR_BI);
    
    \U_ELK16_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0\ : DFN1C0
      port map(D => CLK_40M_GL, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_8, Q => 
        \U_ELK16_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0_net_1\);
    
    \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[6]\ : DFN1C0
      port map(D => \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\);
    
    HIEFFPLA_INST_0_50310 : MX2
      port map(A => \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[0]_net_1\, B
         => \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\, S => 
        \BIT_OS_SEL_5[2]\, Y => HIEFFPLA_NET_0_117979);
    
    \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[10]\ : DFN1C0
      port map(D => 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]_net_1\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\);
    
    HIEFFPLA_INST_0_58311 : AO1A
      port map(A => HIEFFPLA_NET_0_117396, B => 
        HIEFFPLA_NET_0_116593, C => HIEFFPLA_NET_0_116536, Y => 
        HIEFFPLA_NET_0_116537);
    
    HIEFFPLA_INST_0_62409 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_5[2]\, 
        B => HIEFFPLA_NET_0_117131, S => HIEFFPLA_NET_0_117172, Y
         => HIEFFPLA_NET_0_115993);
    
    HIEFFPLA_INST_0_41485 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_7[3]\, B => 
        HIEFFPLA_NET_0_119574, S => HIEFFPLA_NET_0_119289, Y => 
        HIEFFPLA_NET_0_119732);
    
    HIEFFPLA_INST_0_40378 : MX2
      port map(A => HIEFFPLA_NET_0_119578, B => 
        \U50_PATTERNS/ELINK_DINA_11[0]\, S => 
        HIEFFPLA_NET_0_119280, Y => HIEFFPLA_NET_0_119855);
    
    HIEFFPLA_INST_0_54973 : AO1A
      port map(A => HIEFFPLA_NET_0_117082, B => 
        HIEFFPLA_NET_0_117086, C => HIEFFPLA_NET_0_117150, Y => 
        HIEFFPLA_NET_0_117151);
    
    HIEFFPLA_INST_0_38099 : NAND3B
      port map(A => HIEFFPLA_NET_0_120188, B => 
        \U200B_ELINKS/GP_PG_SM[1]_net_1\, C => \OP_MODE_c[6]\, Y
         => HIEFFPLA_NET_0_120153);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_5[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116659, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_11, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_5[2]\);
    
    HIEFFPLA_INST_0_53158 : MX2
      port map(A => HIEFFPLA_NET_0_117538, B => 
        HIEFFPLA_NET_0_117534, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_1[3]\, Y => 
        HIEFFPLA_NET_0_117458);
    
    HIEFFPLA_INST_0_50431 : MX2
      port map(A => HIEFFPLA_NET_0_117953, B => 
        HIEFFPLA_NET_0_117949, S => \BIT_OS_SEL_5[1]\, Y => 
        HIEFFPLA_NET_0_117951);
    
    HIEFFPLA_INST_0_37812 : AND2A
      port map(A => \OP_MODE[4]\, B => 
        \U200B_ELINKS/GP_PG_SM[6]_net_1\, Y => 
        HIEFFPLA_NET_0_120202);
    
    HIEFFPLA_INST_0_37253 : NAND2
      port map(A => HIEFFPLA_NET_0_120327, B => 
        \U200A_TFC/GP_PG_SM[7]_net_1\, Y => HIEFFPLA_NET_0_120313);
    
    HIEFFPLA_INST_0_46308 : NAND3C
      port map(A => HIEFFPLA_NET_0_118790, B => 
        HIEFFPLA_NET_0_118893, C => HIEFFPLA_NET_0_118719, Y => 
        HIEFFPLA_NET_0_118720);
    
    HIEFFPLA_INST_0_47216 : MX2
      port map(A => \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\, 
        B => \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[13]_net_1\, S => 
        \BIT_OS_SEL_4[2]\, Y => HIEFFPLA_NET_0_118533);
    
    HIEFFPLA_INST_0_43386 : MX2
      port map(A => \U50_PATTERNS/SM_BANK_SEL[14]\, B => 
        HIEFFPLA_NET_0_119223, S => HIEFFPLA_NET_0_118691, Y => 
        HIEFFPLA_NET_0_119317);
    
    HIEFFPLA_INST_0_50840 : MX2
      port map(A => 
        \U_ELK8_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]_net_1\, B => 
        \U_ELK8_CH/ELK_TX_DAT[3]\, S => 
        \U_ELK8_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_117882);
    
    \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[4]\ : DFN1C0
      port map(D => \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\);
    
    HIEFFPLA_INST_0_54561 : MX2
      port map(A => HIEFFPLA_NET_0_116496, B => 
        HIEFFPLA_NET_0_116279, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[3]_net_1\, Y => 
        HIEFFPLA_NET_0_117248);
    
    HIEFFPLA_INST_0_51122 : MX2
      port map(A => HIEFFPLA_NET_0_117821, B => 
        HIEFFPLA_NET_0_117817, S => \BIT_OS_SEL_2[1]\, Y => 
        HIEFFPLA_NET_0_117824);
    
    HIEFFPLA_INST_0_49702 : MX2
      port map(A => \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\, B
         => \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[13]_net_1\, S => 
        \BIT_OS_SEL_7[2]\, Y => HIEFFPLA_NET_0_118083);
    
    \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_SEL_4[1]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_BIT_OS_VAL[1]\, CLK
         => CLK_40M_GL, CLR => P_MASTER_POR_B_c_27_0, Q => 
        \BIT_OS_SEL_4[1]\);
    
    HIEFFPLA_INST_0_57150 : XA1B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_2[5]\, B => 
        HIEFFPLA_NET_0_116736, C => HIEFFPLA_NET_0_117179, Y => 
        HIEFFPLA_NET_0_116730);
    
    \U_ELK12_CH/U_SLAVE_1ELK/Q[12]\ : DFN1C0
      port map(D => \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/Q[12]_net_1\);
    
    \U_ELK10_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]\ : DFN1C0
      port map(D => \U_ELK10_CH/U_SLAVE_1ELK/Q[10]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]_net_1\);
    
    HIEFFPLA_INST_0_42101 : MX2
      port map(A => \U50_PATTERNS/OP_MODE[1]\, B => 
        \U50_PATTERNS/OP_MODE_T[1]\, S => HIEFFPLA_NET_0_119472, 
        Y => HIEFFPLA_NET_0_119616);
    
    HIEFFPLA_INST_0_41044 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_1[2]\, B => 
        HIEFFPLA_NET_0_119575, S => HIEFFPLA_NET_0_119243, Y => 
        HIEFFPLA_NET_0_119781);
    
    HIEFFPLA_INST_0_38227 : AND2A
      port map(A => HIEFFPLA_NET_0_119452, B => 
        \U50_PATTERNS/RD_USB_ADBUS[2]\, Y => 
        HIEFFPLA_NET_0_120133);
    
    \U_ELK18_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]\ : DFN1C0
      port map(D => \U_ELK18_CH/U_SLAVE_1ELK/Q[10]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]_net_1\);
    
    \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[7]\ : DFN1C0
      port map(D => 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\);
    
    HIEFFPLA_INST_0_56945 : AND3
      port map(A => HIEFFPLA_NET_0_117415, B => 
        HIEFFPLA_NET_0_117359, C => HIEFFPLA_NET_0_116774, Y => 
        HIEFFPLA_NET_0_116768);
    
    HIEFFPLA_INST_0_44046 : MX2
      port map(A => \U50_PATTERNS/TFC_STOP_ADDR_T[0]\, B => 
        \U50_PATTERNS/RD_USB_ADBUS[0]\, S => 
        HIEFFPLA_NET_0_119492, Y => HIEFFPLA_NET_0_119180);
    
    HIEFFPLA_INST_0_37192 : AND3B
      port map(A => \U200A_TFC/GP_PG_SM[0]_net_1\, B => 
        \U200A_TFC/GP_PG_SM[1]_net_1\, C => HIEFFPLA_NET_0_120334, 
        Y => HIEFFPLA_NET_0_120327);
    
    \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_5[4]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_115935, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_24_0, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_5[4]_net_1\);
    
    \U200B_ELINKS/ADDR_POINTER[6]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120171, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_32, Q => \ELKS_ADDRB[6]\);
    
    HIEFFPLA_INST_0_44641 : XOR2
      port map(A => \ELKS_STOP_ADDR[3]\, B => 
        \U50_PATTERNS/U4D_REGCROSS/SAMP_TWO[3]_net_1\, Y => 
        HIEFFPLA_NET_0_119077);
    
    \U_GEN_REF_CLK/GEN_40M_REFCNT[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117729, CLK => Y, CLR => 
        DEV_RST_B_c, Q => \U_GEN_REF_CLK/GEN_40M_REFCNT[2]_net_1\);
    
    \U_ELK11_CH/U_SLAVE_1ELK/Q[11]\ : DFN1C0
      port map(D => \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/Q[11]_net_1\);
    
    HIEFFPLA_INST_0_50656 : MX2
      port map(A => \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[2]_net_1\, B
         => \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\, S => 
        \BIT_OS_SEL_4[2]\, Y => HIEFFPLA_NET_0_117910);
    
    HIEFFPLA_INST_0_53371 : MX2
      port map(A => HIEFFPLA_NET_0_116325, B => 
        HIEFFPLA_NET_0_116381, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[3]_net_1\, Y
         => HIEFFPLA_NET_0_117419);
    
    HIEFFPLA_INST_0_45659 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_15[1]\, C => 
        \U50_PATTERNS/SM_BANK_SEL[4]\, Y => HIEFFPLA_NET_0_118870);
    
    \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[9]\ : DFN1C0
      port map(D => 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\);
    
    HIEFFPLA_INST_0_55006 : AO1A
      port map(A => HIEFFPLA_NET_0_117215, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_3[6]_net_1\, C => 
        HIEFFPLA_NET_0_117182, Y => HIEFFPLA_NET_0_117142);
    
    HIEFFPLA_INST_0_38231 : AND2A
      port map(A => HIEFFPLA_NET_0_119452, B => 
        \U50_PATTERNS/RD_USB_ADBUS[4]\, Y => 
        HIEFFPLA_NET_0_120131);
    
    HIEFFPLA_INST_0_55434 : AND3B
      port map(A => HIEFFPLA_NET_0_117187, B => 
        HIEFFPLA_NET_0_117087, C => HIEFFPLA_NET_0_117027, Y => 
        HIEFFPLA_NET_0_117038);
    
    HIEFFPLA_INST_0_45877 : AO1
      port map(A => HIEFFPLA_NET_0_119236, B => 
        \U50_PATTERNS/ELINK_DOUTA_0[6]\, C => 
        HIEFFPLA_NET_0_118766, Y => HIEFFPLA_NET_0_118822);
    
    HIEFFPLA_INST_0_57457 : NAND2B
      port map(A => HIEFFPLA_NET_0_116649, B => 
        HIEFFPLA_NET_0_116686, Y => HIEFFPLA_NET_0_116678);
    
    HIEFFPLA_INST_0_58857 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_20[0]\, B => 
        HIEFFPLA_NET_0_116680, S => HIEFFPLA_NET_0_116460, Y => 
        HIEFFPLA_NET_0_116467);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_24[4]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116101, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_8, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_24[4]\);
    
    \U200A_TFC/LOC_STRT_ADDR[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120277, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_4, Q => \U200A_TFC/LOC_STRT_ADDR[5]\);
    
    HIEFFPLA_INST_0_59299 : AND3
      port map(A => HIEFFPLA_NET_0_116620, B => 
        HIEFFPLA_NET_0_117394, C => HIEFFPLA_NET_0_116649, Y => 
        HIEFFPLA_NET_0_116408);
    
    \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM_0[4]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117622, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_22_0, Q => 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM_0[4]_net_1\);
    
    \U_EXEC_MASTER/DEL_CNT[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117790, CLK => CLK_40M_GL, CLR
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i\, Q => 
        \U_EXEC_MASTER/DEL_CNT[5]\);
    
    HIEFFPLA_INST_0_59963 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_4[1]\, B => 
        HIEFFPLA_NET_0_116677, S => HIEFFPLA_NET_0_117155, Y => 
        HIEFFPLA_NET_0_116328);
    
    HIEFFPLA_INST_0_56576 : AND3
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[10]_net_1\, B
         => HIEFFPLA_NET_0_117426, C => HIEFFPLA_NET_0_117425, Y
         => HIEFFPLA_NET_0_116835);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_2[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116752, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_5, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_2[3]\);
    
    HIEFFPLA_INST_0_38795 : MX2
      port map(A => HIEFFPLA_NET_0_119523, B => 
        \U50_PATTERNS/ELINK_ADDRA_13[1]\, S => 
        HIEFFPLA_NET_0_119285, Y => HIEFFPLA_NET_0_120062);
    
    \U50_PATTERNS/ELINK_DINA_18[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119792, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_21, Q => 
        \U50_PATTERNS/ELINK_DINA_18[7]\);
    
    HIEFFPLA_INST_0_46053 : AND3
      port map(A => \U50_PATTERNS/TFC_DOUTA[4]\, B => 
        HIEFFPLA_NET_0_118997, C => HIEFFPLA_NET_0_119365, Y => 
        HIEFFPLA_NET_0_118777);
    
    HIEFFPLA_INST_0_112170 : AO13
      port map(A => HIEFFPLA_NET_0_115817, B => 
        \U200A_TFC/LOC_STOP_ADDR[7]\, C => \TFC_ADDRB[7]\, Y => 
        HIEFFPLA_NET_0_120293);
    
    \U50_PATTERNS/ELINK_DINA_18[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119795, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_21, Q => 
        \U50_PATTERNS/ELINK_DINA_18[4]\);
    
    \U50_PATTERNS/ELINK_DINA_16[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119812, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_18, Q => 
        \U50_PATTERNS/ELINK_DINA_16[3]\);
    
    \U200B_ELINKS/LOC_STRT_ADDR[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120177, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_11, Q => 
        \U200B_ELINKS/LOC_STRT_ADDR[2]\);
    
    HIEFFPLA_INST_0_57169 : AND3
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_2[6]\, B => 
        HIEFFPLA_NET_0_116744, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_2[7]\, Y => 
        HIEFFPLA_NET_0_116726);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_31[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116018, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_10, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_31[2]\);
    
    \U_ELK4_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2\ : IOPADN_BI
      port map(DB => \U_ELK4_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, 
        E => \U_ELK4_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET3\, PAD => 
        ELK4_DAT_N, N2POUT => 
        \U_ELK4_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2_N2P\);
    
    \U50_PATTERNS/U4A_REGCROSS/SAMP_TWO[2]\ : DFN1C0
      port map(D => \U50_PATTERNS/U4A_REGCROSS/SAMP_ONE[2]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_22, Q => 
        \U50_PATTERNS/U4A_REGCROSS/SAMP_TWO[2]_net_1\);
    
    HIEFFPLA_INST_0_56581 : AND3
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[11]_net_1\, B
         => HIEFFPLA_NET_0_117426, C => HIEFFPLA_NET_0_117425, Y
         => HIEFFPLA_NET_0_116834);
    
    HIEFFPLA_INST_0_46204 : AO1
      port map(A => HIEFFPLA_NET_0_119246, B => 
        \U50_PATTERNS/ELINK_DOUTA_3[1]\, C => 
        HIEFFPLA_NET_0_118912, Y => HIEFFPLA_NET_0_118744);
    
    \U_ELK1_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2\ : IOPADN_BI
      port map(DB => \U_ELK1_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, 
        E => \U_ELK1_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET3\, PAD => 
        ELK1_DAT_N, N2POUT => 
        \U_ELK1_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2_N2P\);
    
    \U50_PATTERNS/TFC_DINA[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119196, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_4, Q => \U50_PATTERNS/TFC_DINA[1]\);
    
    HIEFFPLA_INST_0_63069 : AX1
      port map(A => HIEFFPLA_NET_0_115916, B => 
        HIEFFPLA_NET_0_115902, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[11]\, Y => 
        HIEFFPLA_NET_0_115896);
    
    HIEFFPLA_INST_0_47347 : MX2
      port map(A => 
        \U_ELK13_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]_net_1\, B => 
        \U_ELK13_CH/ELK_TX_DAT[6]\, S => 
        \U_ELK13_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118514);
    
    \U_ELK18_CH/U_ELK1_SERDAT_SOURCE/SERDAT[4]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118279, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_13, Q => 
        \U_ELK18_CH/ELK_TX_DAT[4]\);
    
    \U50_PATTERNS/U4E_REGCROSS/LOCAL_REG_VAL_2[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119060, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_1, Q => \OP_MODE_c_2[1]\);
    
    \U50_PATTERNS/ELINK_DINA_10[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119859, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_9, Q => 
        \U50_PATTERNS/ELINK_DINA_10[4]\);
    
    \U_ELK4_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U3\ : IOBI_ID_OD_EB
      port map(DR => \U_ELK4_CH/ELK_OUT_R_i_0\, DF => 
        \U_ELK4_CH/ELK_OUT_F_i_0\, CLR => \GND\, E => 
        \AFLSDF_INV_41\, ICLK => CCC_160M_ADJ, OCLK => 
        CCC_160M_FXD, YIN => 
        \U_ELK4_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\, DOUT => OPEN, 
        EOUT => \U_ELK4_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET3\, YR
         => OPEN, YF => OPEN);
    
    HIEFFPLA_INST_0_43610 : NAND3C
      port map(A => HIEFFPLA_NET_0_119266, B => 
        HIEFFPLA_NET_0_119269, C => HIEFFPLA_NET_0_119252, Y => 
        HIEFFPLA_NET_0_119268);
    
    \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[11]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_115932, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_21, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[11]\);
    
    \U_ELK6_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]\ : DFN1C0
      port map(D => \U_ELK6_CH/U_SLAVE_1ELK/Q[3]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]_net_1\);
    
    \U_ELK6_CH/U_ELK1_SERDAT_SOURCE/SERDAT[5]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117963, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_1, Q => 
        \U_ELK6_CH/ELK_TX_DAT[5]\);
    
    HIEFFPLA_INST_0_54780 : NAND3C
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[1]_net_1\, B => 
        HIEFFPLA_NET_0_117252, C => HIEFFPLA_NET_0_117245, Y => 
        HIEFFPLA_NET_0_117201);
    
    \U_DDR_ELK0/BIBUF_LVDS_0/U0/U2\ : IOPADN_BI
      port map(DB => \U_DDR_ELK0/BIBUF_LVDS_0/U0/NET1\, E => 
        \U_DDR_ELK0/BIBUF_LVDS_0/U0/NET3\, PAD => ELK0_DAT_N, 
        N2POUT => \U_DDR_ELK0/BIBUF_LVDS_0/U0/U2_N2P\);
    
    \U50_PATTERNS/ELINK_DINA_3[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119764, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_11, Q => 
        \U50_PATTERNS/ELINK_DINA_3[3]\);
    
    \U_ELK1_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U3\ : IOBI_ID_OD_EB
      port map(DR => \U_ELK1_CH/ELK_OUT_R_i_0\, DF => 
        \U_ELK1_CH/ELK_OUT_F_i_0\, CLR => \GND\, E => 
        \AFLSDF_INV_35\, ICLK => CCC_160M_ADJ, OCLK => 
        CCC_160M_FXD, YIN => 
        \U_ELK1_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\, DOUT => OPEN, 
        EOUT => \U_ELK1_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET3\, YR
         => OPEN, YF => OPEN);
    
    \U_ELK14_CH/U_SLAVE_1ELK/Q[14]\ : DFN1C0
      port map(D => \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[14]_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/Q[14]_net_1\);
    
    HIEFFPLA_INST_0_55015 : AND3B
      port map(A => HIEFFPLA_NET_0_116768, B => 
        HIEFFPLA_NET_0_117370, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_3[6]_net_1\, Y => 
        HIEFFPLA_NET_0_117140);
    
    \U50_PATTERNS/ELINK_ADDRA_4[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119981, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_2, Q => 
        \U50_PATTERNS/ELINK_ADDRA_4[2]\);
    
    HIEFFPLA_INST_0_49074 : AND2
      port map(A => \U_ELK1_CH/ELK_TX_DAT[0]\, B => 
        \U_ELK1_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118202);
    
    HIEFFPLA_INST_0_55020 : AND3B
      port map(A => HIEFFPLA_NET_0_117339, B => 
        HIEFFPLA_NET_0_117110, C => HIEFFPLA_NET_0_117140, Y => 
        HIEFFPLA_NET_0_117139);
    
    HIEFFPLA_INST_0_40747 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_16[1]\, B => 
        HIEFFPLA_NET_0_119576, S => HIEFFPLA_NET_0_119257, Y => 
        HIEFFPLA_NET_0_119814);
    
    HIEFFPLA_INST_0_52612 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_5[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_6[1]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_2[0]\, Y => 
        HIEFFPLA_NET_0_117539);
    
    HIEFFPLA_INST_0_50519 : MX2
      port map(A => HIEFFPLA_NET_0_117950, B => 
        HIEFFPLA_NET_0_117960, S => \BIT_OS_SEL[0]\, Y => 
        \U_ELK6_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[5]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_6[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116631, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_12, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_6[1]\);
    
    \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[13]\ : DFN1C0
      port map(D => 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[13]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/Q[14]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[14]_net_1\, CLK => 
        CCC_160M_FXD, CLR => P_MASTER_POR_B_c_23, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/Q[14]_net_1\);
    
    \USBCLK60MHZ_pad/U0/U1\ : IOIN_IB
      port map(YIN => \USBCLK60MHZ_pad/U0/NET1\, Y => 
        USBCLK60MHZ_c);
    
    HIEFFPLA_INST_0_53296 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_SEQCNT[4]\, B => 
        HIEFFPLA_NET_0_117433, S => HIEFFPLA_NET_0_117062, Y => 
        HIEFFPLA_NET_0_117438);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_25[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116417, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_20, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_25[3]\);
    
    \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[10]\ : DFN1C0
      port map(D => 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[10]_net_1\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\);
    
    \U_TFC_SERDAT_SOURCE/SERDAT[5]\ : DFN1C0
      port map(D => \U_TFC_SERDAT_SOURCE/N_SERDAT[5]\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \TFC_TX_DAT[5]\);
    
    \U50_PATTERNS/ELINK_ADDRA_13[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120059, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_3, Q => 
        \U50_PATTERNS/ELINK_ADDRA_13[4]\);
    
    \U_ELK11_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U1\ : IOBI_ID_OD_EB
      port map(DR => \U_ELK11_CH/ELK_OUT_R\, DF => 
        \U_ELK11_CH/ELK_OUT_F\, CLR => \GND\, E => 
        \AFLSDF_INV_16\, ICLK => CCC_160M_ADJ, OCLK => 
        CCC_160M_FXD, YIN => 
        \U_ELK11_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\, DOUT => 
        \U_ELK11_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, EOUT => 
        \U_ELK11_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET2\, YR => 
        \U_ELK11_CH/ELK_IN_DDR_R\, YF => 
        \U_ELK11_CH/ELK_IN_DDR_F\);
    
    \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[4]\ : DFN1C0
      port map(D => 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\);
    
    HIEFFPLA_INST_0_45891 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/SM_BANK_SEL[14]\, C => 
        \U50_PATTERNS/ELINK_DOUTA_5[1]\, Y => 
        HIEFFPLA_NET_0_118819);
    
    HIEFFPLA_INST_0_45801 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_12[7]\, C => 
        \U50_PATTERNS/SM_BANK_SEL[7]\, Y => HIEFFPLA_NET_0_118838);
    
    HIEFFPLA_INST_0_47772 : MX2
      port map(A => HIEFFPLA_NET_0_118453, B => 
        HIEFFPLA_NET_0_118450, S => \BIT_OS_SEL_4[0]\, Y => 
        \U_ELK14_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[4]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_SEL_3[1]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_BIT_OS_VAL[1]\, CLK
         => CLK_40M_GL, CLR => P_MASTER_POR_B_c_27_0, Q => 
        \BIT_OS_SEL_3[1]\);
    
    \U62_TS_OE_BUF/_TRIBUFF_F_24U[0]_/U0/U1\ : IOTRI_OB_EB
      port map(D => USB_OE_BI, E => P_USB_MASTER_EN_c, DOUT => 
        \U62_TS_OE_BUF/\\\\TRIBUFF_F_24U[0]\\\\/U0/NET1\, EOUT
         => \U62_TS_OE_BUF/\\\\TRIBUFF_F_24U[0]\\\\/U0/NET2\);
    
    HIEFFPLA_INST_0_44927 : NAND2A
      port map(A => \U50_PATTERNS/USB_RXF_B\, B => 
        \U50_PATTERNS/REG_STATE[3]_net_1\, Y => 
        HIEFFPLA_NET_0_119017);
    
    \DEV_RST_B_pad/U0/U0\ : IOPAD_IN
      port map(PAD => DEV_RST_B, Y => \DEV_RST_B_pad/U0/NET1\);
    
    \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[5]\ : DFN1C0
      port map(D => \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\);
    
    \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[0]\\\\/U0/U0\ : 
        IOPAD_BI_U
      port map(D => 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[0]\\\\/U0/NET1\, 
        E => 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[0]\\\\/U0/NET2\, 
        Y => 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[0]\\\\/U0/NET3\, 
        PAD => BIDIR_USB_ADBUS(0));
    
    HIEFFPLA_INST_0_51671 : XA1
      port map(A => \U_GEN_REF_CLK/GEN_40M_REFCNT[2]_net_1\, B
         => \U_GEN_REF_CLK/GEN_40M_REFCNT[0]_net_1\, C => 
        \U_GEN_REF_CLK/GEN_40M_REFCNT[1]_net_1\, Y => 
        HIEFFPLA_NET_0_117729);
    
    HIEFFPLA_INST_0_48372 : AND2A
      port map(A => \OP_MODE_c_6[1]\, B => \PATT_ELK_DAT_17[6]\, 
        Y => HIEFFPLA_NET_0_118322);
    
    \U_MASTER_DES/U13A_ADJ_160M/SUPDATE/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117614, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_13, Q => \U_MASTER_DES/AUX_SUPDATE\);
    
    HIEFFPLA_INST_0_42029 : AO1A
      port map(A => HIEFFPLA_NET_0_119585, B => 
        HIEFFPLA_NET_0_119579, C => HIEFFPLA_NET_0_119627, Y => 
        HIEFFPLA_NET_0_119628);
    
    \U_MASTER_DES/U13C_MASTER_DESER/BEST_CLKPHASE[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117449, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_10, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_CLKPHASE[3]\);
    
    \U_ELK1_CH/U_SLAVE_1ELK/Q[9]\ : DFN1C0
      port map(D => \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/Q[9]_net_1\);
    
    \U50_PATTERNS/U3_USB_DAT_BUS/_BIBUF_F_24U[3]_/U0/U1\ : 
        IOBI_IRC_OB_EB
      port map(D => \U50_PATTERNS/WR_USB_ADBUS[3]\, CLR => 
        \AFLSDF_INV_7\, E => \U50_PATTERNS/TrienAux\, ICLK => 
        CLK60MHZ, YIN => 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[3]\\\\/U0/NET3\, 
        DOUT => 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[3]\\\\/U0/NET1\, 
        EOUT => 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[3]\\\\/U0/NET2\, 
        Y => \U50_PATTERNS/RD_USB_ADBUS[3]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_26[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116405, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_21, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_26[1]\);
    
    \U_ELK18_CH/U_SLAVE_1ELK/RECD_SER_WORD[0]\ : DFN1C0
      port map(D => \U_ELK18_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[0]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_18[0]\);
    
    \U200B_ELINKS/ADDR_POINTER[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120253, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_31_0, Q => \ELKS_ADDRB[1]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_5[7]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116654, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_11, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_5[7]\);
    
    \U_ELK10_CH/U_SLAVE_1ELK/Q[13]\ : DFN1C0
      port map(D => \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[13]_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/Q[13]_net_1\);
    
    \U_ELK16_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118378, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_10, Q => 
        \U_ELK16_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]_net_1\);
    
    HIEFFPLA_INST_0_45002 : NAND3C
      port map(A => HIEFFPLA_NET_0_119484, B => 
        HIEFFPLA_NET_0_119458, C => HIEFFPLA_NET_0_119002, Y => 
        HIEFFPLA_NET_0_119003);
    
    HIEFFPLA_INST_0_41449 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_6[7]\, B => 
        HIEFFPLA_NET_0_119560, S => HIEFFPLA_NET_0_119258, Y => 
        HIEFFPLA_NET_0_119736);
    
    \U50_PATTERNS/U4A_REGCROSS/SAMP_ONE[0]\ : DFN1C0
      port map(D => \U50_PATTERNS/TFC_STRT_ADDR[0]\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_32, Q => 
        \U50_PATTERNS/U4A_REGCROSS/SAMP_ONE[0]_net_1\);
    
    HIEFFPLA_INST_0_60301 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_9[1]\, B => 
        HIEFFPLA_NET_0_116677, S => HIEFFPLA_NET_0_117130, Y => 
        HIEFFPLA_NET_0_116284);
    
    \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[0]\ : DFN1C0
      port map(D => 
        \U_ELK15_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\);
    
    HIEFFPLA_INST_0_60810 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_15[2]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_16[2]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[0]\, Y => 
        HIEFFPLA_NET_0_116216);
    
    HIEFFPLA_INST_0_51383 : MX2
      port map(A => HIEFFPLA_NET_0_117772, B => 
        \U_EXEC_MASTER/DEL_CNT[6]\, S => HIEFFPLA_NET_0_117796, Y
         => HIEFFPLA_NET_0_117789);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_20[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116464, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_13, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_20[3]\);
    
    HIEFFPLA_INST_0_54729 : AND3B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[2]_net_1\, B => 
        HIEFFPLA_NET_0_117241, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[4]_net_1\, Y => 
        HIEFFPLA_NET_0_117215);
    
    \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[13]\ : DFN1C0
      port map(D => \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\, 
        CLK => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[13]_net_1\);
    
    \U50_PATTERNS/TFC_STOP_ADDR_T[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119174, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_15, Q => 
        \U50_PATTERNS/TFC_STOP_ADDR_T[6]\);
    
    HIEFFPLA_INST_0_61319 : MX2
      port map(A => HIEFFPLA_NET_0_117181, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_21[2]\, S => 
        HIEFFPLA_NET_0_117144, Y => HIEFFPLA_NET_0_116143);
    
    HIEFFPLA_INST_0_42181 : MX2
      port map(A => \U50_PATTERNS/OP_MODE_T[3]\, B => 
        \U50_PATTERNS/RD_USB_ADBUS[3]\, S => 
        HIEFFPLA_NET_0_119440, Y => HIEFFPLA_NET_0_119606);
    
    \U_ELK17_CH/U_ELK1_CMD_TX/SER_OUT_RDEL\ : DFN1C0
      port map(D => \U_ELK17_CH/U_ELK1_CMD_TX/SER_OUT_RI_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_8, Q
         => \U_ELK17_CH/ELK_OUT_R\);
    
    \U50_PATTERNS/SM_BANK_SEL[12]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119319, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_1_0, Q => 
        \U50_PATTERNS/SM_BANK_SEL[12]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_6[4]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116628, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_12, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_6[4]\);
    
    HIEFFPLA_INST_0_49166 : MX2
      port map(A => \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\, B
         => \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\, S => 
        \BIT_OS_SEL[2]\, Y => HIEFFPLA_NET_0_118179);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_4[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116696, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_9, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_4[0]\);
    
    HIEFFPLA_INST_0_57409 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_4[7]\, B => 
        HIEFFPLA_NET_0_116664, S => HIEFFPLA_NET_0_117122, Y => 
        HIEFFPLA_NET_0_116689);
    
    HIEFFPLA_INST_0_56320 : AO1
      port map(A => HIEFFPLA_NET_0_117429, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[3]_net_1\, C => 
        HIEFFPLA_NET_0_116870, Y => HIEFFPLA_NET_0_116894);
    
    \U200A_TFC/RX_SER_WORD_1DEL[2]\ : DFN1C0
      port map(D => \TFC_RX_SER_WORD[2]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_31, Q => 
        \U200A_TFC/RX_SER_WORD_1DEL[2]_net_1\);
    
    HIEFFPLA_INST_0_54093 : MX2
      port map(A => HIEFFPLA_NET_0_116222, B => 
        HIEFFPLA_NET_0_116107, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[3]_net_1\, Y
         => HIEFFPLA_NET_0_117309);
    
    \U_ELK15_CH/U_SLAVE_1ELK/RECD_SER_WORD[2]\ : DFN1C0
      port map(D => \U_ELK15_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[2]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_15[2]\);
    
    HIEFFPLA_INST_0_48941 : MX2
      port map(A => HIEFFPLA_NET_0_118229, B => 
        HIEFFPLA_NET_0_118225, S => \BIT_OS_SEL_0[1]\, Y => 
        HIEFFPLA_NET_0_118221);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_6[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116311, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_2, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_6[3]\);
    
    HIEFFPLA_INST_0_57624 : NAND3B
      port map(A => HIEFFPLA_NET_0_116652, B => 
        HIEFFPLA_NET_0_116646, C => HIEFFPLA_NET_0_116648, Y => 
        HIEFFPLA_NET_0_116649);
    
    HIEFFPLA_INST_0_43085 : NAND2B
      port map(A => HIEFFPLA_NET_0_118994, B => 
        HIEFFPLA_NET_0_119382, Y => HIEFFPLA_NET_0_119383);
    
    HIEFFPLA_INST_0_61784 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_26[2]\, B => 
        HIEFFPLA_NET_0_117131, S => HIEFFPLA_NET_0_117138, Y => 
        HIEFFPLA_NET_0_116078);
    
    \U50_PATTERNS/U4E_REGCROSS/SAMP_TWO[7]\ : DFN1C0
      port map(D => \U50_PATTERNS/U4E_REGCROSS/SAMP_ONE[7]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_24, Q => 
        \U50_PATTERNS/U4E_REGCROSS/SAMP_TWO[7]_net_1\);
    
    HIEFFPLA_INST_0_62215 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_14[3]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_30[3]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[4]_net_1\, Y => 
        HIEFFPLA_NET_0_116021);
    
    HIEFFPLA_INST_0_39902 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_9[4]\, B => 
        HIEFFPLA_NET_0_119519, S => HIEFFPLA_NET_0_119292, Y => 
        HIEFFPLA_NET_0_119939);
    
    \U_ELK18_CH/U_ELK1_CMD_TX/SER_OUT_FDEL\ : DFN1C0
      port map(D => \U_ELK18_CH/U_ELK1_CMD_TX/SER_OUT_FI_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_4, Q
         => \U_ELK18_CH/ELK_OUT_F\);
    
    \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[12]\ : DFN1C0
      port map(D => 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]_net_1\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[12]_net_1\);
    
    HIEFFPLA_INST_0_51991 : MX2A
      port map(A => HIEFFPLA_NET_0_117646, B => 
        HIEFFPLA_NET_0_117645, S => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[1]\, Y => 
        HIEFFPLA_NET_0_117656);
    
    HIEFFPLA_INST_0_60185 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_7[0]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_23[0]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_4[4]_net_1\, Y
         => HIEFFPLA_NET_0_116299);
    
    HIEFFPLA_INST_0_55221 : AOI1D
      port map(A => HIEFFPLA_NET_0_117339, B => 
        HIEFFPLA_NET_0_116812, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[6]_net_1\, Y => 
        HIEFFPLA_NET_0_117082);
    
    HIEFFPLA_INST_0_49090 : MX2
      port map(A => 
        \U_ELK1_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]_net_1\, B => 
        \U_ELK1_CH/ELK_TX_DAT[6]\, S => 
        \U_ELK1_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118199);
    
    \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[9]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_115921, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_9, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[9]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_31[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116342, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_20, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_31[1]\);
    
    \U50_PATTERNS/U4B_REGCROSS/SYNC_SM[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119125, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_23, Q => 
        \U50_PATTERNS/U4B_REGCROSS/SYNC_SM[0]_net_1\);
    
    \U_ELK10_CH/U_SLAVE_1ELK/RECD_SER_WORD[0]\ : DFN1C0
      port map(D => \U_ELK10_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[0]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_10[0]\);
    
    HIEFFPLA_INST_0_56482 : AO1
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[6]_net_1\, B => 
        HIEFFPLA_NET_0_117428, C => HIEFFPLA_NET_0_116838, Y => 
        HIEFFPLA_NET_0_116854);
    
    HIEFFPLA_INST_0_41089 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_1[7]\, B => 
        HIEFFPLA_NET_0_119560, S => HIEFFPLA_NET_0_119243, Y => 
        HIEFFPLA_NET_0_119776);
    
    HIEFFPLA_INST_0_58987 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_22[0]\, B => 
        HIEFFPLA_NET_0_116680, S => HIEFFPLA_NET_0_117095, Y => 
        HIEFFPLA_NET_0_116450);
    
    HIEFFPLA_INST_0_42549 : AND3
      port map(A => HIEFFPLA_NET_0_119371, B => 
        HIEFFPLA_NET_0_119515, C => HIEFFPLA_NET_0_119483, Y => 
        HIEFFPLA_NET_0_119513);
    
    HIEFFPLA_INST_0_41928 : NAND2B
      port map(A => \U50_PATTERNS/ELINK_RWA[13]\, B => 
        HIEFFPLA_NET_0_119657, Y => HIEFFPLA_NET_0_119658);
    
    AFLSDF_INV_11 : INV
      port map(A => P_USB_MASTER_EN_c_22_0, Y => \AFLSDF_INV_11\);
    
    HIEFFPLA_INST_0_61736 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_25[3]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_26[3]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_4[0]\, Y => 
        HIEFFPLA_NET_0_116085);
    
    \U_ELK3_CH/U_ELK1_CMD_TX/SER_OUT_RDEL\ : DFN1P0
      port map(D => \U_ELK3_CH/U_ELK1_CMD_TX/SER_OUT_RI_i\, CLK
         => CCC_160M_FXD, PRE => MASTER_SALT_POR_B_i_0_i_2, Q => 
        \U_ELK3_CH/ELK_OUT_R_i_0\);
    
    \U_ELK16_CH/U_SLAVE_1ELK/Q[9]\ : DFN1C0
      port map(D => \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/Q[9]_net_1\);
    
    HIEFFPLA_INST_0_47117 : MX2
      port map(A => 
        \U_ELK12_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]_net_1\, B => 
        \U_ELK12_CH/ELK_TX_DAT[7]\, S => 
        \U_ELK12_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118555);
    
    HIEFFPLA_INST_0_111788 : MX2C
      port map(A => \U_MASTER_DES/AUX_SDIN\, B => 
        HIEFFPLA_NET_0_117669, S => 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM[2]_net_1\, Y => 
        HIEFFPLA_NET_0_115832);
    
    HIEFFPLA_INST_0_55280 : AND3
      port map(A => HIEFFPLA_NET_0_117119, B => 
        HIEFFPLA_NET_0_117360, C => HIEFFPLA_NET_0_117414, Y => 
        HIEFFPLA_NET_0_117071);
    
    HIEFFPLA_INST_0_55216 : NAND2B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[6]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[8]_net_1\, Y => 
        HIEFFPLA_NET_0_117085);
    
    \U_ELK6_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]\ : DFN1C0
      port map(D => \U_ELK6_CH/U_SLAVE_1ELK/Q[8]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]_net_1\);
    
    HIEFFPLA_INST_0_50286 : MX2
      port map(A => HIEFFPLA_NET_0_118004, B => 
        HIEFFPLA_NET_0_117980, S => \BIT_OS_SEL_0[0]\, Y => 
        \U_ELK5_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[7]\);
    
    \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[8]\ : DFN1C0
      port map(D => \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\);
    
    \U50_PATTERNS/ELINK_ADDRA_7[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119954, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_6, Q => 
        \U50_PATTERNS/ELINK_ADDRA_7[5]\);
    
    \U_ELK2_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]\ : DFN1C0
      port map(D => \U_ELK2_CH/U_SLAVE_1ELK/Q[13]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]_net_1\);
    
    HIEFFPLA_INST_0_40477 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_12[3]\, B => 
        HIEFFPLA_NET_0_119574, S => HIEFFPLA_NET_0_119295, Y => 
        HIEFFPLA_NET_0_119844);
    
    HIEFFPLA_INST_0_37051 : AOI1A
      port map(A => \TFC_STRT_ADDR[5]\, B => 
        HIEFFPLA_NET_0_120349, C => HIEFFPLA_NET_0_120357, Y => 
        HIEFFPLA_NET_0_120358);
    
    HIEFFPLA_INST_0_50080 : MX2
      port map(A => 
        \U_ELK5_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]_net_1\, B => 
        \U_ELK5_CH/ELK_TX_DAT[4]\, S => 
        \U_ELK5_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118020);
    
    \U_ELK7_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]\ : DFN1C0
      port map(D => \U_ELK7_CH/U_SLAVE_1ELK/Q[1]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]_net_1\);
    
    \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[4]\ : DFN1C0
      port map(D => \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\);
    
    HIEFFPLA_INST_0_57268 : NAND2A
      port map(A => HIEFFPLA_NET_0_116713, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_3[0]\, Y => 
        HIEFFPLA_NET_0_116711);
    
    \U50_PATTERNS/U116_PATT_ELINK_BLK/DPRT_512X9_SRAM_R0C0\ : 
        RAM4K9
      generic map(MEMORYFILE => "DPRT_512X9_SRAM_R0C0.mem")

      port map(ADDRA11 => AFLSDF_GND, ADDRA10 => AFLSDF_GND, 
        ADDRA9 => AFLSDF_GND, ADDRA8 => \GND\, ADDRA7 => 
        \U50_PATTERNS/ELINK_ADDRA_16[7]\, ADDRA6 => 
        \U50_PATTERNS/ELINK_ADDRA_16[6]\, ADDRA5 => 
        \U50_PATTERNS/ELINK_ADDRA_16[5]\, ADDRA4 => 
        \U50_PATTERNS/ELINK_ADDRA_16[4]\, ADDRA3 => 
        \U50_PATTERNS/ELINK_ADDRA_16[3]\, ADDRA2 => 
        \U50_PATTERNS/ELINK_ADDRA_16[2]\, ADDRA1 => 
        \U50_PATTERNS/ELINK_ADDRA_16[1]\, ADDRA0 => 
        \U50_PATTERNS/ELINK_ADDRA_16[0]\, ADDRB11 => AFLSDF_GND, 
        ADDRB10 => AFLSDF_GND, ADDRB9 => AFLSDF_GND, ADDRB8 => 
        \GND\, ADDRB7 => \ELKS_ADDRB[7]\, ADDRB6 => 
        \ELKS_ADDRB_0[6]\, ADDRB5 => \ELKS_ADDRB[5]\, ADDRB4 => 
        \ELKS_ADDRB_0[4]\, ADDRB3 => \ELKS_ADDRB[3]\, ADDRB2 => 
        \ELKS_ADDRB_0[2]\, ADDRB1 => \ELKS_ADDRB[1]\, ADDRB0 => 
        \ELKS_ADDRB[0]\, DINA8 => \GND\, DINA7 => 
        \U50_PATTERNS/ELINK_DINA_16[7]\, DINA6 => 
        \U50_PATTERNS/ELINK_DINA_16[6]\, DINA5 => 
        \U50_PATTERNS/ELINK_DINA_16[5]\, DINA4 => 
        \U50_PATTERNS/ELINK_DINA_16[4]\, DINA3 => 
        \U50_PATTERNS/ELINK_DINA_16[3]\, DINA2 => 
        \U50_PATTERNS/ELINK_DINA_16[2]\, DINA1 => 
        \U50_PATTERNS/ELINK_DINA_16[1]\, DINA0 => 
        \U50_PATTERNS/ELINK_DINA_16[0]\, DINB8 => \GND\, DINB7
         => \ELK_RX_SER_WORD_16[7]\, DINB6 => 
        \ELK_RX_SER_WORD_16[6]\, DINB5 => \ELK_RX_SER_WORD_16[5]\, 
        DINB4 => \ELK_RX_SER_WORD_16[4]\, DINB3 => 
        \ELK_RX_SER_WORD_16[3]\, DINB2 => \ELK_RX_SER_WORD_16[2]\, 
        DINB1 => \ELK_RX_SER_WORD_16[1]\, DINB0 => 
        \ELK_RX_SER_WORD_16[0]\, WIDTHA0 => \VCC\, WIDTHA1 => 
        \VCC\, WIDTHB0 => \VCC\, WIDTHB1 => \VCC\, PIPEA => \VCC\, 
        PIPEB => \VCC\, WMODEA => \GND\, WMODEB => \GND\, BLKA
         => \U50_PATTERNS/ELINK_BLKA[16]\, BLKB => 
        ELKS_RAM_BLKB_EN, WENA => \U50_PATTERNS/ELINK_RWA[16]\, 
        WENB => ELKS_RWB, CLKA => CLK60MHZ, CLKB => CLK_40M_GL, 
        RESET => P_USB_MASTER_EN_c_0, DOUTA8 => OPEN, DOUTA7 => 
        \U50_PATTERNS/ELINK_DOUTA_16[7]\, DOUTA6 => 
        \U50_PATTERNS/ELINK_DOUTA_16[6]\, DOUTA5 => 
        \U50_PATTERNS/ELINK_DOUTA_16[5]\, DOUTA4 => 
        \U50_PATTERNS/ELINK_DOUTA_16[4]\, DOUTA3 => 
        \U50_PATTERNS/ELINK_DOUTA_16[3]\, DOUTA2 => 
        \U50_PATTERNS/ELINK_DOUTA_16[2]\, DOUTA1 => 
        \U50_PATTERNS/ELINK_DOUTA_16[1]\, DOUTA0 => 
        \U50_PATTERNS/ELINK_DOUTA_16[0]\, DOUTB8 => OPEN, DOUTB7
         => \PATT_ELK_DAT_16[7]\, DOUTB6 => \PATT_ELK_DAT_16[6]\, 
        DOUTB5 => \PATT_ELK_DAT_16[5]\, DOUTB4 => 
        \PATT_ELK_DAT_16[4]\, DOUTB3 => \PATT_ELK_DAT_16[3]\, 
        DOUTB2 => \PATT_ELK_DAT_16[2]\, DOUTB1 => 
        \PATT_ELK_DAT_16[1]\, DOUTB0 => \PATT_ELK_DAT_16[0]\);
    
    HIEFFPLA_INST_0_37023 : AO1A
      port map(A => \TFC_STRT_ADDR[0]\, B => 
        HIEFFPLA_NET_0_120349, C => HIEFFPLA_NET_0_120348, Y => 
        HIEFFPLA_NET_0_120367);
    
    \U_EXEC_MASTER/MPOR_B_10\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117787, CLK => CLK_40M_GL, CLR
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_1\, Q => 
        P_MASTER_POR_B_c_10);
    
    \U_ELK4_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]\ : DFN1C0
      port map(D => \U_ELK4_CH/U_SLAVE_1ELK/Q[14]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]_net_1\);
    
    HIEFFPLA_INST_0_62674 : XOR2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_SEQCNT[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_CLKPHASE[0]\, Y => 
        HIEFFPLA_NET_0_115959);
    
    HIEFFPLA_INST_0_46607 : MX2
      port map(A => 
        \U_ELK10_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]_net_1\, B => 
        \U_ELK10_CH/ELK_TX_DAT[3]\, S => 
        \U_ELK10_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118647);
    
    HIEFFPLA_INST_0_42313 : AND2A
      port map(A => HIEFFPLA_NET_0_119275, B => 
        \U50_PATTERNS/RD_USB_ADBUS[3]\, Y => 
        HIEFFPLA_NET_0_119574);
    
    \U_ELK10_CH/U_SLAVE_1ELK/Q[9]\ : DFN1C0
      port map(D => \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/Q[9]_net_1\);
    
    HIEFFPLA_INST_0_47630 : MX2
      port map(A => \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[1]_net_1\, 
        B => \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\, S => 
        \BIT_OS_SEL_2[2]\, Y => HIEFFPLA_NET_0_118455);
    
    HIEFFPLA_INST_0_51711 : NAND2B
      port map(A => 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM[4]_net_1\, B => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[34]_net_1\, Y => 
        HIEFFPLA_NET_0_117715);
    
    HIEFFPLA_INST_0_41008 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_19[6]\, B => 
        HIEFFPLA_NET_0_119566, S => HIEFFPLA_NET_0_119293, Y => 
        HIEFFPLA_NET_0_119785);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_14[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116528, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_13, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_14[0]\);
    
    \U_EXEC_MASTER/USB_MASTER_EN/TERMCNT_FG40M0S\ : DFN1C0
      port map(D => 
        \U_EXEC_MASTER/USB_MASTER_EN/TERMCNT_FG60M_net_1\, CLK
         => CLK_40M_GL, CLR => P_MASTER_POR_B_c_32_0, Q => 
        \U_EXEC_MASTER/USB_MASTER_EN/TERMCNT_FG40M0S_net_1\);
    
    \U_ELK15_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]\ : DFN1C0
      port map(D => \U_ELK15_CH/U_SLAVE_1ELK/Q[9]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]_net_1\);
    
    \U50_PATTERNS/ELINK_DINA_0[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119867, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_5, Q => 
        \U50_PATTERNS/ELINK_DINA_0[4]\);
    
    \U_ELK18_CH/U_SLAVE_1ELK/Q[6]\ : DFN1C0
      port map(D => \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/Q[6]_net_1\);
    
    \U_ELK10_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL\ : DFN1C0
      port map(D => 
        \U_ELK10_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL_net_1\);
    
    HIEFFPLA_INST_0_62454 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_5[1]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_6[1]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_2[0]\, Y => 
        HIEFFPLA_NET_0_115987);
    
    \U_ELK2_CH/U_SLAVE_1ELK/Q[3]\ : DFN1C0
      port map(D => \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/Q[3]_net_1\);
    
    HIEFFPLA_INST_0_46566 : MX2
      port map(A => \U_ELK0_CMD_TX/SER_CMD_WORD_R[1]_net_1\, B
         => \ELK0_TX_DAT[5]\, S => 
        \U_ELK0_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118663);
    
    HIEFFPLA_INST_0_44854 : AOI1C
      port map(A => HIEFFPLA_NET_0_119032, B => 
        HIEFFPLA_NET_0_119026, C => HIEFFPLA_NET_0_119034, Y => 
        HIEFFPLA_NET_0_119035);
    
    HIEFFPLA_INST_0_41602 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_9[0]\, B => 
        HIEFFPLA_NET_0_119578, S => HIEFFPLA_NET_0_119292, Y => 
        HIEFFPLA_NET_0_119719);
    
    \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[4]\ : DFN1C0
      port map(D => 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\);
    
    HIEFFPLA_INST_0_61259 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_19[3]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_20[3]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_4[0]\, Y => 
        HIEFFPLA_NET_0_116152);
    
    HIEFFPLA_INST_0_42945 : AO1A
      port map(A => HIEFFPLA_NET_0_119405, B => 
        HIEFFPLA_NET_0_119366, C => HIEFFPLA_NET_0_119397, Y => 
        HIEFFPLA_NET_0_119418);
    
    \U_ELK1_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]\ : DFN1C0
      port map(D => \U_ELK1_CH/U_SLAVE_1ELK/Q[9]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]_net_1\);
    
    HIEFFPLA_INST_0_48371 : AND2A
      port map(A => \OP_MODE_c_6[1]\, B => \PATT_ELK_DAT_17[5]\, 
        Y => HIEFFPLA_NET_0_118323);
    
    HIEFFPLA_INST_0_38146 : MX2
      port map(A => \U50_PATTERNS/CHKSUM[0]\, B => 
        HIEFFPLA_NET_0_120135, S => HIEFFPLA_NET_0_119470, Y => 
        HIEFFPLA_NET_0_120143);
    
    \U_ELK19_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]\ : DFN1C0
      port map(D => \U_ELK19_CH/U_SLAVE_1ELK/Q[2]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]_net_1\);
    
    HIEFFPLA_INST_0_56529 : AND3A
      port map(A => HIEFFPLA_NET_0_117430, B => \BIT_OS_SEL_1[2]\, 
        C => \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[9]_net_1\, 
        Y => HIEFFPLA_NET_0_116845);
    
    HIEFFPLA_INST_0_49119 : AND2A
      port map(A => \OP_MODE_c_5[1]\, B => \PATT_ELK_DAT_1[6]\, Y
         => HIEFFPLA_NET_0_118187);
    
    \U50_PATTERNS/ELINK_DINA_6[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119739, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_16, Q => 
        \U50_PATTERNS/ELINK_DINA_6[4]\);
    
    HIEFFPLA_INST_0_42051 : AND3
      port map(A => \U50_PATTERNS/TFC_DOUTA[7]\, B => 
        HIEFFPLA_NET_0_118997, C => HIEFFPLA_NET_0_119365, Y => 
        HIEFFPLA_NET_0_119623);
    
    HIEFFPLA_INST_0_39966 : MX2
      port map(A => HIEFFPLA_NET_0_119907, B => 
        \U50_PATTERNS/ELINK_BLKA[13]\, S => 
        \U50_PATTERNS/SM_BANK_SEL[20]\, Y => 
        HIEFFPLA_NET_0_119931);
    
    \U_ELK19_CH/U_SLAVE_1ELK/Q[0]\ : DFN1C0
      port map(D => \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/Q[0]_net_1\);
    
    \U50_PATTERNS/U4D_REGCROSS/LOCAL_REG_VAL[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119087, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_3, Q => \ELKS_STOP_ADDR[4]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[5]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_WRD_40M_FIXED[5]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_27, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[5]_net_1\);
    
    HIEFFPLA_INST_0_62209 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_14[2]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_30[2]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[4]_net_1\, Y => 
        HIEFFPLA_NET_0_116022);
    
    \U_ELK18_CH/U_SLAVE_1ELK/RECD_SER_WORD[2]\ : DFN1C0
      port map(D => \U_ELK18_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[2]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_18[2]\);
    
    HIEFFPLA_INST_0_52169 : AO1A
      port map(A => \U_MASTER_DES/CCC2_CONFIG_TRIG\, B => 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM[6]_net_1\, C => 
        HIEFFPLA_NET_0_117625, Y => HIEFFPLA_NET_0_117617);
    
    HIEFFPLA_INST_0_54899 : AO1A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_0[6]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_0[8]_net_1\, C => 
        HIEFFPLA_NET_0_117175, Y => HIEFFPLA_NET_0_117176);
    
    \U_ELK4_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118060, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_17, Q => 
        \U_ELK4_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]_net_1\);
    
    HIEFFPLA_INST_0_50202 : MX2
      port map(A => \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\, B
         => \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[12]_net_1\, S => 
        \BIT_OS_SEL_6[2]\, Y => HIEFFPLA_NET_0_117993);
    
    HIEFFPLA_INST_0_42249 : AND3B
      port map(A => \U50_PATTERNS/RD_USB_ADBUS[4]\, B => 
        HIEFFPLA_NET_0_119590, C => 
        \U50_PATTERNS/RD_USB_ADBUS[5]\, Y => 
        HIEFFPLA_NET_0_119591);
    
    \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[0]\ : DFN1C0
      port map(D => 
        \U_ELK1_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\);
    
    \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[12]\ : DFN1C0
      port map(D => 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]_net_1\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[12]_net_1\);
    
    \U_ELK16_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U0\ : IOPADP_BI
      port map(N2PIN => 
        \U_ELK16_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2_N2P\, D => 
        \U_ELK16_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, E => 
        \U_ELK16_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET2\, PAD => 
        ELK16_DAT_P, Y => 
        \U_ELK16_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\);
    
    \U_GEN_REF_CLK/GEN_40M_REFCNT[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117730, CLK => Y, CLR => 
        DEV_RST_B_c, Q => \U_GEN_REF_CLK/GEN_40M_REFCNT[0]_net_1\);
    
    \U50_PATTERNS/ELINK_DINA_1[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119779, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_7, Q => 
        \U50_PATTERNS/ELINK_DINA_1[4]\);
    
    AFLSDF_INV_45 : INV
      port map(A => DCB_SALT_SEL_c, Y => \AFLSDF_INV_45\);
    
    \U_ELK11_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]\ : DFN1C0
      port map(D => \U_ELK11_CH/U_SLAVE_1ELK/Q[6]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]_net_1\);
    
    HIEFFPLA_INST_0_62845 : AOI1B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[8]_net_1\, B => 
        \OP_MODE_c[5]\, C => HIEFFPLA_NET_0_115942, Y => 
        HIEFFPLA_NET_0_115937);
    
    HIEFFPLA_INST_0_57760 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_6[6]\, B => 
        HIEFFPLA_NET_0_116609, S => HIEFFPLA_NET_0_117599, Y => 
        HIEFFPLA_NET_0_116626);
    
    HIEFFPLA_INST_0_45319 : AO1A
      port map(A => HIEFFPLA_NET_0_118832, B => 
        \U50_PATTERNS/SM_BANK_SEL[7]\, C => HIEFFPLA_NET_0_118941, 
        Y => HIEFFPLA_NET_0_118942);
    
    HIEFFPLA_INST_0_39803 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_8[1]\, B => 
        HIEFFPLA_NET_0_119523, S => HIEFFPLA_NET_0_119291, Y => 
        HIEFFPLA_NET_0_119950);
    
    \U50_PATTERNS/ELINK_DINA_9[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119717, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_19, Q => 
        \U50_PATTERNS/ELINK_DINA_9[2]\);
    
    HIEFFPLA_INST_0_56671 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_0[4]\, B => 
        HIEFFPLA_NET_0_116796, S => HIEFFPLA_NET_0_117602, Y => 
        HIEFFPLA_NET_0_116820);
    
    \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[0]\ : DFN1C0
      port map(D => 
        \U_ELK19_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\);
    
    \U50_PATTERNS/U4C_REGCROSS/DELCNT[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119113, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_28, Q => 
        \U50_PATTERNS/U4C_REGCROSS/DELCNT[0]_net_1\);
    
    HIEFFPLA_INST_0_38777 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_12[7]\, B => 
        HIEFFPLA_NET_0_119516, S => HIEFFPLA_NET_0_119295, Y => 
        HIEFFPLA_NET_0_120064);
    
    HIEFFPLA_INST_0_48053 : MX2
      port map(A => HIEFFPLA_NET_0_118384, B => 
        HIEFFPLA_NET_0_118409, S => \BIT_OS_SEL_2[1]\, Y => 
        HIEFFPLA_NET_0_118386);
    
    HIEFFPLA_INST_0_42007 : NAND3A
      port map(A => HIEFFPLA_NET_0_119450, B => 
        \U50_PATTERNS/REG_STATE_0[1]_net_1\, C => 
        HIEFFPLA_NET_0_119630, Y => HIEFFPLA_NET_0_119633);
    
    HIEFFPLA_INST_0_48911 : MX2
      port map(A => \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\, 
        B => \U_ELK19_CH/U_SLAVE_1ELK/ARB_BYTE[11]_net_1\, S => 
        \BIT_OS_SEL[2]\, Y => HIEFFPLA_NET_0_118225);
    
    \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[12]\ : DFN1C0
      port map(D => \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\);
    
    \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[0]\ : DFN1C0
      port map(D => 
        \U_ELK4_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\);
    
    HIEFFPLA_INST_0_57499 : XA1B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_4[3]\, B => 
        HIEFFPLA_NET_0_116683, C => HIEFFPLA_NET_0_117179, Y => 
        HIEFFPLA_NET_0_116668);
    
    HIEFFPLA_INST_0_37530 : MX2
      port map(A => HIEFFPLA_NET_0_120265, B => TFC_RAM_BLKB_EN, 
        S => HIEFFPLA_NET_0_120264, Y => HIEFFPLA_NET_0_120266);
    
    \U_ELK6_CH/U_SLAVE_1ELK/Q[14]\ : DFN1C0
      port map(D => \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[14]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/Q[14]_net_1\);
    
    \U50_PATTERNS/ELINK_DINA_8[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119724, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_18, Q => 
        \U50_PATTERNS/ELINK_DINA_8[3]\);
    
    HIEFFPLA_INST_0_61973 : MX2
      port map(A => HIEFFPLA_NET_0_117075, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_28[3]\, S => 
        HIEFFPLA_NET_0_117146, Y => HIEFFPLA_NET_0_116052);
    
    HIEFFPLA_INST_0_51426 : XA1
      port map(A => \U_EXEC_MASTER/DEL_CNT[1]\, B => 
        \U_EXEC_MASTER/DEL_CNT[0]\, C => 
        \U_EXEC_MASTER/CCC_1_LOCK_STAT_1D_net_1\, Y => 
        HIEFFPLA_NET_0_117777);
    
    \U_ELK13_CH/U_SLAVE_1ELK/RECD_SER_WORD[0]\ : DFN1C0
      port map(D => \U_ELK13_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[0]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_13[0]\);
    
    \U200B_ELINKS/LOC_STOP_ADDR[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120185, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_7, Q => 
        \U200B_ELINKS/LOC_STOP_ADDR[2]\);
    
    \U_ELK17_CH/U_SLAVE_1ELK/Q[1]\ : DFN1C0
      port map(D => \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/Q[1]_net_1\);
    
    HIEFFPLA_INST_0_55548 : AO1
      port map(A => HIEFFPLA_NET_0_117087, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_1[3]\, C => 
        HIEFFPLA_NET_0_117008, Y => HIEFFPLA_NET_0_117022);
    
    HIEFFPLA_INST_0_54301 : MX2
      port map(A => HIEFFPLA_NET_0_116446, B => 
        HIEFFPLA_NET_0_116523, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_2[3]_net_1\, Y
         => HIEFFPLA_NET_0_117283);
    
    \U50_PATTERNS/ELINK_DINA_11[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119855, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_11, Q => 
        \U50_PATTERNS/ELINK_DINA_11[0]\);
    
    HIEFFPLA_INST_0_40657 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_14[7]\, B => 
        HIEFFPLA_NET_0_119560, S => HIEFFPLA_NET_0_119249, Y => 
        HIEFFPLA_NET_0_119824);
    
    HIEFFPLA_INST_0_37583 : AOI1A
      port map(A => HIEFFPLA_NET_0_120246, B => 
        HIEFFPLA_NET_0_120220, C => HIEFFPLA_NET_0_120254, Y => 
        HIEFFPLA_NET_0_120255);
    
    \U_ELK16_CH/U_SLAVE_1ELK/Q[10]\ : DFN1C0
      port map(D => \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/Q[10]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_0[6]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117099, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_27_1, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_0[6]_net_1\);
    
    \U_ELK12_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]\ : DFN1C0
      port map(D => \U_ELK12_CH/U_SLAVE_1ELK/Q[1]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]_net_1\);
    
    \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[0]\ : DFN1C0
      port map(D => 
        \U_ELK16_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\);
    
    \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[9]\ : DFN1C0
      port map(D => \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\);
    
    HIEFFPLA_INST_0_41116 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_2[2]\, B => 
        HIEFFPLA_NET_0_119575, S => HIEFFPLA_NET_0_119278, Y => 
        HIEFFPLA_NET_0_119773);
    
    \U_ELK13_CH/U_SLAVE_1ELK/RECD_SER_WORD[1]\ : DFN1C0
      port map(D => \U_ELK13_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[1]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_13[1]\);
    
    \U200B_ELINKS/RX_SER_WORD_2DEL[7]\ : DFN1C0
      port map(D => \U200B_ELINKS/RX_SER_WORD_1DEL[7]_net_1\, CLK
         => CLK_40M_GL, CLR => P_MASTER_POR_B_c_26, Q => 
        \U200B_ELINKS/RX_SER_WORD_2DEL[7]_net_1\);
    
    HIEFFPLA_INST_0_42957 : AO1A
      port map(A => HIEFFPLA_NET_0_119388, B => 
        HIEFFPLA_NET_0_118995, C => HIEFFPLA_NET_0_119390, Y => 
        HIEFFPLA_NET_0_119416);
    
    HIEFFPLA_INST_0_39515 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_4[1]\, B => 
        HIEFFPLA_NET_0_119523, S => HIEFFPLA_NET_0_119284, Y => 
        HIEFFPLA_NET_0_119982);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_19[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116178, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_11, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_19[2]\);
    
    HIEFFPLA_INST_0_58085 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_0[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_16[1]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_1[4]_net_1\, Y
         => HIEFFPLA_NET_0_116566);
    
    HIEFFPLA_INST_0_54776 : NAND3B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[4]_net_1\, B => 
        HIEFFPLA_NET_0_117241, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[2]_net_1\, Y => 
        HIEFFPLA_NET_0_117202);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_1[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116786, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_4, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_1[2]\);
    
    \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[11]\ : DFN1C0
      port map(D => \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\);
    
    \U_ELK12_CH/U_SLAVE_1ELK/RECD_SER_WORD[4]\ : DFN1C0
      port map(D => \U_ELK12_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[4]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_12[4]\);
    
    \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[10]\ : DFN1C0
      port map(D => \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\);
    
    HIEFFPLA_INST_0_57552 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_5[2]\, B => 
        HIEFFPLA_NET_0_116643, S => HIEFFPLA_NET_0_117121, Y => 
        HIEFFPLA_NET_0_116659);
    
    HIEFFPLA_INST_0_51498 : NAND3
      port map(A => \U_EXEC_MASTER/PRESCALE[2]\, B => 
        \U_EXEC_MASTER/PRESCALE[3]\, C => 
        \U_EXEC_MASTER/PRESCALE[1]\, Y => HIEFFPLA_NET_0_117764);
    
    \U_ELK3_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]\ : DFN1C0
      port map(D => \U_ELK3_CH/U_SLAVE_1ELK/Q[5]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]_net_1\);
    
    HIEFFPLA_INST_0_39443 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_3[1]\, B => 
        HIEFFPLA_NET_0_119523, S => HIEFFPLA_NET_0_119247, Y => 
        HIEFFPLA_NET_0_119990);
    
    \U_EXEC_MASTER/MPOR_B_9\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117787, CLK => CLK_40M_GL, CLR
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_1\, Q => 
        P_MASTER_POR_B_c_9);
    
    \U50_PATTERNS/ELINK_ADDRA_10[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120083, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_22, Q => 
        \U50_PATTERNS/ELINK_ADDRA_10[4]\);
    
    \U_ELK15_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]\ : DFN1C0
      port map(D => \U_ELK15_CH/U_SLAVE_1ELK/Q[1]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]_net_1\);
    
    HIEFFPLA_INST_0_59552 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_12[3]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_28[3]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[4]_net_1\, Y
         => HIEFFPLA_NET_0_116379);
    
    HIEFFPLA_INST_0_55818 : MX2
      port map(A => HIEFFPLA_NET_0_116146, B => 
        HIEFFPLA_NET_0_116060, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[3]\, Y => 
        HIEFFPLA_NET_0_116986);
    
    HIEFFPLA_INST_0_48503 : MX2
      port map(A => HIEFFPLA_NET_0_118306, B => 
        HIEFFPLA_NET_0_118320, S => \BIT_OS_SEL_3[0]\, Y => 
        \U_ELK17_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[2]\);
    
    \U_ELK17_CH/U_SLAVE_1ELK/Q[2]\ : DFN1C0
      port map(D => \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/Q[2]_net_1\);
    
    HIEFFPLA_INST_0_49234 : MX2
      port map(A => HIEFFPLA_NET_0_118161, B => 
        HIEFFPLA_NET_0_118172, S => \BIT_OS_SEL_1[0]\, Y => 
        \U_ELK1_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[0]\);
    
    HIEFFPLA_INST_0_44442 : XOR2
      port map(A => \U50_PATTERNS/U4B_REGCROSS/DELCNT[0]_net_1\, 
        B => \U50_PATTERNS/U4B_REGCROSS/DELCNT[1]_net_1\, Y => 
        HIEFFPLA_NET_0_119115);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_9[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116284, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_6, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_9[1]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/MAX_CNT[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_116950, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_16, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/MAX_CNT[4]\);
    
    \U_ELK1_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118202, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_7, Q => 
        \U_ELK1_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]_net_1\);
    
    HIEFFPLA_INST_0_59125 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_24[2]\, B => 
        HIEFFPLA_NET_0_116428, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_2[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116432);
    
    HIEFFPLA_INST_0_52409 : MX2
      port map(A => HIEFFPLA_NET_0_117519, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_29[1]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[3]\, Y => 
        HIEFFPLA_NET_0_117567);
    
    \U_ELK14_CH/U_SLAVE_1ELK/Q[7]\ : DFN1C0
      port map(D => \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/Q[7]_net_1\);
    
    \U50_PATTERNS/ELINK_ADDRA_11[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120076, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_2, Q => 
        \U50_PATTERNS/ELINK_ADDRA_11[3]\);
    
    \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[79]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117702, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_34, Q => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[79]_net_1\);
    
    HIEFFPLA_INST_0_53086 : MX2
      port map(A => HIEFFPLA_NET_0_117555, B => 
        HIEFFPLA_NET_0_117551, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[2]\, Y => 
        HIEFFPLA_NET_0_117467);
    
    HIEFFPLA_INST_0_48863 : AND2
      port map(A => CLK_40M_GL, B => 
        \U_ELK19_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0_net_1\, Y => 
        HIEFFPLA_NET_0_118239);
    
    \U50_PATTERNS/ELINKS_STRT_ADDR_T[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120103, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_21, Q => 
        \U50_PATTERNS/ELINKS_STRT_ADDR_T[0]\);
    
    HIEFFPLA_INST_0_57514 : XA1B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_4[6]\, B => 
        HIEFFPLA_NET_0_116672, C => HIEFFPLA_NET_0_117179, Y => 
        HIEFFPLA_NET_0_116665);
    
    HIEFFPLA_INST_0_55293 : AOI1A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[6]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[8]_net_1\, C => 
        HIEFFPLA_NET_0_117393, Y => HIEFFPLA_NET_0_117069);
    
    HIEFFPLA_INST_0_40076 : AOI1A
      port map(A => \U50_PATTERNS/ELINK_BLKA[0]\, B => 
        HIEFFPLA_NET_0_119664, C => HIEFFPLA_NET_0_119914, Y => 
        HIEFFPLA_NET_0_119915);
    
    HIEFFPLA_INST_0_55203 : AND3A
      port map(A => HIEFFPLA_NET_0_117247, B => 
        HIEFFPLA_NET_0_117240, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[6]_net_1\, Y => 
        HIEFFPLA_NET_0_117093);
    
    HIEFFPLA_INST_0_52734 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_21[0]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_22[0]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[0]\, Y => 
        HIEFFPLA_NET_0_117520);
    
    HIEFFPLA_INST_0_42768 : AO1D
      port map(A => \U50_PATTERNS/REG_STATE_0[1]_net_1\, B => 
        HIEFFPLA_NET_0_119366, C => HIEFFPLA_NET_0_119425, Y => 
        HIEFFPLA_NET_0_119466);
    
    \U_ELK19_CH/U_SLAVE_1ELK/Q[13]\ : DFN1C0
      port map(D => \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[13]_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/Q[13]_net_1\);
    
    \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[13]\ : DFN1C0
      port map(D => 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[13]_net_1\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[13]_net_1\);
    
    HIEFFPLA_INST_0_111268 : AND3A
      port map(A => HIEFFPLA_NET_0_115845, B => 
        HIEFFPLA_NET_0_116344, C => HIEFFPLA_NET_0_117357, Y => 
        HIEFFPLA_NET_0_116347);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_2[5]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116750, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_5, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_2[5]\);
    
    \U_ELK1_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118196, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_4, Q => 
        \U_ELK1_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]_net_1\);
    
    \U50_PATTERNS/U4D_REGCROSS/SYNC_SM[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119083, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_25, Q => 
        \U50_PATTERNS/U4D_REGCROSS/SYNC_SM[0]_net_1\);
    
    HIEFFPLA_INST_0_44150 : MX2
      port map(A => \U50_PATTERNS/TFC_STRT_ADDR[5]\, B => 
        \U50_PATTERNS/TFC_STRT_ADDR_T[5]\, S => 
        HIEFFPLA_NET_0_119472, Y => HIEFFPLA_NET_0_119167);
    
    HIEFFPLA_INST_0_52624 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_5[3]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_6[3]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_2[0]\, Y => 
        HIEFFPLA_NET_0_117537);
    
    \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[6]\ : DFN1C0
      port map(D => 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\);
    
    HIEFFPLA_INST_0_49804 : MX2
      port map(A => HIEFFPLA_NET_0_118085, B => 
        HIEFFPLA_NET_0_118068, S => \BIT_OS_SEL_0[1]\, Y => 
        HIEFFPLA_NET_0_118070);
    
    HIEFFPLA_INST_0_48324 : MX2
      port map(A => \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\, 
        B => \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[14]_net_1\, S => 
        \BIT_OS_SEL_3[2]\, Y => HIEFFPLA_NET_0_118338);
    
    \U_ELK3_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]\ : DFN1C0
      port map(D => \U_ELK3_CH/U_SLAVE_1ELK/Q[11]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]_net_1\);
    
    HIEFFPLA_INST_0_48605 : MX2
      port map(A => 
        \U_ELK18_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]_net_1\, B => 
        \U_ELK18_CH/ELK_TX_DAT[5]\, S => 
        \U_ELK18_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118286);
    
    HIEFFPLA_INST_0_44070 : MX2
      port map(A => \U50_PATTERNS/TFC_STOP_ADDR_T[3]\, B => 
        \U50_PATTERNS/RD_USB_ADBUS[3]\, S => 
        HIEFFPLA_NET_0_119492, Y => HIEFFPLA_NET_0_119177);
    
    HIEFFPLA_INST_0_41170 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_3[0]\, B => 
        HIEFFPLA_NET_0_119578, S => HIEFFPLA_NET_0_119247, Y => 
        HIEFFPLA_NET_0_119767);
    
    \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[12]\ : DFN1C0
      port map(D => 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[12]_net_1\);
    
    \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[3]\ : DFN1C0
      port map(D => 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[3]_net_1\);
    
    HIEFFPLA_INST_0_55332 : AOI1C
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[5]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[3]_net_1\, C => 
        HIEFFPLA_NET_0_117053, Y => HIEFFPLA_NET_0_117058);
    
    HIEFFPLA_INST_0_52842 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_15[2]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_16[2]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_2[0]\, Y => 
        HIEFFPLA_NET_0_117502);
    
    \U_MASTER_DES/U13C_MASTER_DESER/BEST_SEQCNT[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117439, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_9, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_SEQCNT[3]\);
    
    HIEFFPLA_INST_0_46584 : AND2
      port map(A => \U_ELK10_CH/ELK_TX_DAT[0]\, B => 
        \U_ELK10_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118652);
    
    HIEFFPLA_INST_0_54877 : NAND3B
      port map(A => HIEFFPLA_NET_0_117139, B => 
        HIEFFPLA_NET_0_117069, C => HIEFFPLA_NET_0_117179, Y => 
        HIEFFPLA_NET_0_117183);
    
    \U_ELK11_CH/U_SLAVE_1ELK/Q[2]\ : DFN1C0
      port map(D => \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/Q[2]_net_1\);
    
    \U_ELK13_CH/U_ELK1_CMD_TX/SER_OUT_RI\ : DFN1C0
      port map(D => 
        \U_ELK13_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[3]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_1, Q => 
        \U_ELK13_CH/U_ELK1_CMD_TX/SER_OUT_RI_net_1\);
    
    HIEFFPLA_INST_0_62442 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_5[4]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_6[4]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_2[0]\, Y => 
        HIEFFPLA_NET_0_115989);
    
    HIEFFPLA_INST_0_62289 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_3[2]\, 
        B => HIEFFPLA_NET_0_117131, S => HIEFFPLA_NET_0_117178, Y
         => HIEFFPLA_NET_0_116008);
    
    HIEFFPLA_INST_0_62493 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_6[3]\, 
        B => HIEFFPLA_NET_0_117075, S => HIEFFPLA_NET_0_117132, Y
         => HIEFFPLA_NET_0_115982);
    
    HIEFFPLA_INST_0_44736 : MX2
      port map(A => \OP_MODE_c_3[1]\, B => 
        \U50_PATTERNS/U4E_REGCROSS/SAMP_TWO[1]_net_1\, S => 
        HIEFFPLA_NET_0_119072, Y => HIEFFPLA_NET_0_119059);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_21[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116453, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_14, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_21[3]\);
    
    HIEFFPLA_INST_0_54684 : MX2
      port map(A => HIEFFPLA_NET_0_117297, B => 
        HIEFFPLA_NET_0_117279, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[2]_net_1\, Y => 
        HIEFFPLA_NET_0_117223);
    
    HIEFFPLA_INST_0_48576 : AND2
      port map(A => \U_ELK18_CH/ELK_TX_DAT[0]\, B => 
        \U_ELK18_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118292);
    
    \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[11]\ : DFN1C0
      port map(D => 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]_net_1\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[11]_net_1\);
    
    \U50_PATTERNS/OP_MODE_T[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119605, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_17, Q => 
        \U50_PATTERNS/OP_MODE_T[4]\);
    
    HIEFFPLA_INST_0_50338 : AND2
      port map(A => \U_ELK6_CH/ELK_TX_DAT[1]\, B => 
        \U_ELK6_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_117973);
    
    HIEFFPLA_INST_0_49748 : MX2
      port map(A => HIEFFPLA_NET_0_118081, B => 
        HIEFFPLA_NET_0_118080, S => \BIT_OS_SEL_1[0]\, Y => 
        \U_ELK3_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[2]\);
    
    HIEFFPLA_INST_0_37287 : NAND3C
      port map(A => \U200A_TFC/GP_PG_SM[6]_net_1\, B => 
        \U200A_TFC/GP_PG_SM[7]_net_1\, C => \OP_MODE[0]\, Y => 
        HIEFFPLA_NET_0_120305);
    
    \U_EXEC_MASTER/MPOR_B_29\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117787, CLK => CLK_40M_GL, CLR
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_0\, Q => 
        P_MASTER_POR_B_c_29);
    
    HIEFFPLA_INST_0_40468 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_12[2]\, B => 
        HIEFFPLA_NET_0_119575, S => HIEFFPLA_NET_0_119295, Y => 
        HIEFFPLA_NET_0_119845);
    
    HIEFFPLA_INST_0_48278 : MX2
      port map(A => HIEFFPLA_NET_0_118359, B => 
        HIEFFPLA_NET_0_118354, S => \BIT_OS_SEL_3[0]\, Y => 
        \U_ELK16_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[5]\);
    
    \U50_PATTERNS/ELINK_DINA_19[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119788, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_1, Q => 
        \U50_PATTERNS/ELINK_DINA_19[3]\);
    
    HIEFFPLA_INST_0_56242 : AND2
      port map(A => DCB_SALT_SEL_c, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/RECD_SER_WORD[4]_net_1\, 
        Y => \ELK_RX_SER_WORD_0[4]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_12[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116254, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_21, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_12[1]\);
    
    \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[4]\ : DFN1C0
      port map(D => 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\);
    
    HIEFFPLA_INST_0_55675 : MX2
      port map(A => HIEFFPLA_NET_0_115989, B => 
        HIEFFPLA_NET_0_116245, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_2[3]\, Y => 
        HIEFFPLA_NET_0_117005);
    
    HIEFFPLA_INST_0_46419 : NOR3A
      port map(A => \U50_PATTERNS/WR_XFER_TYPE[0]_net_1\, B => 
        HIEFFPLA_NET_0_118692, C => 
        \U50_PATTERNS/WR_XFER_TYPE[1]_net_1\, Y => 
        HIEFFPLA_NET_0_118694);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_6[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116312, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_2, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_6[2]\);
    
    \U_ELK5_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]\ : DFN1C0
      port map(D => \U_ELK5_CH/U_SLAVE_1ELK/Q[8]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_29[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116045, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_16_0, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_29[0]\);
    
    \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_40M\ : DFN1C0
      port map(D => 
        \U_EXEC_MASTER/USB_MASTER_EN/TEST_SM[4]_net_1\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_29, Q => 
        \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_40M_net_1\);
    
    \U50_PATTERNS/U3_USB_DAT_BUS/_BIBUF_F_24U[5]_/U0/U1\ : 
        IOBI_IRC_OB_EB
      port map(D => \U50_PATTERNS/WR_USB_ADBUS[5]\, CLR => 
        \AFLSDF_INV_9\, E => \U50_PATTERNS/TrienAux\, ICLK => 
        CLK60MHZ, YIN => 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[5]\\\\/U0/NET3\, 
        DOUT => 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[5]\\\\/U0/NET1\, 
        EOUT => 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[5]\\\\/U0/NET2\, 
        Y => \U50_PATTERNS/RD_USB_ADBUS[5]\);
    
    HIEFFPLA_INST_0_46874 : NAND2B
      port map(A => \OP_MODE_c[1]\, B => \PATT_ELK_DAT_11[2]\, Y
         => HIEFFPLA_NET_0_118596);
    
    HIEFFPLA_INST_0_42727 : AND3B
      port map(A => HIEFFPLA_NET_0_119379, B => 
        \U50_PATTERNS/REG_STATE_0[2]_net_1\, C => 
        HIEFFPLA_NET_0_119431, Y => HIEFFPLA_NET_0_119474);
    
    HIEFFPLA_INST_0_38876 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_14[2]\, B => 
        HIEFFPLA_NET_0_119522, S => HIEFFPLA_NET_0_119249, Y => 
        HIEFFPLA_NET_0_120053);
    
    \U_ELK14_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118469, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_5, Q => 
        \U_ELK14_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]_net_1\);
    
    \U_ELK7_CH/U_ELK1_SERDAT_SOURCE/SERDAT[7]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117916, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_3, Q => 
        \U_ELK7_CH/ELK_TX_DAT[7]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_3[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116336, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_19, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_3[3]\);
    
    HIEFFPLA_INST_0_51684 : MX2
      port map(A => \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[47]\, B
         => \U_MASTER_DES/PHASE_ADJ_160_L[1]\, S => 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM_0[4]_net_1\, Y => 
        HIEFFPLA_NET_0_117725);
    
    HIEFFPLA_INST_0_41978 : NAND2B
      port map(A => \U50_PATTERNS/ELINK_RWA[8]\, B => 
        HIEFFPLA_NET_0_119638, Y => HIEFFPLA_NET_0_119639);
    
    HIEFFPLA_INST_0_60171 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_7[2]\, B => 
        HIEFFPLA_NET_0_116295, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_0[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116301);
    
    \U50_PATTERNS/USB_SIWU_BI/U1\ : DFN1P0
      port map(D => HIEFFPLA_NET_0_119013, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_8, Q => USB_SIWU_BI);
    
    HIEFFPLA_INST_0_49220 : MX2
      port map(A => \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\, B
         => \U_ELK1_CH/U_SLAVE_1ELK/ARB_BYTE[13]_net_1\, S => 
        \BIT_OS_SEL[2]\, Y => HIEFFPLA_NET_0_118171);
    
    \U0A_40M_REFCLK/_BIBUF_LVDS[0]_/U0/U1\ : IOBI_IB_OB_EB
      port map(D => CLK40M_10NS_REF, E => \AFLSDF_INV_2\, YIN => 
        \U0A_40M_REFCLK/\\\\BIBUF_LVDS[0]\\\\/U0/NET4\, DOUT => 
        \U0A_40M_REFCLK/\\\\BIBUF_LVDS[0]\\\\/U0/NET1\, EOUT => 
        \U0A_40M_REFCLK/\\\\BIBUF_LVDS[0]\\\\/U0/NET2\, Y => 
        CLK_40M_BUF_RECD);
    
    HIEFFPLA_INST_0_49093 : AND2
      port map(A => HIEFFPLA_NET_0_161288, B => 
        HIEFFPLA_NET_0_161287, Y => HIEFFPLA_NET_0_118198);
    
    HIEFFPLA_INST_0_39596 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_5[2]\, B => 
        HIEFFPLA_NET_0_119522, S => HIEFFPLA_NET_0_119251, Y => 
        HIEFFPLA_NET_0_119973);
    
    HIEFFPLA_INST_0_37297 : AOI1B
      port map(A => \OP_MODE[0]\, B => 
        \U200A_TFC/GP_PG_SM[6]_net_1\, C => HIEFFPLA_NET_0_120295, 
        Y => HIEFFPLA_NET_0_120301);
    
    \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[13]\ : DFN1C0
      port map(D => \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[11]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[13]_net_1\);
    
    \U_ELK18_CH/U_SLAVE_1ELK/Q[3]\ : DFN1C0
      port map(D => \U_ELK18_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/Q[3]_net_1\);
    
    HIEFFPLA_INST_0_40873 : MX2
      port map(A => HIEFFPLA_NET_0_119560, B => 
        \U50_PATTERNS/ELINK_DINA_17[7]\, S => 
        HIEFFPLA_NET_0_119260, Y => HIEFFPLA_NET_0_119800);
    
    HIEFFPLA_INST_0_48367 : NAND2B
      port map(A => \OP_MODE_c_6[1]\, B => \PATT_ELK_DAT_17[1]\, 
        Y => HIEFFPLA_NET_0_118327);
    
    \U_ELK16_CH/U_ELK1_SERDAT_SOURCE/SERDAT[4]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118369, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_9, Q => 
        \U_ELK16_CH/ELK_TX_DAT[4]\);
    
    HIEFFPLA_INST_0_48535 : MX2
      port map(A => HIEFFPLA_NET_0_118308, B => 
        HIEFFPLA_NET_0_118305, S => \BIT_OS_SEL_3[0]\, Y => 
        \U_ELK17_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[6]\);
    
    HIEFFPLA_INST_0_43765 : AND3B
      port map(A => \U50_PATTERNS/RD_USB_ADBUS[3]\, B => 
        \U50_PATTERNS/RD_USB_ADBUS[2]\, C => 
        HIEFFPLA_NET_0_119593, Y => HIEFFPLA_NET_0_119219);
    
    \U50_PATTERNS/U4C_REGCROSS/SAMP_ONE[4]\ : DFN1C0
      port map(D => \U50_PATTERNS/ELINKS_STRT_ADDR[4]\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_33, Q => 
        \U50_PATTERNS/U4C_REGCROSS/SAMP_ONE[4]_net_1\);
    
    HIEFFPLA_INST_0_56934 : NAND2B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_1[4]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_1[5]\, Y => 
        HIEFFPLA_NET_0_116771);
    
    HIEFFPLA_INST_0_60612 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_13[0]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_29[0]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_2[4]_net_1\, Y
         => HIEFFPLA_NET_0_116244);
    
    HIEFFPLA_INST_0_47945 : MX2
      port map(A => HIEFFPLA_NET_0_118403, B => 
        HIEFFPLA_NET_0_118398, S => \BIT_OS_SEL_2[1]\, Y => 
        HIEFFPLA_NET_0_118400);
    
    HIEFFPLA_INST_0_49186 : MX2
      port map(A => HIEFFPLA_NET_0_118178, B => 
        HIEFFPLA_NET_0_118174, S => \BIT_OS_SEL_0[1]\, Y => 
        HIEFFPLA_NET_0_118176);
    
    HIEFFPLA_INST_0_47874 : AND2A
      port map(A => \OP_MODE_c_6[1]\, B => \PATT_ELK_DAT_15[6]\, 
        Y => HIEFFPLA_NET_0_118412);
    
    HIEFFPLA_INST_0_42629 : AO1
      port map(A => HIEFFPLA_NET_0_119557, B => 
        HIEFFPLA_NET_0_119465, C => HIEFFPLA_NET_0_119481, Y => 
        HIEFFPLA_NET_0_119496);
    
    \U_ELK3_CH/U_SLAVE_1ELK/Q[5]\ : DFN1C0
      port map(D => \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/Q[5]_net_1\);
    
    \U_ELK2_CH/U_SLAVE_1ELK/Q[6]\ : DFN1C0
      port map(D => \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/Q[6]_net_1\);
    
    \U_ELK14_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]\ : DFN1C0
      port map(D => \U_ELK14_CH/U_SLAVE_1ELK/Q[0]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[0]_net_1\);
    
    HIEFFPLA_INST_0_63144 : AX1C
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[2]_net_1\, B => 
        HIEFFPLA_NET_0_115876, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[3]_net_1\, Y => 
        HIEFFPLA_NET_0_115877);
    
    \U_EXEC_MASTER/MPOR_SALT_B_7\ : DFI1P0
      port map(D => HIEFFPLA_NET_0_117781, CLK => CLK_40M_GL, PRE
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_2\, QN => 
        MASTER_SALT_POR_B_i_0_i_7);
    
    HIEFFPLA_INST_0_39101 : MX2
      port map(A => HIEFFPLA_NET_0_119520, B => 
        \U50_PATTERNS/ELINK_ADDRA_17[3]\, S => 
        HIEFFPLA_NET_0_119260, Y => HIEFFPLA_NET_0_120028);
    
    HIEFFPLA_INST_0_43332 : XA1C
      port map(A => HIEFFPLA_NET_0_119330, B => 
        \U50_PATTERNS/SI_CNT[3]\, C => HIEFFPLA_NET_0_119452, Y
         => HIEFFPLA_NET_0_119324);
    
    HIEFFPLA_INST_0_51949 : MX2A
      port map(A => HIEFFPLA_NET_0_117652, B => 
        HIEFFPLA_NET_0_117651, S => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[6]\, Y => 
        HIEFFPLA_NET_0_117660);
    
    HIEFFPLA_INST_0_44710 : MX2
      port map(A => \U50_PATTERNS/U4E_REGCROSS/LOCAL_REG_VAL[7]\, 
        B => \U50_PATTERNS/U4E_REGCROSS/SAMP_TWO[7]_net_1\, S => 
        HIEFFPLA_NET_0_119072, Y => HIEFFPLA_NET_0_119063);
    
    \U_ELK14_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118471, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_5, Q => 
        \U_ELK14_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/TUNE_CLKPHASE[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_115948, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_12, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/TUNE_CLKPHASE[1]\);
    
    \U_ELK2_CH/U_SLAVE_1ELK/Q[14]\ : DFN1C0
      port map(D => \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[14]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/Q[14]_net_1\);
    
    HIEFFPLA_INST_0_56155 : NAND2A
      port map(A => HIEFFPLA_NET_0_116941, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/MAX_CNT[4]\, Y => 
        HIEFFPLA_NET_0_116940);
    
    HIEFFPLA_INST_0_53688 : MX2
      port map(A => HIEFFPLA_NET_0_117322, B => 
        HIEFFPLA_NET_0_117267, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[1]_net_1\, Y
         => HIEFFPLA_NET_0_117372);
    
    HIEFFPLA_INST_0_42896 : NAND2
      port map(A => \U50_PATTERNS/REG_STATE[5]_net_1\, B => 
        \U50_PATTERNS/REG_STATE[2]_net_1\, Y => 
        HIEFFPLA_NET_0_119432);
    
    HIEFFPLA_INST_0_53306 : AND2A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_0[8]_net_1\, B => 
        HIEFFPLA_NET_0_116977, Y => HIEFFPLA_NET_0_117435);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_7[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116602, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_14, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_7[1]\);
    
    HIEFFPLA_INST_0_55965 : MX2
      port map(A => HIEFFPLA_NET_0_116985, B => 
        HIEFFPLA_NET_0_116969, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[4]\, Y => 
        HIEFFPLA_NET_0_116967);
    
    \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_2S_5\ : DFN1C0
      port map(D => 
        \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_1S_net_1\, CLK
         => CLK60MHZ, CLR => P_MASTER_POR_B_c_0_0, Q => 
        P_USB_MASTER_EN_c_5);
    
    \U_ELK1_CH/U_ELK1_SERDAT_SOURCE/SERDAT[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118192, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_11, Q => 
        \U_ELK1_CH/ELK_TX_DAT[1]\);
    
    \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[1]\ : DFN1C0
      port map(D => 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[1]_net_1\);
    
    HIEFFPLA_INST_0_61457 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_6[2]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_22[2]\, S
         => \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_5[4]_net_1\, 
        Y => HIEFFPLA_NET_0_116124);
    
    HIEFFPLA_INST_0_38298 : MX2
      port map(A => \U50_PATTERNS/ELINKS_STOP_ADDR[7]\, B => 
        \U50_PATTERNS/ELINKS_STOP_ADDR_T[7]\, S => 
        HIEFFPLA_NET_0_119472, Y => HIEFFPLA_NET_0_120120);
    
    HIEFFPLA_INST_0_53412 : MX2
      port map(A => HIEFFPLA_NET_0_117199, B => 
        HIEFFPLA_NET_0_117346, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[2]_net_1\, Y
         => HIEFFPLA_NET_0_117412);
    
    \U50_PATTERNS/ELINK_DINA_16[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119809, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_18, Q => 
        \U50_PATTERNS/ELINK_DINA_16[6]\);
    
    HIEFFPLA_INST_0_59268 : AO1
      port map(A => HIEFFPLA_NET_0_116589, B => 
        HIEFFPLA_NET_0_117394, C => HIEFFPLA_NET_0_116408, Y => 
        HIEFFPLA_NET_0_116411);
    
    HIEFFPLA_INST_0_40531 : MX2
      port map(A => HIEFFPLA_NET_0_119576, B => 
        \U50_PATTERNS/ELINK_DINA_13[1]\, S => 
        HIEFFPLA_NET_0_119285, Y => HIEFFPLA_NET_0_119838);
    
    \U_ELK8_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117884, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]_net_1\);
    
    \U_ELK5_CH/U_SLAVE_1ELK/Q[8]\ : DFN1C0
      port map(D => \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/Q[8]_net_1\);
    
    HIEFFPLA_INST_0_37190 : NAND2B
      port map(A => \U200A_TFC/GP_PG_SM[2]_net_1\, B => 
        \U200A_TFC/GP_PG_SM[3]_net_1\, Y => HIEFFPLA_NET_0_120328);
    
    HIEFFPLA_INST_0_37952 : MX2
      port map(A => \U200B_ELINKS/LOC_STOP_ADDR[3]\, B => 
        \ELKS_STOP_ADDR[3]\, S => 
        \U200B_ELINKS/GP_PG_SM_0[10]_net_1\, Y => 
        HIEFFPLA_NET_0_120184);
    
    HIEFFPLA_INST_0_62009 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_12[3]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_28[3]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_3[4]_net_1\, Y
         => HIEFFPLA_NET_0_116047);
    
    HIEFFPLA_INST_0_41458 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_7[0]\, B => 
        HIEFFPLA_NET_0_119578, S => HIEFFPLA_NET_0_119289, Y => 
        HIEFFPLA_NET_0_119735);
    
    HIEFFPLA_INST_0_44166 : MX2
      port map(A => \U50_PATTERNS/TFC_STRT_ADDR[7]\, B => 
        \U50_PATTERNS/TFC_STRT_ADDR_T[7]\, S => 
        HIEFFPLA_NET_0_119472, Y => HIEFFPLA_NET_0_119165);
    
    HIEFFPLA_INST_0_43249 : AND2A
      port map(A => \U50_PATTERNS/RD_XFER_TYPE[0]_net_1\, B => 
        \U50_PATTERNS/RD_XFER_TYPE[1]_net_1\, Y => 
        HIEFFPLA_NET_0_119338);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_0[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116822, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_3, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_0[2]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_5[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116660, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_11, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_5[1]\);
    
    \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_2S_2_0\ : DFN1C0
      port map(D => 
        \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_1S_0_net_1\, CLK
         => CLK60MHZ, CLR => P_MASTER_POR_B_c_0_0, Q => 
        P_USB_MASTER_EN_c_2_0);
    
    HIEFFPLA_INST_0_52363 : AND2A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[8]_net_1\, B => 
        HIEFFPLA_NET_0_117570, Y => HIEFFPLA_NET_0_117574);
    
    HIEFFPLA_INST_0_39952 : MX2
      port map(A => HIEFFPLA_NET_0_119911, B => 
        \U50_PATTERNS/ELINK_BLKA[11]\, S => 
        \U50_PATTERNS/SM_BANK_SEL[20]\, Y => 
        HIEFFPLA_NET_0_119933);
    
    HIEFFPLA_INST_0_58523 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_16[2]\, B => 
        HIEFFPLA_NET_0_116506, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_1[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116510);
    
    HIEFFPLA_INST_0_52164 : OA1A
      port map(A => HIEFFPLA_NET_0_117689, B => 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM[6]_net_1\, C => 
        HIEFFPLA_NET_0_117616, Y => HIEFFPLA_NET_0_117618);
    
    \U_ELK16_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]\ : DFN1C0
      port map(D => \U_ELK16_CH/U_SLAVE_1ELK/Q[3]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[3]_net_1\);
    
    \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[5]\ : DFN1C0
      port map(D => 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\);
    
    HIEFFPLA_INST_0_60636 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_13[0]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_14[0]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_3[0]\, Y => 
        HIEFFPLA_NET_0_116240);
    
    HIEFFPLA_INST_0_37107 : AND3B
      port map(A => \U200A_TFC/LOC_STRT_ADDR[2]\, B => 
        HIEFFPLA_NET_0_120293, C => HIEFFPLA_NET_0_120328, Y => 
        HIEFFPLA_NET_0_120346);
    
    \U_ELK12_CH/U_SLAVE_1ELK/RECD_SER_WORD[0]\ : DFN1C0
      port map(D => \U_ELK12_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[0]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_12[0]\);
    
    HIEFFPLA_INST_0_54770 : AND3B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[3]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[0]_net_1\, C => 
        HIEFFPLA_NET_0_117236, Y => HIEFFPLA_NET_0_117204);
    
    HIEFFPLA_INST_0_39821 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_8[3]\, B => 
        HIEFFPLA_NET_0_119520, S => HIEFFPLA_NET_0_119291, Y => 
        HIEFFPLA_NET_0_119948);
    
    HIEFFPLA_INST_0_37621 : XO1
      port map(A => HIEFFPLA_NET_0_120150, B => \ELKS_ADDRB[1]\, 
        C => \U200B_ELINKS/GP_PG_SM[10]_net_1\, Y => 
        HIEFFPLA_NET_0_120245);
    
    \U_ELK8_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]\ : DFN1C0
      port map(D => \U_ELK8_CH/U_SLAVE_1ELK/Q[9]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_14[4]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116231, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_2, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_14[4]\);
    
    \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[6]\ : DFN1C0
      port map(D => 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[6]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\);
    
    \U_ELK7_CH/U_SLAVE_1ELK/RECD_SER_WORD[7]\ : DFN1C0
      port map(D => \U_ELK7_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[7]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_7[7]\);
    
    \U_ELK12_CH/U_SLAVE_1ELK/RECD_SER_WORD[1]\ : DFN1C0
      port map(D => \U_ELK12_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[1]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_12[1]\);
    
    HIEFFPLA_INST_0_59979 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_4[3]\, B => 
        HIEFFPLA_NET_0_116323, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_2[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116326);
    
    HIEFFPLA_INST_0_54618 : MX2
      port map(A => HIEFFPLA_NET_0_117306, B => 
        HIEFFPLA_NET_0_117296, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[2]_net_1\, Y => 
        HIEFFPLA_NET_0_117232);
    
    HIEFFPLA_INST_0_54373 : MX2
      port map(A => HIEFFPLA_NET_0_116140, B => 
        HIEFFPLA_NET_0_116239, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_2[3]_net_1\, Y
         => HIEFFPLA_NET_0_117274);
    
    \U50_PATTERNS/U4C_REGCROSS/SAMP_ONE[7]\ : DFN1C0
      port map(D => \U50_PATTERNS/ELINKS_STRT_ADDR[7]\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_33, Q => 
        \U50_PATTERNS/U4C_REGCROSS/SAMP_ONE[7]_net_1\);
    
    \U_ELK7_CH/U_SLAVE_1ELK/Q[9]\ : DFN1C0
      port map(D => \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/Q[9]_net_1\);
    
    HIEFFPLA_INST_0_45174 : NAND3C
      port map(A => HIEFFPLA_NET_0_118878, B => 
        HIEFFPLA_NET_0_118730, C => HIEFFPLA_NET_0_118800, Y => 
        HIEFFPLA_NET_0_118972);
    
    HIEFFPLA_INST_0_50399 : MX2
      port map(A => HIEFFPLA_NET_0_117954, B => 
        HIEFFPLA_NET_0_117952, S => \BIT_OS_SEL_5[1]\, Y => 
        HIEFFPLA_NET_0_117956);
    
    HIEFFPLA_INST_0_51716 : NAND2B
      port map(A => 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM[4]_net_1\, B => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[42]_net_1\, Y => 
        HIEFFPLA_NET_0_117710);
    
    \U_ELK16_CH/U_SLAVE_1ELK/Q[0]\ : DFN1C0
      port map(D => \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/Q[0]_net_1\);
    
    HIEFFPLA_INST_0_45127 : MX2
      port map(A => HIEFFPLA_NET_0_118970, B => 
        \U50_PATTERNS/WR_USB_ADBUS[5]\, S => 
        HIEFFPLA_NET_0_119486, Y => HIEFFPLA_NET_0_118980);
    
    HIEFFPLA_INST_0_39272 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_19[6]\, B => 
        HIEFFPLA_NET_0_119517, S => HIEFFPLA_NET_0_119293, Y => 
        HIEFFPLA_NET_0_120009);
    
    \U_ELK14_CH/U_ELK1_SERDAT_SOURCE/SERDAT[7]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118456, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_6, Q => 
        \U_ELK14_CH/ELK_TX_DAT[7]\);
    
    HIEFFPLA_INST_0_45249 : AO1
      port map(A => HIEFFPLA_NET_0_119290, B => 
        \U50_PATTERNS/ELINK_DOUTA_17[0]\, C => 
        HIEFFPLA_NET_0_118837, Y => HIEFFPLA_NET_0_118958);
    
    HIEFFPLA_INST_0_45791 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/SM_BANK_SEL[16]\, C => 
        \U50_PATTERNS/ELINK_DOUTA_3[4]\, Y => 
        HIEFFPLA_NET_0_118841);
    
    \U_ELK6_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]\ : DFN1C0
      port map(D => \U_ELK6_CH/U_SLAVE_1ELK/Q[9]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]_net_1\);
    
    HIEFFPLA_INST_0_45701 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_19[5]\, C => 
        \U50_PATTERNS/SM_BANK_SEL[0]\, Y => HIEFFPLA_NET_0_118862);
    
    HIEFFPLA_INST_0_44830 : NOR3A
      port map(A => HIEFFPLA_NET_0_119370, B => 
        \U50_PATTERNS/REG_STATE[4]_net_1\, C => 
        \U50_PATTERNS/REG_STATE[3]_net_1\, Y => 
        HIEFFPLA_NET_0_119039);
    
    HIEFFPLA_INST_0_37821 : AND3B
      port map(A => HIEFFPLA_NET_0_120188, B => 
        \U200B_ELINKS/GP_PG_SM[9]_net_1\, C => \OP_MODE_c[6]\, Y
         => HIEFFPLA_NET_0_120198);
    
    \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_2S_18\ : DFN1C0
      port map(D => 
        \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_1S_0_net_1\, CLK
         => CLK60MHZ, CLR => \U_EXEC_MASTER/P_MASTER_POR_B_c_0\, 
        Q => P_USB_MASTER_EN_c_18);
    
    \U_EXEC_MASTER/MPOR_B_25\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117787, CLK => CLK_40M_GL, CLR
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_0\, Q => 
        P_MASTER_POR_B_c_25);
    
    HIEFFPLA_INST_0_56395 : NAND3C
      port map(A => HIEFFPLA_NET_0_116830, B => 
        HIEFFPLA_NET_0_116846, C => HIEFFPLA_NET_0_116854, Y => 
        HIEFFPLA_NET_0_116878);
    
    \U50_PATTERNS/ELINK_DINA_6[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119741, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_16, Q => 
        \U50_PATTERNS/ELINK_DINA_6[2]\);
    
    HIEFFPLA_INST_0_53233 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_CLKPHASE[3]\, B => 
        HIEFFPLA_NET_0_117444, S => HIEFFPLA_NET_0_117111, Y => 
        HIEFFPLA_NET_0_117449);
    
    HIEFFPLA_INST_0_45298 : AO1
      port map(A => HIEFFPLA_NET_0_119277, B => 
        \U50_PATTERNS/ELINK_DOUTA_11[1]\, C => 
        HIEFFPLA_NET_0_118827, Y => HIEFFPLA_NET_0_118948);
    
    HIEFFPLA_INST_0_45051 : NAND3C
      port map(A => HIEFFPLA_NET_0_119432, B => 
        \U50_PATTERNS/USB_TXE_B\, C => HIEFFPLA_NET_0_119379, Y
         => HIEFFPLA_NET_0_118991);
    
    HIEFFPLA_INST_0_50419 : MX2
      port map(A => \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\, B
         => \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\, S => 
        \BIT_OS_SEL_5[2]\, Y => HIEFFPLA_NET_0_117953);
    
    HIEFFPLA_INST_0_37441 : MX2
      port map(A => \U200A_TFC/LOC_STOP_ADDR[6]\, B => 
        \TFC_STOP_ADDR[6]\, S => \U200A_TFC/GP_PG_SM_0[10]_net_1\, 
        Y => HIEFFPLA_NET_0_120284);
    
    \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[8]\ : DFN1C0
      port map(D => 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\);
    
    \U50_PATTERNS/ELINK_ADDRA_1[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120006, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_20, Q => 
        \U50_PATTERNS/ELINK_ADDRA_1[1]\);
    
    \U_ELK10_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]\ : DFN1C0
      port map(D => \U_ELK10_CH/U_SLAVE_1ELK/Q[9]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]_net_1\);
    
    \U_ELK0_SERDAT_SOURCE/SERDAT[7]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118653, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_10, Q => \ELK0_TX_DAT[7]\);
    
    HIEFFPLA_INST_0_56340 : AO1
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[7]_net_1\, B => 
        HIEFFPLA_NET_0_117429, C => HIEFFPLA_NET_0_116866, Y => 
        HIEFFPLA_NET_0_116890);
    
    \U_ELK18_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]\ : DFN1C0
      port map(D => \U_ELK18_CH/U_SLAVE_1ELK/Q[5]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]_net_1\);
    
    HIEFFPLA_INST_0_56988 : XA1C
      port map(A => HIEFFPLA_NET_0_116778, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_1[8]\, C => 
        HIEFFPLA_NET_0_117179, Y => HIEFFPLA_NET_0_116759);
    
    \U_ELK19_CH/U_ELK1_SERDAT_SOURCE/SERDAT[7]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118231, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_15, Q => 
        \U_ELK19_CH/ELK_TX_DAT[7]\);
    
    HIEFFPLA_INST_0_43197 : AND3A
      port map(A => \U50_PATTERNS/REG_STATE_0[2]_net_1\, B => 
        HIEFFPLA_NET_0_119377, C => 
        \U50_PATTERNS/REG_STATE_0[4]_net_1\, Y => 
        HIEFFPLA_NET_0_119349);
    
    \U200A_TFC/GP_PG_SM[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120318, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_28, Q => 
        \U200A_TFC/GP_PG_SM[3]_net_1\);
    
    HIEFFPLA_INST_0_57860 : AOI1A
      port map(A => HIEFFPLA_NET_0_116622, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_6[5]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_6[6]\, Y => 
        HIEFFPLA_NET_0_116605);
    
    \U_ELK3_CH/U_ELK1_CMD_TX/START_RISE\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118104, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_3, Q => 
        \U_ELK3_CH/U_ELK1_CMD_TX/START_RISE_net_1\);
    
    \U_ELK4_CH/U_ELK1_SERDAT_SOURCE/SERDAT[7]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118051, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_16, Q => 
        \U_ELK4_CH/ELK_TX_DAT[7]\);
    
    \U_ELK10_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0\ : DFN1C0
      port map(D => CLK_40M_GL, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_5, Q => 
        \U_ELK10_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0_net_1\);
    
    HIEFFPLA_INST_0_56970 : AND3B
      port map(A => HIEFFPLA_NET_0_117085, B => 
        HIEFFPLA_NET_0_116757, C => HIEFFPLA_NET_0_116777, Y => 
        HIEFFPLA_NET_0_116762);
    
    \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[14]\ : DFN1C0
      port map(D => 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[14]_net_1\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[14]_net_1\);
    
    \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM[5]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117618, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_22_0, Q => 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM[5]_net_1\);
    
    \U_ELK9_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL\ : DFN1C0
      port map(D => \U_ELK9_CH/ELK_IN_F_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL_net_1\);
    
    \U_ELK19_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118241, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_4, Q => 
        \U_ELK19_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]_net_1\);
    
    HIEFFPLA_INST_0_56804 : XA1C
      port map(A => HIEFFPLA_NET_0_116807, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_0[7]\, C => 
        HIEFFPLA_NET_0_117179, Y => HIEFFPLA_NET_0_116793);
    
    HIEFFPLA_INST_0_39812 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_8[2]\, B => 
        HIEFFPLA_NET_0_119522, S => HIEFFPLA_NET_0_119291, Y => 
        HIEFFPLA_NET_0_119949);
    
    \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117620, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_22, Q => 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM[1]_net_1\);
    
    \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[14]\ : DFN1C0
      port map(D => \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\, 
        CLK => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[14]_net_1\);
    
    HIEFFPLA_INST_0_57481 : AND2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_4[3]\, B => 
        HIEFFPLA_NET_0_116683, Y => HIEFFPLA_NET_0_116673);
    
    HIEFFPLA_INST_0_52660 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_17[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_18[1]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_3[0]\, Y => 
        HIEFFPLA_NET_0_117531);
    
    \U_ELK1_CH/U_ELK1_SERDAT_SOURCE/SERDAT[4]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118189, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_11, Q => 
        \U_ELK1_CH/ELK_TX_DAT[4]\);
    
    HIEFFPLA_INST_0_50827 : MX2
      port map(A => 
        \U_ELK8_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]_net_1\, B => 
        \U_ELK8_CH/ELK_TX_DAT[4]\, S => 
        \U_ELK8_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_117885);
    
    \U50_PATTERNS/ELINKS_STOP_ADDR[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120121, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_14, Q => 
        \U50_PATTERNS/ELINKS_STOP_ADDR[6]\);
    
    HIEFFPLA_INST_0_52125 : NAND3C
      port map(A => HIEFFPLA_NET_0_117627, B => 
        HIEFFPLA_NET_0_117629, C => 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM_0[4]_net_1\, Y => 
        HIEFFPLA_NET_0_117631);
    
    HIEFFPLA_INST_0_44464 : MX2
      port map(A => \ELKS_STRT_ADDR[2]\, B => 
        \U50_PATTERNS/U4C_REGCROSS/SAMP_TWO[2]_net_1\, S => 
        HIEFFPLA_NET_0_119114, Y => HIEFFPLA_NET_0_119110);
    
    HIEFFPLA_INST_0_38258 : MX2
      port map(A => \U50_PATTERNS/ELINKS_STOP_ADDR[2]\, B => 
        \U50_PATTERNS/ELINKS_STOP_ADDR_T[2]\, S => 
        HIEFFPLA_NET_0_119472, Y => HIEFFPLA_NET_0_120125);
    
    \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_2S_14\ : DFN1C0
      port map(D => 
        \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_1S_0_net_1\, CLK
         => CLK60MHZ, CLR => \U_EXEC_MASTER/P_MASTER_POR_B_c_0\, 
        Q => P_USB_MASTER_EN_c_14);
    
    HIEFFPLA_INST_0_54540 : MX2
      port map(A => HIEFFPLA_NET_0_117250, B => 
        HIEFFPLA_NET_0_117323, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[1]_net_1\, Y => 
        HIEFFPLA_NET_0_117253);
    
    HIEFFPLA_INST_0_51741 : MX2
      port map(A => \U_MASTER_DES/U13A_ADJ_160M/BITCNT[1]\, B => 
        HIEFFPLA_NET_0_117680, S => HIEFFPLA_NET_0_117630, Y => 
        HIEFFPLA_NET_0_117697);
    
    HIEFFPLA_INST_0_49049 : MX2
      port map(A => HIEFFPLA_NET_0_118204, B => 
        HIEFFPLA_NET_0_118219, S => \BIT_OS_SEL_0[1]\, Y => 
        HIEFFPLA_NET_0_118206);
    
    \U50_PATTERNS/ELINK_ADDRA_17[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120030, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_10, Q => 
        \U50_PATTERNS/ELINK_ADDRA_17[1]\);
    
    HIEFFPLA_INST_0_60893 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_17[3]\, B => 
        HIEFFPLA_NET_0_117186, S => HIEFFPLA_NET_0_117169, Y => 
        HIEFFPLA_NET_0_116202);
    
    \U50_PATTERNS/U4A_REGCROSS/SAMP_ONE[5]\ : DFN1C0
      port map(D => \U50_PATTERNS/TFC_STRT_ADDR[5]\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_32_0, Q => 
        \U50_PATTERNS/U4A_REGCROSS/SAMP_ONE[5]_net_1\);
    
    HIEFFPLA_INST_0_38957 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_15[3]\, B => 
        HIEFFPLA_NET_0_119520, S => HIEFFPLA_NET_0_119297, Y => 
        HIEFFPLA_NET_0_120044);
    
    \U_MASTER_DES/U13C_MASTER_DESER/ARB_WRD_40M_FIXED[5]\ : 
        DFN1C0
      port map(D => \U_MASTER_DES/U13C_MASTER_DESER/Q[5]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_26, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_WRD_40M_FIXED[5]_net_1\);
    
    \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[14]\ : DFN1C0
      port map(D => \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/ADJ_Q[14]_net_1\);
    
    \U_ELK19_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]\ : DFN1C0
      port map(D => \U_ELK19_CH/U_SLAVE_1ELK/Q[7]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]_net_1\);
    
    HIEFFPLA_INST_0_50254 : MX2
      port map(A => HIEFFPLA_NET_0_118002, B => 
        HIEFFPLA_NET_0_117997, S => \BIT_OS_SEL_0[0]\, Y => 
        \U_ELK5_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[3]\);
    
    HIEFFPLA_INST_0_47796 : MX2
      port map(A => HIEFFPLA_NET_0_118442, B => 
        HIEFFPLA_NET_0_118430, S => \BIT_OS_SEL_4[0]\, Y => 
        \U_ELK14_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[7]\);
    
    HIEFFPLA_INST_0_63056 : AND2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[12]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[8]\, Y => 
        HIEFFPLA_NET_0_115900);
    
    \U_MAINCLKGEN/Core\ : DYNCCC
      generic map(VCOFREQUENCY => 160.0)

      port map(CLKA => CLK_40M_BUF_RECD, EXTFB => \GND\, 
        POWERDOWN => \VCC\, GLA => CLK_40M_GL, LOCK => 
        CCC_MAIN_LOCK, CLKB => \GND\, GLB => CCC_160M_FXD, YB => 
        OPEN, CLKC => USBCLK60MHZ_c, GLC => CLK60MHZ, YC => OPEN, 
        SDIN => \GND\, SCLK => \GND\, SSHIFT => \GND\, SUPDATE
         => \GND\, MODE => \GND\, SDOUT => OPEN, OADIV0 => \VCC\, 
        OADIV1 => \VCC\, OADIV2 => \GND\, OADIV3 => \GND\, OADIV4
         => \GND\, OAMUX0 => \GND\, OAMUX1 => \GND\, OAMUX2 => 
        \VCC\, DLYGLA0 => \GND\, DLYGLA1 => \GND\, DLYGLA2 => 
        \GND\, DLYGLA3 => \GND\, DLYGLA4 => \GND\, OBDIV0 => 
        \GND\, OBDIV1 => \GND\, OBDIV2 => \GND\, OBDIV3 => \GND\, 
        OBDIV4 => \GND\, OBMUX0 => \GND\, OBMUX1 => \GND\, OBMUX2
         => \VCC\, DLYYB0 => \GND\, DLYYB1 => \GND\, DLYYB2 => 
        \GND\, DLYYB3 => \GND\, DLYYB4 => \GND\, DLYGLB0 => \GND\, 
        DLYGLB1 => \GND\, DLYGLB2 => \VCC\, DLYGLB3 => \VCC\, 
        DLYGLB4 => \GND\, OCDIV0 => \GND\, OCDIV1 => \GND\, 
        OCDIV2 => \GND\, OCDIV3 => \GND\, OCDIV4 => \GND\, OCMUX0
         => \GND\, OCMUX1 => \GND\, OCMUX2 => \GND\, DLYYC0 => 
        \GND\, DLYYC1 => \GND\, DLYYC2 => \GND\, DLYYC3 => \GND\, 
        DLYYC4 => \GND\, DLYGLC0 => \VCC\, DLYGLC1 => \GND\, 
        DLYGLC2 => \VCC\, DLYGLC3 => \VCC\, DLYGLC4 => \VCC\, 
        FINDIV0 => \VCC\, FINDIV1 => \VCC\, FINDIV2 => \VCC\, 
        FINDIV3 => \GND\, FINDIV4 => \GND\, FINDIV5 => \GND\, 
        FINDIV6 => \GND\, FBDIV0 => \VCC\, FBDIV1 => \VCC\, 
        FBDIV2 => \VCC\, FBDIV3 => \VCC\, FBDIV4 => \VCC\, FBDIV5
         => \GND\, FBDIV6 => \GND\, FBDLY0 => \GND\, FBDLY1 => 
        \GND\, FBDLY2 => \VCC\, FBDLY3 => \GND\, FBDLY4 => \GND\, 
        FBSEL0 => \GND\, FBSEL1 => \VCC\, XDLYSEL => \GND\, 
        VCOSEL0 => \GND\, VCOSEL1 => \GND\, VCOSEL2 => \VCC\);
    
    HIEFFPLA_INST_0_46355 : AO1A
      port map(A => HIEFFPLA_NET_0_118857, B => 
        \U50_PATTERNS/SM_BANK_SEL[1]\, C => HIEFFPLA_NET_0_118849, 
        Y => HIEFFPLA_NET_0_118709);
    
    HIEFFPLA_INST_0_44656 : MX2
      port map(A => \OP_MODE[0]\, B => 
        \U50_PATTERNS/U4E_REGCROSS/SAMP_TWO[0]_net_1\, S => 
        HIEFFPLA_NET_0_119072, Y => HIEFFPLA_NET_0_119070);
    
    \U50_PATTERNS/ELINK_DINA_16[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119810, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_18, Q => 
        \U50_PATTERNS/ELINK_DINA_16[5]\);
    
    HIEFFPLA_INST_0_57970 : NAND3C
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_7[7]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_7[8]\, C => 
        HIEFFPLA_NET_0_116587, Y => HIEFFPLA_NET_0_116588);
    
    \U_ELK7_CH/U_SLAVE_1ELK/RECD_SER_WORD[5]\ : DFN1C0
      port map(D => \U_ELK7_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[5]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_7[5]\);
    
    \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[76]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117705, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_33, Q => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[76]_net_1\);
    
    HIEFFPLA_INST_0_54946 : AND2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_3[6]_net_1\, B => 
        HIEFFPLA_NET_0_117217, Y => HIEFFPLA_NET_0_117162);
    
    HIEFFPLA_INST_0_52117 : MX2
      port map(A => HIEFFPLA_NET_0_117663, B => 
        HIEFFPLA_NET_0_117662, S => 
        \U_MASTER_DES/U13A_ADJ_160M/BITCNT[5]\, Y => 
        HIEFFPLA_NET_0_117633);
    
    \U0B_TX40M_REFCLK/\\\\OUTBUF_LVDS[0]\\\\/U0/U2\ : IOPADN_OUT
      port map(DB => 
        \U0B_TX40M_REFCLK/\\\\OUTBUF_LVDS[0]\\\\/U0/NET1\, PAD
         => TX_CLK40M_N);
    
    \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_2[4]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_115935, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_24_0, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_2[4]_net_1\);
    
    HIEFFPLA_INST_0_56297 : NAND3C
      port map(A => HIEFFPLA_NET_0_116874, B => 
        HIEFFPLA_NET_0_116882, C => HIEFFPLA_NET_0_116890, Y => 
        HIEFFPLA_NET_0_116898);
    
    HIEFFPLA_INST_0_37187 : AND3B
      port map(A => \U200A_TFC/GP_PG_SM[4]_net_1\, B => 
        \U200A_TFC/GP_PG_SM[5]_net_1\, C => HIEFFPLA_NET_0_120326, 
        Y => HIEFFPLA_NET_0_120330);
    
    \U50_PATTERNS/ELINK_RWA[15]/U1\ : DFN1P0
      port map(D => HIEFFPLA_NET_0_119705, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_12, Q => 
        \U50_PATTERNS/ELINK_RWA[15]\);
    
    HIEFFPLA_INST_0_61802 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_26[4]\, B => 
        HIEFFPLA_NET_0_117100, S => HIEFFPLA_NET_0_117138, Y => 
        HIEFFPLA_NET_0_116076);
    
    HIEFFPLA_INST_0_59694 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_2[0]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_18[0]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_1[4]_net_1\, Y
         => HIEFFPLA_NET_0_116360);
    
    HIEFFPLA_INST_0_43252 : AO1
      port map(A => \U50_PATTERNS/REG_STATE[5]_net_1\, B => 
        \U50_PATTERNS/REG_STATE[1]_net_1\, C => 
        HIEFFPLA_NET_0_119015, Y => HIEFFPLA_NET_0_119337);
    
    HIEFFPLA_INST_0_50447 : MX2
      port map(A => \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\, B
         => \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\, S => 
        \BIT_OS_SEL_5[2]\, Y => HIEFFPLA_NET_0_117949);
    
    HIEFFPLA_INST_0_55842 : MX2
      port map(A => HIEFFPLA_NET_0_116966, B => 
        HIEFFPLA_NET_0_117000, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[2]\, Y => 
        HIEFFPLA_NET_0_116983);
    
    \DCB_SALT_SEL_pad/U0/U0\ : IOPAD_IN_U
      port map(PAD => DCB_SALT_SEL, Y => 
        \DCB_SALT_SEL_pad/U0/NET1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_9[4]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_115961, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_20, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_9[4]\);
    
    HIEFFPLA_INST_0_56335 : AO1
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[6]_net_1\, B => 
        HIEFFPLA_NET_0_117429, C => HIEFFPLA_NET_0_116867, Y => 
        HIEFFPLA_NET_0_116891);
    
    HIEFFPLA_INST_0_55064 : AND2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[6]_net_1\, B => 
        HIEFFPLA_NET_0_117393, Y => HIEFFPLA_NET_0_117130);
    
    \U_ELK4_CH/U_SLAVE_1ELK/Q[5]\ : DFN1C0
      port map(D => \U_ELK4_CH/U_SLAVE_1ELK/ADJ_Q[5]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK4_CH/U_SLAVE_1ELK/Q[5]_net_1\);
    
    \U50_PATTERNS/ELK_N_ACTIVE\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119628, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_22, Q => 
        \U50_PATTERNS/ELK_N_ACTIVE_net_1\);
    
    HIEFFPLA_INST_0_54269 : MX2
      port map(A => HIEFFPLA_NET_0_116208, B => 
        HIEFFPLA_NET_0_116098, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_2[3]_net_1\, Y
         => HIEFFPLA_NET_0_117287);
    
    \U50_PATTERNS/U4C_REGCROSS/SAMP_ONE[5]\ : DFN1C0
      port map(D => \U50_PATTERNS/ELINKS_STRT_ADDR[5]\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_33, Q => 
        \U50_PATTERNS/U4C_REGCROSS/SAMP_ONE[5]_net_1\);
    
    HIEFFPLA_INST_0_61241 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_4[3]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_20[3]\, S
         => \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_5[4]_net_1\, 
        Y => HIEFFPLA_NET_0_116155);
    
    HIEFFPLA_INST_0_50037 : MX2
      port map(A => HIEFFPLA_NET_0_118050, B => 
        HIEFFPLA_NET_0_118025, S => \BIT_OS_SEL_1[0]\, Y => 
        \U_ELK4_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[7]\);
    
    \U_ELK17_CH/ELK_IN_R\ : DFN1C0
      port map(D => \U_ELK17_CH/ELK_IN_DDR_R\, CLK => 
        CCC_160M_ADJ, CLR => DEV_RST_B_c, Q => 
        \U_ELK17_CH/ELK_IN_R_net_1\);
    
    HIEFFPLA_INST_0_51451 : OA1A
      port map(A => HIEFFPLA_NET_0_117779, B => 
        \U_EXEC_MASTER/DEL_CNT[7]\, C => 
        \U_EXEC_MASTER/CCC_1_LOCK_STAT_1D_net_1\, Y => 
        HIEFFPLA_NET_0_117770);
    
    \U_ELK17_CH/U_SLAVE_1ELK/Q[3]\ : DFN1C0
      port map(D => \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/Q[3]_net_1\);
    
    \U200B_ELINKS/GP_PG_SM[6]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120209, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_29, Q => 
        \U200B_ELINKS/GP_PG_SM[6]_net_1\);
    
    AFLSDF_INV_7 : INV
      port map(A => P_USB_MASTER_EN_c_22, Y => \AFLSDF_INV_7\);
    
    \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[12]\ : DFN1C0
      port map(D => \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\, 
        CLK => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\);
    
    \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[6]\ : DFN1C0
      port map(D => \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\);
    
    HIEFFPLA_INST_0_53919 : MX2
      port map(A => HIEFFPLA_NET_0_117399, B => 
        HIEFFPLA_NET_0_117315, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[1]_net_1\, Y
         => HIEFFPLA_NET_0_117333);
    
    HIEFFPLA_INST_0_42706 : AND3
      port map(A => HIEFFPLA_NET_0_119511, B => 
        \U50_PATTERNS/REG_STATE_0[4]_net_1\, C => 
        HIEFFPLA_NET_0_119448, Y => HIEFFPLA_NET_0_119478);
    
    HIEFFPLA_INST_0_43121 : AO1A
      port map(A => \U50_PATTERNS/REG_STATE[0]_net_1\, B => 
        \U50_PATTERNS/REG_STATE[1]_net_1\, C => 
        \U50_PATTERNS/REG_STATE[3]_net_1\, Y => 
        HIEFFPLA_NET_0_119368);
    
    HIEFFPLA_INST_0_42265 : NAND2B
      port map(A => \U50_PATTERNS/RD_USB_ADBUS[6]\, B => 
        HIEFFPLA_NET_0_119020, Y => HIEFFPLA_NET_0_119585);
    
    \U50_PATTERNS/ELINK_DINA_3[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119763, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_11, Q => 
        \U50_PATTERNS/ELINK_DINA_3[4]\);
    
    HIEFFPLA_INST_0_56549 : AND3A
      port map(A => HIEFFPLA_NET_0_117430, B => \BIT_OS_SEL_1[2]\, 
        C => \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[13]_net_1\, 
        Y => HIEFFPLA_NET_0_116841);
    
    HIEFFPLA_INST_0_48869 : AND2A
      port map(A => \OP_MODE_c_6[1]\, B => \PATT_ELK_DAT_19[5]\, 
        Y => HIEFFPLA_NET_0_118233);
    
    \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[8]\ : DFN1C0
      port map(D => \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\);
    
    \U200B_ELINKS/LOC_STRT_ADDR[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120175, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_11, Q => 
        \U200B_ELINKS/LOC_STRT_ADDR[4]\);
    
    HIEFFPLA_INST_0_45931 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_7[4]\, C => 
        \U50_PATTERNS/SM_BANK_SEL[12]\, Y => 
        HIEFFPLA_NET_0_118808);
    
    \U_ELK2_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]\ : DFN1C0
      port map(D => \U_ELK2_CH/U_SLAVE_1ELK/Q[2]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]_net_1\);
    
    \U_ELK8_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U1\ : IOBI_ID_OD_EB
      port map(DR => \U_ELK8_CH/ELK_OUT_R\, DF => 
        \U_ELK8_CH/ELK_OUT_F\, CLR => \GND\, E => \AFLSDF_INV_48\, 
        ICLK => CCC_160M_ADJ, OCLK => CCC_160M_FXD, YIN => 
        \U_ELK8_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\, DOUT => 
        \U_ELK8_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, EOUT => 
        \U_ELK8_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET2\, YR => 
        \U_ELK8_CH/ELK_IN_DDR_R\, YF => \U_ELK8_CH/ELK_IN_DDR_F\);
    
    HIEFFPLA_INST_0_46979 : MX2
      port map(A => HIEFFPLA_NET_0_118589, B => 
        HIEFFPLA_NET_0_118585, S => \BIT_OS_SEL_4[1]\, Y => 
        HIEFFPLA_NET_0_118576);
    
    \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[1]\\\\/U0/U0\ : 
        IOPAD_BI_U
      port map(D => 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[1]\\\\/U0/NET1\, 
        E => 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[1]\\\\/U0/NET2\, 
        Y => 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[1]\\\\/U0/NET3\, 
        PAD => BIDIR_USB_ADBUS(1));
    
    HIEFFPLA_INST_0_53502 : MX2
      port map(A => HIEFFPLA_NET_0_117275, B => 
        HIEFFPLA_NET_0_117260, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[2]_net_1\, Y
         => HIEFFPLA_NET_0_117399);
    
    \U_ELK11_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118601, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_7, Q => 
        \U_ELK11_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]_net_1\);
    
    \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[2]\ : DFN1C0
      port map(D => \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK15_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\);
    
    \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[49]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117723, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_19, Q => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[49]\);
    
    \U_ELK18_CH/U_SLAVE_1ELK/RECD_SER_WORD[6]\ : DFN1C0
      port map(D => \U_ELK18_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[6]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_18[6]\);
    
    \U_ELK14_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118472, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_5, Q => 
        \U_ELK14_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]_net_1\);
    
    \U50_PATTERNS/ELINK_ADDRA_3[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119987, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_1, Q => 
        \U50_PATTERNS/ELINK_ADDRA_3[4]\);
    
    HIEFFPLA_INST_0_61556 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_23[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_24[1]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[0]\, Y => 
        HIEFFPLA_NET_0_116110);
    
    HIEFFPLA_INST_0_38975 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_15[5]\, B => 
        HIEFFPLA_NET_0_119518, S => HIEFFPLA_NET_0_119297, Y => 
        HIEFFPLA_NET_0_120042);
    
    AFLSDF_INV_41 : INV
      port map(A => DCB_SALT_SEL_c, Y => \AFLSDF_INV_41\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_7[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_115979, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_17_0, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_7[1]\);
    
    \U_ELK18_CH/U_ELK1_CMD_TX/SER_OUT_FI\ : DFN1C0
      port map(D => 
        \U_ELK18_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_9, Q => 
        \U_ELK18_CH/U_ELK1_CMD_TX/SER_OUT_FI_net_1\);
    
    HIEFFPLA_INST_0_37934 : MX2
      port map(A => \U200B_ELINKS/LOC_STOP_ADDR[0]\, B => 
        \ELKS_STOP_ADDR[0]\, S => 
        \U200B_ELINKS/GP_PG_SM_0[10]_net_1\, Y => 
        HIEFFPLA_NET_0_120187);
    
    \U_ELK3_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118110, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_16, Q => 
        \U_ELK3_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_23[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116439, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_17_0, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_23[3]\);
    
    \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[1]\ : DFN1C0
      port map(D => 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/ARB_BYTE[1]_net_1\);
    
    \U_ELK6_CH/U_SLAVE_1ELK/Q[6]\ : DFN1C0
      port map(D => \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/Q[6]_net_1\);
    
    HIEFFPLA_INST_0_53255 : AND2A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[8]_net_1\, B => 
        HIEFFPLA_NET_0_115873, Y => HIEFFPLA_NET_0_117443);
    
    HIEFFPLA_INST_0_37268 : AND3
      port map(A => HIEFFPLA_NET_0_120327, B => 
        HIEFFPLA_NET_0_120333, C => HIEFFPLA_NET_0_120302, Y => 
        HIEFFPLA_NET_0_120310);
    
    \U_ELK2_CH/U_ELK1_CMD_TX/SER_OUT_FDEL\ : DFN1C0
      port map(D => \U_ELK2_CH/U_ELK1_CMD_TX/SER_OUT_FI_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_12, Q
         => \U_ELK2_CH/ELK_OUT_F\);
    
    \U_ELK11_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118603, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_7, Q => 
        \U_ELK11_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[0]_net_1\);
    
    \U50_PATTERNS/ELINKS_STOP_ADDR_T[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120112, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_7, Q => 
        \U50_PATTERNS/ELINKS_STOP_ADDR_T[7]\);
    
    HIEFFPLA_INST_0_44280 : MX2
      port map(A => \TFC_STRT_ADDR[5]\, B => 
        \U50_PATTERNS/U4A_REGCROSS/SAMP_TWO[5]_net_1\, S => 
        HIEFFPLA_NET_0_119156, Y => HIEFFPLA_NET_0_119149);
    
    HIEFFPLA_INST_0_42173 : MX2
      port map(A => \U50_PATTERNS/OP_MODE_T[2]\, B => 
        \U50_PATTERNS/RD_USB_ADBUS[2]\, S => 
        HIEFFPLA_NET_0_119440, Y => HIEFFPLA_NET_0_119607);
    
    \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[9]\ : DFN1C0
      port map(D => 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[9]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\);
    
    HIEFFPLA_INST_0_54952 : AND2A
      port map(A => HIEFFPLA_NET_0_117219, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_3[6]_net_1\, Y => 
        HIEFFPLA_NET_0_117159);
    
    HIEFFPLA_INST_0_60019 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_5[1]\, B => 
        HIEFFPLA_NET_0_116677, S => HIEFFPLA_NET_0_117156, Y => 
        HIEFFPLA_NET_0_116321);
    
    HIEFFPLA_INST_0_47618 : AND2
      port map(A => CLK_40M_GL, B => 
        \U_ELK14_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0_net_1\, Y => 
        HIEFFPLA_NET_0_118464);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_1[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116473, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_17_0, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_1[2]\);
    
    \U_ELK0_CMD_TX/SER_OUT_RDEL\ : DFN1P0
      port map(D => \U_ELK0_CMD_TX/SER_OUT_RI_i\, CLK => 
        CCC_160M_FXD, PRE => MASTER_SALT_POR_B_i_0_i_7, Q => 
        ELK0_OUT_R_i_0);
    
    \U50_PATTERNS/OP_MODE_T[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119608, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_17, Q => 
        \U50_PATTERNS/OP_MODE_T[1]\);
    
    HIEFFPLA_INST_0_48318 : MX2
      port map(A => \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[0]_net_1\, 
        B => \U_ELK16_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\, S => 
        \BIT_OS_SEL_1[2]\, Y => HIEFFPLA_NET_0_118339);
    
    HIEFFPLA_INST_0_54434 : MX2
      port map(A => HIEFFPLA_NET_0_117331, B => 
        HIEFFPLA_NET_0_117303, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[2]_net_1\, Y => 
        HIEFFPLA_NET_0_117266);
    
    HIEFFPLA_INST_0_51725 : NAND2B
      port map(A => 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM[4]_net_1\, B => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[7]_net_1\, Y => 
        HIEFFPLA_NET_0_117701);
    
    HIEFFPLA_INST_0_50578 : MX2
      port map(A => 
        \U_ELK7_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]_net_1\, B => 
        \U_ELK7_CH/ELK_TX_DAT[4]\, S => 
        \U_ELK7_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_117930);
    
    \U_EXEC_MASTER/USB_MASTER_EN/TEST_SM[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117750, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_24, Q => 
        \U_EXEC_MASTER/USB_MASTER_EN/TEST_SM[3]_net_1\);
    
    HIEFFPLA_INST_0_54842 : NAND3B
      port map(A => HIEFFPLA_NET_0_117378, B => 
        HIEFFPLA_NET_0_117127, C => HIEFFPLA_NET_0_117180, Y => 
        HIEFFPLA_NET_0_117191);
    
    HIEFFPLA_INST_0_48286 : MX2
      port map(A => HIEFFPLA_NET_0_118354, B => 
        HIEFFPLA_NET_0_118351, S => \BIT_OS_SEL_3[0]\, Y => 
        \U_ELK16_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[6]\);
    
    \U50_PATTERNS/ELINK_DINA_2[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119771, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_9, Q => 
        \U50_PATTERNS/ELINK_DINA_2[4]\);
    
    HIEFFPLA_INST_0_56237 : AND2A
      port map(A => DCB_SALT_SEL_c, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/RECD_SER_WORD[1]_net_1\, 
        Y => \TFC_RX_SER_WORD[1]\);
    
    \U0_200M_BUF/\\\\INBUF_LVDS[0]\\\\/U0/U0\ : IOPADP_IN
      port map(N2PIN => 
        \U0_200M_BUF/\\\\INBUF_LVDS[0]\\\\/U0/U2_N2P\, PAD => 
        CLK200_P, Y => 
        \U0_200M_BUF/\\\\INBUF_LVDS[0]\\\\/U0/NET1\);
    
    \U_ELK9_CH/U_ELK1_SERDAT_SOURCE/SERDAT[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117830, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_7, Q => 
        \U_ELK9_CH/ELK_TX_DAT[3]\);
    
    \U_ELK8_CH/U_ELK1_CMD_TX/SER_OUT_FDEL\ : DFN1C0
      port map(D => \U_ELK8_CH/U_ELK1_CMD_TX/SER_OUT_FI_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_5, Q
         => \U_ELK8_CH/ELK_OUT_F\);
    
    HIEFFPLA_INST_0_60417 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_9[1]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_10[1]\, S
         => \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_1[0]\, Y
         => HIEFFPLA_NET_0_116269);
    
    HIEFFPLA_INST_0_61811 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_10[0]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_26[0]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_4[4]_net_1\, Y
         => HIEFFPLA_NET_0_116075);
    
    HIEFFPLA_INST_0_37223 : AOI1
      port map(A => \OP_MODE_c[2]\, B => HIEFFPLA_NET_0_120328, C
         => HIEFFPLA_NET_0_120320, Y => HIEFFPLA_NET_0_120321);
    
    \U50_PATTERNS/ELINK_ADDRA_10[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120086, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_22, Q => 
        \U50_PATTERNS/ELINK_ADDRA_10[1]\);
    
    HIEFFPLA_INST_0_42325 : NAND3B
      port map(A => \U50_PATTERNS/RD_USB_ADBUS[6]\, B => 
        HIEFFPLA_NET_0_119020, C => 
        \U50_PATTERNS/RD_USB_ADBUS[7]\, Y => 
        HIEFFPLA_NET_0_119571);
    
    HIEFFPLA_INST_0_51860 : AOI1D
      port map(A => HIEFFPLA_NET_0_117629, B => 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM_0[4]_net_1\, C => 
        HIEFFPLA_NET_0_117672, Y => HIEFFPLA_NET_0_117675);
    
    HIEFFPLA_INST_0_50720 : MX2
      port map(A => HIEFFPLA_NET_0_117912, B => 
        HIEFFPLA_NET_0_117909, S => \BIT_OS_SEL_4[1]\, Y => 
        HIEFFPLA_NET_0_117900);
    
    \U50_PATTERNS/ELINK_DINA_5[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119749, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_14, Q => 
        \U50_PATTERNS/ELINK_DINA_5[2]\);
    
    HIEFFPLA_INST_0_63238 : NAND2B
      port map(A => \OP_MODE_c_0[1]\, B => \PATT_TFC_DAT[1]\, Y
         => \U_TFC_SERDAT_SOURCE/N_SERDAT[1]\);
    
    HIEFFPLA_INST_0_52494 : MX2
      port map(A => HIEFFPLA_NET_0_117500, B => 
        HIEFFPLA_NET_0_117496, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_1[3]\, Y => 
        HIEFFPLA_NET_0_117556);
    
    \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[10]\ : DFN1C0
      port map(D => \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\);
    
    HIEFFPLA_INST_0_55188 : AND2A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[8]_net_1\, B => 
        HIEFFPLA_NET_0_115868, Y => HIEFFPLA_NET_0_117100);
    
    \U_ELK11_CH/U_ELK1_CMD_TX/SER_OUT_RDEL\ : DFN1C0
      port map(D => \U_ELK11_CH/U_ELK1_CMD_TX/SER_OUT_RI_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_16, Q
         => \U_ELK11_CH/ELK_OUT_R\);
    
    HIEFFPLA_INST_0_54213 : MX2
      port map(A => HIEFFPLA_NET_0_116361, B => 
        HIEFFPLA_NET_0_116555, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_1[3]_net_1\, Y
         => HIEFFPLA_NET_0_117294);
    
    \U_EXEC_MASTER/USB_MASTER_EN/T_CNT60M[4]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117739, CLK => CLK60MHZ, CLR
         => P_MASTER_POR_B_c_28, Q => 
        \U_EXEC_MASTER/USB_MASTER_EN/T_CNT60M[4]_net_1\);
    
    HIEFFPLA_INST_0_53981 : MX2
      port map(A => HIEFFPLA_NET_0_116223, B => 
        HIEFFPLA_NET_0_116109, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[3]_net_1\, Y
         => HIEFFPLA_NET_0_117324);
    
    HIEFFPLA_INST_0_161263 : DFN1C0
      port map(D => DCB_SALT_SEL_c, CLK => CCC_160M_ADJ, CLR => 
        P_MASTER_POR_B_c_31_0, Q => HIEFFPLA_NET_0_161292);
    
    HIEFFPLA_INST_0_43350 : MX2
      port map(A => \U50_PATTERNS/SM_BANK_SEL[10]\, B => 
        HIEFFPLA_NET_0_119227, S => HIEFFPLA_NET_0_118691, Y => 
        HIEFFPLA_NET_0_119321);
    
    HIEFFPLA_INST_0_51710 : NAND2B
      port map(A => 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM[4]_net_1\, B => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[31]_net_1\, Y => 
        HIEFFPLA_NET_0_117716);
    
    HIEFFPLA_INST_0_51095 : MX2
      port map(A => HIEFFPLA_NET_0_161291, B => 
        HIEFFPLA_NET_0_161290, S => HIEFFPLA_NET_0_161289, Y => 
        HIEFFPLA_NET_0_117836);
    
    HIEFFPLA_INST_0_50323 : MX2
      port map(A => 
        \U_ELK6_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[0]_net_1\, B => 
        \U_ELK6_CH/ELK_TX_DAT[2]\, S => 
        \U_ELK6_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_117976);
    
    HIEFFPLA_INST_0_46411 : AO1
      port map(A => HIEFFPLA_NET_0_119241, B => 
        \U50_PATTERNS/ELINK_DOUTA_1[7]\, C => 
        HIEFFPLA_NET_0_118846, Y => HIEFFPLA_NET_0_118696);
    
    HIEFFPLA_INST_0_46169 : AO1
      port map(A => HIEFFPLA_NET_0_119290, B => 
        \U50_PATTERNS/ELINK_DOUTA_17[3]\, C => 
        HIEFFPLA_NET_0_118750, Y => HIEFFPLA_NET_0_118751);
    
    HIEFFPLA_INST_0_43561 : NAND2B
      port map(A => \U50_PATTERNS/SM_BANK_SEL_0[21]\, B => 
        \U50_PATTERNS/SM_BANK_SEL[0]\, Y => HIEFFPLA_NET_0_119293);
    
    HIEFFPLA_INST_0_46234 : AO1A
      port map(A => HIEFFPLA_NET_0_118915, B => 
        \U50_PATTERNS/SM_BANK_SEL[0]\, C => HIEFFPLA_NET_0_118907, 
        Y => HIEFFPLA_NET_0_118735);
    
    \U_ELK15_CH/U_SLAVE_1ELK/RECD_SER_WORD[3]\ : DFN1C0
      port map(D => \U_ELK15_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[3]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_15[3]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_2[6]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117099, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_27_1, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_2[6]_net_1\);
    
    \U_ELK2_CH/U_SLAVE_1ELK/RECD_SER_WORD[5]\ : DFN1C0
      port map(D => \U_ELK2_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[5]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_2[5]\);
    
    \U50_PATTERNS/SM_BANK_SEL[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119311, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_7, Q => 
        \U50_PATTERNS/SM_BANK_SEL[1]\);
    
    HIEFFPLA_INST_0_49788 : MX2
      port map(A => HIEFFPLA_NET_0_118090, B => 
        HIEFFPLA_NET_0_118070, S => \BIT_OS_SEL_1[0]\, Y => 
        \U_ELK3_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[7]\);
    
    HIEFFPLA_INST_0_45372 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_7[2]\, C => 
        \U50_PATTERNS/SM_BANK_SEL[12]\, Y => 
        HIEFFPLA_NET_0_118927);
    
    HIEFFPLA_INST_0_56919 : NAND2A
      port map(A => HIEFFPLA_NET_0_116779, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_1[0]\, Y => 
        HIEFFPLA_NET_0_116775);
    
    HIEFFPLA_INST_0_39884 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_9[2]\, B => 
        HIEFFPLA_NET_0_119522, S => HIEFFPLA_NET_0_119292, Y => 
        HIEFFPLA_NET_0_119941);
    
    HIEFFPLA_INST_0_161264 : DFN1C0
      port map(D => 
        \U_ELK9_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_0, Q => 
        HIEFFPLA_NET_0_161291);
    
    \U_MASTER_DES/U13C_MASTER_DESER/Q[12]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[12]_net_1\, CLK => 
        CCC_160M_FXD, CLR => P_MASTER_POR_B_c_23, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/Q[12]_net_1\);
    
    HIEFFPLA_INST_0_40765 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_16[3]\, B => 
        HIEFFPLA_NET_0_119574, S => HIEFFPLA_NET_0_119257, Y => 
        HIEFFPLA_NET_0_119812);
    
    HIEFFPLA_INST_0_39911 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_9[5]\, B => 
        HIEFFPLA_NET_0_119518, S => HIEFFPLA_NET_0_119292, Y => 
        HIEFFPLA_NET_0_119938);
    
    \P_USB_MASTER_EN_pad/U0/U1\ : IOTRI_OB_EB
      port map(D => P_USB_MASTER_EN_c, E => \VCC\, DOUT => 
        \P_USB_MASTER_EN_pad/U0/NET1\, EOUT => 
        \P_USB_MASTER_EN_pad/U0/NET2\);
    
    \U_TFC_CMD_TX/CLK40M_GEN_DEL0\ : DFN1C0
      port map(D => CLK_40M_GL, CLK => CCC_160M_FXD, CLR => 
        MASTER_DCB_POR_B_i_0_i, Q => 
        \U_TFC_CMD_TX/CLK40M_GEN_DEL0_net_1\);
    
    \U_ELK2_CH/U_ELK1_SERDAT_SOURCE/SERDAT[7]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118141, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_13, Q => 
        \U_ELK2_CH/ELK_TX_DAT[7]\);
    
    \U_ELK4_CH/U_SLAVE_1ELK/RECD_SER_WORD[5]\ : DFN1C0
      port map(D => \U_ELK4_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[5]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_4[5]\);
    
    \U_ELK17_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]\ : DFN1C0
      port map(D => \U_ELK17_CH/U_SLAVE_1ELK/Q[4]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]_net_1\);
    
    \U50_PATTERNS/ELINK_RWA[12]/U1\ : DFN1P0
      port map(D => HIEFFPLA_NET_0_119708, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_11, Q => 
        \U50_PATTERNS/ELINK_RWA[12]\);
    
    HIEFFPLA_INST_0_49117 : AND2A
      port map(A => \OP_MODE_c_5[1]\, B => \PATT_ELK_DAT_1[4]\, Y
         => HIEFFPLA_NET_0_118189);
    
    HIEFFPLA_INST_0_62048 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_29[3]\, B => 
        HIEFFPLA_NET_0_117075, S => HIEFFPLA_NET_0_117072, Y => 
        HIEFFPLA_NET_0_116042);
    
    HIEFFPLA_INST_0_55612 : MX2
      port map(A => HIEFFPLA_NET_0_116194, B => 
        HIEFFPLA_NET_0_116085, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_1[3]\, Y => 
        HIEFFPLA_NET_0_117014);
    
    HIEFFPLA_INST_0_48214 : MX2
      port map(A => HIEFFPLA_NET_0_118364, B => 
        HIEFFPLA_NET_0_118362, S => \BIT_OS_SEL_1[1]\, Y => 
        HIEFFPLA_NET_0_118352);
    
    \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_115928, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_9, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/WAITCNT[2]\);
    
    \U50_PATTERNS/U4B_REGCROSS/SAMP_TWO[7]\ : DFN1C0
      port map(D => \U50_PATTERNS/U4B_REGCROSS/SAMP_ONE[7]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_29, Q => 
        \U50_PATTERNS/U4B_REGCROSS/SAMP_TWO[7]_net_1\);
    
    \U_ELK17_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL\ : DFN1C0
      port map(D => 
        \U_ELK17_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_0DEL_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL_net_1\);
    
    HIEFFPLA_INST_0_56786 : XA1B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_0[3]\, B => 
        HIEFFPLA_NET_0_116790, C => HIEFFPLA_NET_0_117085, Y => 
        HIEFFPLA_NET_0_116797);
    
    \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[4]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_WRD_40M_FIXED[4]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_27, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[4]_net_1\);
    
    HIEFFPLA_INST_0_52860 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_19[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_20[1]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_1[0]\, Y => 
        HIEFFPLA_NET_0_117499);
    
    HIEFFPLA_INST_0_48622 : NAND2B
      port map(A => \OP_MODE_c_2[1]\, B => \PATT_ELK_DAT_18[7]\, 
        Y => HIEFFPLA_NET_0_118276);
    
    \U_ELK14_CH/U_SLAVE_1ELK/Q[6]\ : DFN1C0
      port map(D => \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/Q[6]_net_1\);
    
    HIEFFPLA_INST_0_46514 : AND3B
      port map(A => \U50_PATTERNS/RD_USB_ADBUS[5]\, B => 
        \U50_PATTERNS/WR_XFER_TYPE[1]_net_1\, C => 
        \U50_PATTERNS/RD_USB_ADBUS[0]\, Y => 
        HIEFFPLA_NET_0_118675);
    
    \U_ELK5_CH/U_SLAVE_1ELK/RECD_SER_WORD[7]\ : DFN1C0
      port map(D => \U_ELK5_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[7]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_5[7]\);
    
    \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[1]\ : DFN1C0
      port map(D => 
        \U_ELK17_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_1DEL_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[1]_net_1\);
    
    HIEFFPLA_INST_0_49818 : MX2
      port map(A => \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\, 
        B => \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[14]_net_1\, S => 
        \BIT_OS_SEL_0[2]\, Y => HIEFFPLA_NET_0_118068);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_8[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116290, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_5, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_8[3]\);
    
    \U50_PATTERNS/RD_XFER_TYPE[6]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119543, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c, Q => 
        \U50_PATTERNS/RD_XFER_TYPE[6]_net_1\);
    
    HIEFFPLA_INST_0_54911 : AO1A
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_0[6]_net_1\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_0[8]_net_1\, C => 
        HIEFFPLA_NET_0_117171, Y => HIEFFPLA_NET_0_117172);
    
    HIEFFPLA_INST_0_40029 : MX2
      port map(A => HIEFFPLA_NET_0_119892, B => 
        \U50_PATTERNS/ELINK_BLKA[3]\, S => 
        \U50_PATTERNS/SM_BANK_SEL[20]\, Y => 
        HIEFFPLA_NET_0_119922);
    
    \U_EXEC_MASTER/MPOR_SALT_B_10\ : DFI1P0
      port map(D => HIEFFPLA_NET_0_117781, CLK => CLK_40M_GL, PRE
         => \U_EXEC_MASTER/SYNC_BRD_RST_BI_i_0_i_2\, QN => 
        MASTER_SALT_POR_B_i_0_i_10);
    
    \U_ELK1_CH/U_SLAVE_1ELK/RECD_SER_WORD[1]\ : DFN1C0
      port map(D => \U_ELK1_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[1]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_1[1]\);
    
    \U_ELK11_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]\ : DFN1C0
      port map(D => \U_ELK11_CH/U_SLAVE_1ELK/Q[4]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[4]_net_1\);
    
    HIEFFPLA_INST_0_62699 : AO13
      port map(A => HIEFFPLA_NET_0_115958, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_CLKPHASE[2]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_SEQCNT[3]\, Y => 
        HIEFFPLA_NET_0_115955);
    
    HIEFFPLA_INST_0_46676 : MX2
      port map(A => HIEFFPLA_NET_0_118621, B => 
        HIEFFPLA_NET_0_118635, S => \BIT_OS_SEL_5[1]\, Y => 
        HIEFFPLA_NET_0_118629);
    
    AFLSDF_INV_55 : INV
      port map(A => \U_ELK1_CH/U_DDR_ELK1/ELK_IN_DDR_F\, Y => 
        \AFLSDF_INV_55\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_CNT_6[6]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116626, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_12, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_6[6]\);
    
    HIEFFPLA_INST_0_46370 : AO1
      port map(A => HIEFFPLA_NET_0_119263, B => 
        \U50_PATTERNS/ELINK_DOUTA_8[7]\, C => 
        HIEFFPLA_NET_0_118704, Y => HIEFFPLA_NET_0_118705);
    
    HIEFFPLA_INST_0_37151 : XO1
      port map(A => HIEFFPLA_NET_0_120258, B => \TFC_ADDRB[4]\, C
         => \U200A_TFC/GP_PG_SM[10]_net_1\, Y => 
        HIEFFPLA_NET_0_120339);
    
    HIEFFPLA_INST_0_61859 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_27[2]\, B => 
        HIEFFPLA_NET_0_117131, S => HIEFFPLA_NET_0_117196, Y => 
        HIEFFPLA_NET_0_116068);
    
    HIEFFPLA_INST_0_54557 : AOI1B
      port map(A => HIEFFPLA_NET_0_117208, B => 
        HIEFFPLA_NET_0_116678, C => HIEFFPLA_NET_0_117263, Y => 
        HIEFFPLA_NET_0_117249);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_22[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116449, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_15, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_22[1]\);
    
    HIEFFPLA_INST_0_46497 : AND3C
      port map(A => \U50_PATTERNS/RD_USB_ADBUS[3]\, B => 
        HIEFFPLA_NET_0_119596, C => HIEFFPLA_NET_0_119571, Y => 
        HIEFFPLA_NET_0_118678);
    
    \U_ELK5_CH/U_SLAVE_1ELK/Q[3]\ : DFN1C0
      port map(D => \U_ELK5_CH/U_SLAVE_1ELK/ADJ_Q[3]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK5_CH/U_SLAVE_1ELK/Q[3]_net_1\);
    
    \U_ELK7_CH/U_SLAVE_1ELK/Q[14]\ : DFN1C0
      port map(D => \U_ELK7_CH/U_SLAVE_1ELK/ADJ_Q[14]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK7_CH/U_SLAVE_1ELK/Q[14]_net_1\);
    
    HIEFFPLA_INST_0_55098 : AO1
      port map(A => HIEFFPLA_NET_0_117126, B => 
        HIEFFPLA_NET_0_117588, C => HIEFFPLA_NET_0_117179, Y => 
        HIEFFPLA_NET_0_117122);
    
    HIEFFPLA_INST_0_41575 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_8[5]\, B => 
        HIEFFPLA_NET_0_119567, S => HIEFFPLA_NET_0_119291, Y => 
        HIEFFPLA_NET_0_119722);
    
    \U_ELK14_CH/U_ELK1_CMD_TX/SER_OUT_RDEL\ : DFN1C0
      port map(D => \U_ELK14_CH/U_ELK1_CMD_TX/SER_OUT_RI_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_12, Q
         => \U_ELK14_CH/ELK_OUT_R\);
    
    HIEFFPLA_INST_0_49103 : MX2
      port map(A => 
        \U_ELK1_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[1]_net_1\, B => 
        \U_ELK1_CH/ELK_TX_DAT[5]\, S => 
        \U_ELK1_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118196);
    
    HIEFFPLA_INST_0_62586 : MX2
      port map(A => HIEFFPLA_NET_0_117096, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_8[0]\, S => 
        HIEFFPLA_NET_0_117153, Y => HIEFFPLA_NET_0_115970);
    
    \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[2]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_WRD_40M_FIXED[2]_net_1\, 
        CLK => CLK_40M_GL, CLR => P_MASTER_POR_B_c_27, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[2]_net_1\);
    
    HIEFFPLA_INST_0_40158 : AOI1C
      port map(A => \U50_PATTERNS/ELINK_BLKA[6]\, B => 
        HIEFFPLA_NET_0_119641, C => HIEFFPLA_NET_0_119885, Y => 
        HIEFFPLA_NET_0_119886);
    
    \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[12]\ : DFN1C0
      port map(D => \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\, 
        CLK => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\);
    
    \U50_PATTERNS/ELINK_ADDRA_2[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119996, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_21, Q => 
        \U50_PATTERNS/ELINK_ADDRA_2[3]\);
    
    HIEFFPLA_INST_0_57165 : XA1B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_2[8]\, B => 
        HIEFFPLA_NET_0_116726, C => HIEFFPLA_NET_0_117179, Y => 
        HIEFFPLA_NET_0_116727);
    
    HIEFFPLA_INST_0_52938 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_31[2]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_0[2]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_3[0]\, Y => 
        HIEFFPLA_NET_0_117486);
    
    HIEFFPLA_INST_0_37763 : AO1
      port map(A => HIEFFPLA_NET_0_120223, B => 
        HIEFFPLA_NET_0_120203, C => HIEFFPLA_NET_0_120196, Y => 
        HIEFFPLA_NET_0_120213);
    
    \U_ELK5_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118021, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_5, Q => 
        \U_ELK5_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[1]_net_1\);
    
    HIEFFPLA_INST_0_63176 : AX1C
      port map(A => HIEFFPLA_NET_0_115869, B => 
        HIEFFPLA_NET_0_117225, C => HIEFFPLA_NET_0_117220, Y => 
        HIEFFPLA_NET_0_115868);
    
    HIEFFPLA_INST_0_55556 : MX2
      port map(A => HIEFFPLA_NET_0_116164, B => 
        HIEFFPLA_NET_0_116269, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_1[3]\, Y => 
        HIEFFPLA_NET_0_117021);
    
    HIEFFPLA_INST_0_47676 : MX2
      port map(A => \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[6]_net_1\, 
        B => \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[10]_net_1\, S => 
        \BIT_OS_SEL_2[2]\, Y => HIEFFPLA_NET_0_118448);
    
    HIEFFPLA_INST_0_47370 : AND2A
      port map(A => \OP_MODE_c_6[1]\, B => \PATT_ELK_DAT_13[0]\, 
        Y => HIEFFPLA_NET_0_118508);
    
    \U50_PATTERNS/U4C_REGCROSS/LOCAL_REG_VAL[1]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119111, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_21, Q => \ELKS_STRT_ADDR[1]\);
    
    HIEFFPLA_INST_0_57117 : AND3
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_2[5]\, B => 
        HIEFFPLA_NET_0_116736, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_2[6]\, Y => 
        HIEFFPLA_NET_0_116737);
    
    HIEFFPLA_INST_0_55514 : NAND3A
      port map(A => HIEFFPLA_NET_0_116971, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[0]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[3]\, Y => 
        HIEFFPLA_NET_0_117027);
    
    HIEFFPLA_INST_0_55400 : AO1
      port map(A => HIEFFPLA_NET_0_117087, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[2]\, C => 
        HIEFFPLA_NET_0_117038, Y => HIEFFPLA_NET_0_117043);
    
    HIEFFPLA_INST_0_50584 : MX2
      port map(A => 
        \U_ELK7_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[2]_net_1\, B => 
        \U_ELK7_CH/ELK_TX_DAT[6]\, S => 
        \U_ELK7_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_117929);
    
    \U_ELK13_CH/U_ELK1_CMD_TX/SER_OUT_FDEL\ : DFN1C0
      port map(D => \U_ELK13_CH/U_ELK1_CMD_TX/SER_OUT_FI_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_4, Q
         => \U_ELK13_CH/ELK_OUT_F\);
    
    \U200A_TFC/RX_SER_WORD_1DEL[3]\ : DFN1C0
      port map(D => \TFC_RX_SER_WORD[3]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_31, Q => 
        \U200A_TFC/RX_SER_WORD_1DEL[3]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/MAX_CNT[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_116948, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_16, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/MAX_CNT[6]\);
    
    \U50_PATTERNS/ELINKS_STOP_ADDR[4]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120123, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_14, Q => 
        \U50_PATTERNS/ELINKS_STOP_ADDR[4]\);
    
    HIEFFPLA_INST_0_60525 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_12[1]\, B => 
        HIEFFPLA_NET_0_117114, S => HIEFFPLA_NET_0_117133, Y => 
        HIEFFPLA_NET_0_116254);
    
    HIEFFPLA_INST_0_38037 : AO1A
      port map(A => \ELKS_STRT_ADDR[2]\, B => 
        HIEFFPLA_NET_0_120219, C => HIEFFPLA_NET_0_120167, Y => 
        HIEFFPLA_NET_0_120168);
    
    HIEFFPLA_INST_0_59644 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_2[0]\, B => 
        HIEFFPLA_NET_0_116680, S => HIEFFPLA_NET_0_117090, Y => 
        HIEFFPLA_NET_0_116367);
    
    HIEFFPLA_INST_0_58613 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_17[3]\, B => 
        HIEFFPLA_NET_0_116815, S => HIEFFPLA_NET_0_117161, Y => 
        HIEFFPLA_NET_0_116498);
    
    HIEFFPLA_INST_0_55997 : MX2
      port map(A => HIEFFPLA_NET_0_116959, B => 
        HIEFFPLA_NET_0_117036, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[4]\, Y => 
        HIEFFPLA_NET_0_116963);
    
    HIEFFPLA_INST_0_45346 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_18[3]\, C => 
        \U50_PATTERNS/SM_BANK_SEL[1]\, Y => HIEFFPLA_NET_0_118934);
    
    \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[10]\ : DFN1C0
      port map(D => \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[10]_net_1\);
    
    \U50_PATTERNS/U4E_REGCROSS/LOCAL_REG_VAL[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119065, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_6, Q => \OP_MODE_c[5]\);
    
    \U50_PATTERNS/U4A_REGCROSS/LOCAL_REG_VAL[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119147, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_17, Q => \TFC_STRT_ADDR[7]\);
    
    HIEFFPLA_INST_0_38114 : AX1C
      port map(A => \ELKS_ADDRB[2]\, B => HIEFFPLA_NET_0_120145, 
        C => \ELKS_ADDRB[3]\, Y => HIEFFPLA_NET_0_120149);
    
    \U_ELK6_CH/U_SLAVE_1ELK/Q[7]\ : DFN1C0
      port map(D => \U_ELK6_CH/U_SLAVE_1ELK/ADJ_Q[7]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/Q[7]_net_1\);
    
    HIEFFPLA_INST_0_48443 : MX2
      port map(A => HIEFFPLA_NET_0_118319, B => 
        HIEFFPLA_NET_0_118317, S => \BIT_OS_SEL_1[1]\, Y => 
        HIEFFPLA_NET_0_118310);
    
    \U_ELK15_CH/ELK_IN_R\ : DFN1C0
      port map(D => \U_ELK15_CH/ELK_IN_DDR_R\, CLK => 
        CCC_160M_ADJ, CLR => DEV_RST_B_c, Q => 
        \U_ELK15_CH/ELK_IN_R_net_1\);
    
    HIEFFPLA_INST_0_39785 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_7[7]\, B => 
        HIEFFPLA_NET_0_119516, S => HIEFFPLA_NET_0_119289, Y => 
        HIEFFPLA_NET_0_119952);
    
    HIEFFPLA_INST_0_38651 : MX2
      port map(A => HIEFFPLA_NET_0_119523, B => 
        \U50_PATTERNS/ELINK_ADDRA_11[1]\, S => 
        HIEFFPLA_NET_0_119280, Y => HIEFFPLA_NET_0_120078);
    
    \U_ELK17_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]\ : DFN1C0
      port map(D => \U_ELK17_CH/U_SLAVE_1ELK/Q[7]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]_net_1\);
    
    \U_ELK10_CH/U_SLAVE_1ELK/RECD_SER_WORD[2]\ : DFN1C0
      port map(D => \U_ELK10_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[2]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_10[2]\);
    
    HIEFFPLA_INST_0_58250 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_12[3]\, B => 
        HIEFFPLA_NET_0_116543, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_0[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116545);
    
    HIEFFPLA_INST_0_56457 : AOI1D
      port map(A => HIEFFPLA_NET_0_117432, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_SEL[3]_net_1\, C
         => \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[2]_net_1\, Y
         => HIEFFPLA_NET_0_116862);
    
    \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117718, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_31, Q => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[1]_net_1\);
    
    \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[7]\ : DFN1C0
      port map(D => 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[7]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\);
    
    HIEFFPLA_INST_0_57308 : XA1C
      port map(A => HIEFFPLA_NET_0_116716, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_3[5]\, C => 
        HIEFFPLA_NET_0_117179, Y => HIEFFPLA_NET_0_116702);
    
    \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[1]\ : DFN1C0
      port map(D => 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_BYTE[1]_net_1\);
    
    HIEFFPLA_INST_0_58966 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_21[3]\, B => 
        HIEFFPLA_NET_0_116815, S => HIEFFPLA_NET_0_117093, Y => 
        HIEFFPLA_NET_0_116453);
    
    HIEFFPLA_INST_0_43586 : NAND2B
      port map(A => \U50_PATTERNS/SM_BANK_SEL[21]\, B => 
        \U50_PATTERNS/SM_BANK_SEL[17]\, Y => 
        HIEFFPLA_NET_0_119278);
    
    \U50_PATTERNS/ELINK_BLKA[15]/U1\ : DFN1P0
      port map(D => HIEFFPLA_NET_0_119929, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_20, Q => 
        \U50_PATTERNS/ELINK_BLKA[15]\);
    
    HIEFFPLA_INST_0_43116 : AND2A
      port map(A => \U50_PATTERNS/REG_STATE[2]_net_1\, B => 
        \U50_PATTERNS/REG_STATE[0]_net_1\, Y => 
        HIEFFPLA_NET_0_119371);
    
    HIEFFPLA_INST_0_55262 : AO1C
      port map(A => HIEFFPLA_NET_0_117107, B => 
        HIEFFPLA_NET_0_117208, C => HIEFFPLA_NET_0_117086, Y => 
        HIEFFPLA_NET_0_117074);
    
    HIEFFPLA_INST_0_37702 : AO1C
      port map(A => \U200B_ELINKS/GP_PG_SM[0]_net_1\, B => 
        HIEFFPLA_NET_0_120188, C => \OP_MODE_c[6]\, Y => 
        HIEFFPLA_NET_0_120225);
    
    HIEFFPLA_INST_0_56913 : NAND3A
      port map(A => HIEFFPLA_NET_0_116775, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_1[5]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_1[4]\, Y => 
        HIEFFPLA_NET_0_116777);
    
    \U_ELK5_CH/U_SLAVE_1ELK/RECD_SER_WORD[1]\ : DFN1C0
      port map(D => \U_ELK5_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[1]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_5[1]\);
    
    \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[0]\ : DFN1C0
      port map(D => 
        \U_ELK12_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/Q[8]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/ADJ_Q[8]_net_1\, CLK => 
        CCC_160M_FXD, CLR => P_MASTER_POR_B_c_34, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/Q[8]_net_1\);
    
    HIEFFPLA_INST_0_55866 : MX2
      port map(A => HIEFFPLA_NET_0_116002, B => 
        HIEFFPLA_NET_0_116258, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[3]\, Y => 
        HIEFFPLA_NET_0_116980);
    
    \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_2S_16\ : DFN1C0
      port map(D => 
        \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_1S_0_net_1\, CLK
         => CLK60MHZ, CLR => \U_EXEC_MASTER/P_MASTER_POR_B_c_0\, 
        Q => P_USB_MASTER_EN_c_16);
    
    HIEFFPLA_INST_0_59612 : MX2
      port map(A => HIEFFPLA_NET_0_116677, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_29[1]\, S => 
        HIEFFPLA_NET_0_117395, Y => HIEFFPLA_NET_0_116370);
    
    HIEFFPLA_INST_0_56153 : NAND2A
      port map(A => HIEFFPLA_NET_0_116942, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/MAX_CNT[3]\, Y => 
        HIEFFPLA_NET_0_116941);
    
    HIEFFPLA_INST_0_56711 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_0[8]\, B => 
        HIEFFPLA_NET_0_116792, S => HIEFFPLA_NET_0_117602, Y => 
        HIEFFPLA_NET_0_116816);
    
    \U200B_ELINKS/RX_SER_WORD_3DEL[2]\ : DFN1P0
      port map(D => \AFLSDF_INV_67\, CLK => CLK_40M_GL, PRE => 
        P_MASTER_POR_B_c_31_0, Q => 
        \U200B_ELINKS/RX_SER_WORD_3DEL_i_0[2]\);
    
    HIEFFPLA_INST_0_44392 : MX2
      port map(A => \TFC_STOP_ADDR[6]\, B => 
        \U50_PATTERNS/U4B_REGCROSS/SAMP_TWO[6]_net_1\, S => 
        HIEFFPLA_NET_0_119135, Y => HIEFFPLA_NET_0_119127);
    
    HIEFFPLA_INST_0_45416 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_15[7]\, C => 
        \U50_PATTERNS/SM_BANK_SEL[4]\, Y => HIEFFPLA_NET_0_118917);
    
    HIEFFPLA_INST_0_44928 : AND2B
      port map(A => \U50_PATTERNS/REG_STATE[3]_net_1\, B => 
        \U50_PATTERNS/USB_RXF_B\, Y => HIEFFPLA_NET_0_119016);
    
    HIEFFPLA_INST_0_37746 : AND3C
      port map(A => HIEFFPLA_NET_0_120234, B => 
        \U200B_ELINKS/GP_PG_SM[0]_net_1\, C => 
        HIEFFPLA_NET_0_120231, Y => HIEFFPLA_NET_0_120218);
    
    HIEFFPLA_INST_0_40486 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_12[4]\, B => 
        HIEFFPLA_NET_0_119570, S => HIEFFPLA_NET_0_119295, Y => 
        HIEFFPLA_NET_0_119843);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_2[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116034, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_10, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_2[1]\);
    
    \U_ELK16_CH/U_SLAVE_1ELK/RECD_SER_WORD[7]\ : DFN1C0
      port map(D => \U_ELK16_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[7]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_16[7]\);
    
    HIEFFPLA_INST_0_54792 : MX2
      port map(A => HIEFFPLA_NET_0_116184, B => 
        HIEFFPLA_NET_0_116073, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[3]_net_1\, Y => 
        HIEFFPLA_NET_0_117199);
    
    HIEFFPLA_INST_0_50196 : MX2
      port map(A => \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[7]_net_1\, B
         => \U_ELK5_CH/U_SLAVE_1ELK/ARB_BYTE[11]_net_1\, S => 
        \BIT_OS_SEL_6[2]\, Y => HIEFFPLA_NET_0_117994);
    
    HIEFFPLA_INST_0_40225 : NAND3C
      port map(A => HIEFFPLA_NET_0_119389, B => 
        HIEFFPLA_NET_0_119464, C => \U50_PATTERNS/SM_BANK_SEL[0]\, 
        Y => HIEFFPLA_NET_0_119873);
    
    \U50_PATTERNS/U3_USB_DAT_BUS/_BIBUF_F_24U[7]_/U0/U1\ : 
        IOBI_IRC_OB_EB
      port map(D => \U50_PATTERNS/WR_USB_ADBUS[7]\, CLR => 
        \AFLSDF_INV_11\, E => \U50_PATTERNS/TrienAux\, ICLK => 
        CLK60MHZ, YIN => 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[7]\\\\/U0/NET3\, 
        DOUT => 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[7]\\\\/U0/NET1\, 
        EOUT => 
        \U50_PATTERNS/U3_USB_DAT_BUS/\\\\BIBUF_F_24U[7]\\\\/U0/NET2\, 
        Y => \U50_PATTERNS/RD_USB_ADBUS[7]\);
    
    HIEFFPLA_INST_0_56261 : NAND3C
      port map(A => HIEFFPLA_NET_0_116880, B => 
        HIEFFPLA_NET_0_116888, C => HIEFFPLA_NET_0_116896, Y => 
        HIEFFPLA_NET_0_116904);
    
    HIEFFPLA_INST_0_111893 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_4[1]\, C => 
        \U50_PATTERNS/SM_BANK_SEL[15]\, Y => 
        HIEFFPLA_NET_0_115826);
    
    \U50_PATTERNS/ELINK_ADDRA_5[0]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119975, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_3, Q => 
        \U50_PATTERNS/ELINK_ADDRA_5[0]\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_19[0]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116180, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_10, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_19[0]\);
    
    \U_DDR_ELK0/BIBUF_LVDS_0/U0/U0\ : IOPADP_BI
      port map(N2PIN => \U_DDR_ELK0/BIBUF_LVDS_0/U0/U2_N2P\, D
         => \U_DDR_ELK0/BIBUF_LVDS_0/U0/NET1\, E => 
        \U_DDR_ELK0/BIBUF_LVDS_0/U0/NET2\, PAD => ELK0_DAT_P, Y
         => \U_DDR_ELK0/BIBUF_LVDS_0/U0/NET4\);
    
    HIEFFPLA_INST_0_42669 : NAND3C
      port map(A => HIEFFPLA_NET_0_118998, B => 
        HIEFFPLA_NET_0_119462, C => HIEFFPLA_NET_0_119391, Y => 
        HIEFFPLA_NET_0_119487);
    
    \U50_PATTERNS/SM_BANK_SEL[8]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119302, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_8, Q => 
        \U50_PATTERNS/SM_BANK_SEL[8]\);
    
    HIEFFPLA_INST_0_42434 : AND2
      port map(A => HIEFFPLA_NET_0_119473, B => 
        \U50_PATTERNS/RD_XFER_TYPE[7]_net_1\, Y => 
        HIEFFPLA_NET_0_119534);
    
    HIEFFPLA_INST_0_41215 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_3[5]\, B => 
        HIEFFPLA_NET_0_119567, S => HIEFFPLA_NET_0_119247, Y => 
        HIEFFPLA_NET_0_119762);
    
    \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[14]\ : DFN1C0
      port map(D => \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[12]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/ADJ_Q[14]_net_1\);
    
    HIEFFPLA_INST_0_59905 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_3[3]\, B => 
        HIEFFPLA_NET_0_116330, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_2[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116336);
    
    HIEFFPLA_INST_0_45313 : AO1
      port map(A => HIEFFPLA_NET_0_119250, B => 
        \U50_PATTERNS/ELINK_DOUTA_5[4]\, C => 
        HIEFFPLA_NET_0_118943, Y => HIEFFPLA_NET_0_118944);
    
    \U200B_ELINKS/ADDR_POINTER_0[4]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120164, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_32_0, Q => \ELKS_ADDRB_0[4]\);
    
    HIEFFPLA_INST_0_37548 : OA1A
      port map(A => HIEFFPLA_NET_0_120334, B => 
        \U200A_TFC/GP_PG_SM[10]_net_1\, C => \TFC_ADDRB[0]\, Y
         => HIEFFPLA_NET_0_120262);
    
    HIEFFPLA_INST_0_60516 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_12[0]\, B => 
        HIEFFPLA_NET_0_117096, S => HIEFFPLA_NET_0_117133, Y => 
        HIEFFPLA_NET_0_116255);
    
    HIEFFPLA_INST_0_60209 : MX2
      port map(A => HIEFFPLA_NET_0_116687, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_7[2]\, S => 
        HIEFFPLA_NET_0_117212, Y => HIEFFPLA_NET_0_116295);
    
    \U_ELK2_CH/U_SLAVE_1ELK/Q[9]\ : DFN1C0
      port map(D => \U_ELK2_CH/U_SLAVE_1ELK/ADJ_Q[9]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/Q[9]_net_1\);
    
    HIEFFPLA_INST_0_57972 : NAND3C
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_7[6]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_7[5]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_7[4]\, Y => 
        HIEFFPLA_NET_0_116587);
    
    \U_ELK3_CH/U_SLAVE_1ELK/Q[2]\ : DFN1C0
      port map(D => \U_ELK3_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/Q[2]_net_1\);
    
    HIEFFPLA_INST_0_52152 : NAND2A
      port map(A => HIEFFPLA_NET_0_117689, B => 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM[5]_net_1\, Y => 
        HIEFFPLA_NET_0_117623);
    
    HIEFFPLA_INST_0_45655 : AO1A
      port map(A => HIEFFPLA_NET_0_119475, B => 
        \U50_PATTERNS/ELINKS_STOP_ADDR[0]\, C => 
        HIEFFPLA_NET_0_118773, Y => HIEFFPLA_NET_0_118871);
    
    HIEFFPLA_INST_0_48417 : MX2
      port map(A => \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\, 
        B => \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\, S => 
        \BIT_OS_SEL_0[2]\, Y => HIEFFPLA_NET_0_118314);
    
    \U_ELK8_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]\ : DFN1C0
      port map(D => \U_ELK8_CH/U_SLAVE_1ELK/Q[5]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK8_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]_net_1\);
    
    HIEFFPLA_INST_0_59507 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_28[1]\, B => 
        HIEFFPLA_NET_0_116677, S => HIEFFPLA_NET_0_117094, Y => 
        HIEFFPLA_NET_0_116385);
    
    \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_SEL[0]\ : DFN1C0
      port map(D => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_BIT_OS_VAL[0]\, CLK
         => CLK_40M_GL, CLR => P_MASTER_POR_B_c_27_1, Q => 
        \BIT_OS_SEL[0]\);
    
    HIEFFPLA_INST_0_43555 : NAND2B
      port map(A => \U50_PATTERNS/SM_BANK_SEL_0[21]\, B => 
        \U50_PATTERNS/SM_BANK_SEL[4]\, Y => HIEFFPLA_NET_0_119297);
    
    \U_ELK10_CH/U_ELK1_CMD_TX/SER_OUT_FDEL\ : DFN1C0
      port map(D => \U_ELK10_CH/U_ELK1_CMD_TX/SER_OUT_FI_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_8, Q
         => \U_ELK10_CH/ELK_OUT_F\);
    
    HIEFFPLA_INST_0_56453 : AOI1D
      port map(A => HIEFFPLA_NET_0_117432, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_SEL[3]_net_1\, C
         => \U_MASTER_DES/U13C_MASTER_DESER/ARB_BYTE[0]_net_1\, Y
         => HIEFFPLA_NET_0_116864);
    
    \U_ELK12_CH/U_SLAVE_1ELK/Q[0]\ : DFN1C0
      port map(D => \U_ELK12_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK12_CH/U_SLAVE_1ELK/Q[0]_net_1\);
    
    HIEFFPLA_INST_0_48617 : NAND2B
      port map(A => \OP_MODE_c_1[1]\, B => \PATT_ELK_DAT_18[2]\, 
        Y => HIEFFPLA_NET_0_118281);
    
    HIEFFPLA_INST_0_37021 : AOI1A
      port map(A => HIEFFPLA_NET_0_120353, B => 
        HIEFFPLA_NET_0_120325, C => HIEFFPLA_NET_0_120367, Y => 
        HIEFFPLA_NET_0_120368);
    
    HIEFFPLA_INST_0_43027 : AO1D
      port map(A => HIEFFPLA_NET_0_119328, B => 
        HIEFFPLA_NET_0_119376, C => HIEFFPLA_NET_0_119430, Y => 
        HIEFFPLA_NET_0_119398);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_2[4]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116031, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_10, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_2[4]\);
    
    \U50_PATTERNS/ELINK_ADDRA_14[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120052, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_5, Q => 
        \U50_PATTERNS/ELINK_ADDRA_14[3]\);
    
    HIEFFPLA_INST_0_45913 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_12[0]\, C => 
        \U50_PATTERNS/SM_BANK_SEL[7]\, Y => HIEFFPLA_NET_0_118812);
    
    \U_ELK4_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118064, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_1, Q => 
        \U_ELK4_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_14[1]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116527, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_13, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_14[1]\);
    
    HIEFFPLA_INST_0_57731 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_6[3]\, B => 
        HIEFFPLA_NET_0_116613, S => HIEFFPLA_NET_0_117599, Y => 
        HIEFFPLA_NET_0_116629);
    
    HIEFFPLA_INST_0_57494 : XA1B
      port map(A => HIEFFPLA_NET_0_116671, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_4[2]\, C => 
        HIEFFPLA_NET_0_117179, Y => HIEFFPLA_NET_0_116669);
    
    HIEFFPLA_INST_0_42880 : NAND2B
      port map(A => \U50_PATTERNS/REG_STATE[5]_net_1\, B => 
        \U50_PATTERNS/REG_STATE[1]_net_1\, Y => 
        HIEFFPLA_NET_0_119438);
    
    HIEFFPLA_INST_0_54418 : MX2
      port map(A => HIEFFPLA_NET_0_116334, B => 
        HIEFFPLA_NET_0_116389, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[3]_net_1\, Y => 
        HIEFFPLA_NET_0_117268);
    
    HIEFFPLA_INST_0_37672 : NAND2B
      port map(A => \U200B_ELINKS/GP_PG_SM[0]_net_1\, B => 
        \U200B_ELINKS/GP_PG_SM[1]_net_1\, Y => 
        HIEFFPLA_NET_0_120235);
    
    HIEFFPLA_INST_0_56759 : NAND3A
      port map(A => HIEFFPLA_NET_0_116802, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_0[0]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_0[4]\, Y => 
        HIEFFPLA_NET_0_116805);
    
    HIEFFPLA_INST_0_46096 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_15[4]\, C => 
        \U50_PATTERNS/SM_BANK_SEL[4]\, Y => HIEFFPLA_NET_0_118767);
    
    HIEFFPLA_INST_0_49290 : MX2
      port map(A => HIEFFPLA_NET_0_118184, B => 
        HIEFFPLA_NET_0_118160, S => \BIT_OS_SEL_2[0]\, Y => 
        \U_ELK1_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[7]\);
    
    HIEFFPLA_INST_0_44929 : AND2A
      port map(A => \U50_PATTERNS/REG_STATE[4]_net_1\, B => 
        \U50_PATTERNS/USB_RXF_B\, Y => HIEFFPLA_NET_0_119015);
    
    HIEFFPLA_INST_0_40279 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_0[5]\, B => 
        HIEFFPLA_NET_0_119567, S => HIEFFPLA_NET_0_119272, Y => 
        HIEFFPLA_NET_0_119866);
    
    \U50_PATTERNS/U4D_REGCROSS/SAMP_ONE[0]\ : DFN1C0
      port map(D => \U50_PATTERNS/ELINKS_STOP_ADDR[0]\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_25, Q => 
        \U50_PATTERNS/U4D_REGCROSS/SAMP_ONE[0]_net_1\);
    
    HIEFFPLA_INST_0_39794 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_8[0]\, B => 
        HIEFFPLA_NET_0_119524, S => HIEFFPLA_NET_0_119291, Y => 
        HIEFFPLA_NET_0_119951);
    
    \U_ELK19_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]\ : DFN1C0
      port map(D => \U_ELK19_CH/U_SLAVE_1ELK/Q[12]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK19_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]_net_1\);
    
    HIEFFPLA_INST_0_49959 : MX2
      port map(A => \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[9]_net_1\, B
         => \U_ELK4_CH/U_SLAVE_1ELK/ARB_BYTE[13]_net_1\, S => 
        \BIT_OS_SEL_7[2]\, Y => HIEFFPLA_NET_0_118037);
    
    HIEFFPLA_INST_0_60875 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_17[1]\, B => 
        HIEFFPLA_NET_0_117167, S => HIEFFPLA_NET_0_117169, Y => 
        HIEFFPLA_NET_0_116204);
    
    HIEFFPLA_INST_0_51606 : MX2
      port map(A => 
        \U_EXEC_MASTER/USB_MASTER_EN/CNT_EN_60M2S_net_1\, B => 
        \U_EXEC_MASTER/USB_MASTER_EN/T_CNT60M[1]_net_1\, S => 
        HIEFFPLA_NET_0_117753, Y => HIEFFPLA_NET_0_117735);
    
    HIEFFPLA_INST_0_44038 : MX2
      port map(A => \U50_PATTERNS/TFC_STOP_ADDR[7]\, B => 
        \U50_PATTERNS/TFC_STOP_ADDR_T[7]\, S => 
        HIEFFPLA_NET_0_119472, Y => HIEFFPLA_NET_0_119181);
    
    \U_ELK6_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117974, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_9, Q => 
        \U_ELK6_CH/U_ELK1_CMD_TX/SER_CMD_WORD_F[3]_net_1\);
    
    HIEFFPLA_INST_0_39659 : MX2
      port map(A => \U50_PATTERNS/ELINK_ADDRA_6[1]\, B => 
        HIEFFPLA_NET_0_119523, S => HIEFFPLA_NET_0_119258, Y => 
        HIEFFPLA_NET_0_119966);
    
    \U_ELK18_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118286, CLK => CCC_160M_FXD, 
        CLR => MASTER_SALT_POR_B_i_0_i_0, Q => 
        \U_ELK18_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]_net_1\);
    
    HIEFFPLA_INST_0_51717 : NAND2B
      port map(A => 
        \U_MASTER_DES/U13A_ADJ_160M/SHIFT_SM[4]_net_1\, B => 
        \U_MASTER_DES/U13A_ADJ_160M/ALL81BITS[44]_net_1\, Y => 
        HIEFFPLA_NET_0_117709);
    
    HIEFFPLA_INST_0_41916 : NAND2B
      port map(A => \U50_PATTERNS/ELINK_RWA[10]\, B => 
        HIEFFPLA_NET_0_119662, Y => HIEFFPLA_NET_0_119663);
    
    HIEFFPLA_INST_0_54293 : MX2
      port map(A => HIEFFPLA_NET_0_116149, B => 
        HIEFFPLA_NET_0_116049, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_2[3]_net_1\, Y
         => HIEFFPLA_NET_0_117284);
    
    HIEFFPLA_INST_0_44222 : MX2
      port map(A => \U50_PATTERNS/TFC_STRT_ADDR_T[6]\, B => 
        \U50_PATTERNS/RD_USB_ADBUS[6]\, S => 
        HIEFFPLA_NET_0_119491, Y => HIEFFPLA_NET_0_119158);
    
    \U50_PATTERNS/ELINK_DINA_7[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119728, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_17, Q => 
        \U50_PATTERNS/ELINK_DINA_7[7]\);
    
    HIEFFPLA_INST_0_55095 : AOI1D
      port map(A => HIEFFPLA_NET_0_116768, B => 
        HIEFFPLA_NET_0_117370, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[6]_net_1\, Y => 
        HIEFFPLA_NET_0_117123);
    
    \U_ELK9_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0\ : DFN1C0
      port map(D => CLK_40M_GL, CLK => CCC_160M_FXD, CLR => 
        MASTER_SALT_POR_B_i_0_i_12, Q => 
        \U_ELK9_CH/U_ELK1_CMD_TX/CLK40M_GEN_DEL0_net_1\);
    
    \U200A_TFC/RX_SER_WORD_1DEL[0]\ : DFN1C0
      port map(D => \TFC_RX_SER_WORD[0]\, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_30, Q => 
        \U200A_TFC/RX_SER_WORD_1DEL[0]_net_1\);
    
    \U_ELK5_CH/U_ELK1_CMD_TX/SER_OUT_RDEL\ : DFN1C0
      port map(D => \U_ELK5_CH/U_ELK1_CMD_TX/SER_OUT_RI_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_SALT_POR_B_i_0_i_5, Q
         => \U_ELK5_CH/ELK_OUT_R\);
    
    \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[6]\ : DFN1C0
      port map(D => \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[4]_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\);
    
    \U50_PATTERNS/ELINKS_STRT_ADDR_T[3]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120100, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_21, Q => 
        \U50_PATTERNS/ELINKS_STRT_ADDR_T[3]\);
    
    \U50_PATTERNS/TFC_ADDRA[6]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119201, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_10, Q => 
        \U50_PATTERNS/TFC_ADDRA[6]\);
    
    AFLSDF_INV_22 : INV
      port map(A => DCB_SALT_SEL_c, Y => \AFLSDF_INV_22\);
    
    \U_ELK13_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]\ : DFN1C0
      port map(D => \U_ELK13_CH/U_SLAVE_1ELK/Q[2]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK13_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[2]_net_1\);
    
    HIEFFPLA_INST_0_46575 : AND2
      port map(A => CLK_40M_GL, B => 
        \U_ELK0_CMD_TX/CLK40M_GEN_DEL0_net_1\, Y => 
        HIEFFPLA_NET_0_118661);
    
    \U50_PATTERNS/ELINK_DINA_7[2]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119733, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_17, Q => 
        \U50_PATTERNS/ELINK_DINA_7[2]\);
    
    HIEFFPLA_INST_0_37782 : NAND2
      port map(A => HIEFFPLA_NET_0_120223, B => 
        \U200B_ELINKS/GP_PG_SM[7]_net_1\, Y => 
        HIEFFPLA_NET_0_120208);
    
    HIEFFPLA_INST_0_37778 : AND3A
      port map(A => HIEFFPLA_NET_0_120201, B => 
        \U200B_ELINKS/GP_PG_SM[8]_net_1\, C => 
        HIEFFPLA_NET_0_120218, Y => HIEFFPLA_NET_0_120210);
    
    HIEFFPLA_INST_0_111416 : MX2
      port map(A => HIEFFPLA_NET_0_116735, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_13[0]\, S => 
        HIEFFPLA_NET_0_117396, Y => HIEFFPLA_NET_0_116531);
    
    \U_ELK1_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL\ : DFN1C0
      port map(D => \U_ELK1_CH/ELK_IN_F_net_1\, CLK => 
        CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK1_CH/U_SLAVE_1ELK/ADJ_SER_IN_F_0DEL_net_1\);
    
    HIEFFPLA_INST_0_61868 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_27[3]\, B => 
        HIEFFPLA_NET_0_117075, S => HIEFFPLA_NET_0_117196, Y => 
        HIEFFPLA_NET_0_116067);
    
    HIEFFPLA_INST_0_61568 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_23[2]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_24[2]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[0]\, Y => 
        HIEFFPLA_NET_0_116108);
    
    \U_EXEC_MASTER/USB_MASTER_EN/T_CNT60M[7]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117736, CLK => CLK60MHZ, CLR
         => P_MASTER_POR_B_c_29, Q => 
        \U_EXEC_MASTER/USB_MASTER_EN/T_CNT60M[7]_net_1\);
    
    \U_ELK6_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]\ : DFN1C0
      port map(D => \U_ELK6_CH/U_SLAVE_1ELK/Q[12]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK6_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[12]_net_1\);
    
    HIEFFPLA_INST_0_42740 : AND3A
      port map(A => \U50_PATTERNS/REG_STATE_0[2]_net_1\, B => 
        \U50_PATTERNS/REG_STATE_0[5]_net_1\, C => 
        \U50_PATTERNS/REG_STATE_0[1]_net_1\, Y => 
        HIEFFPLA_NET_0_119471);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.SEQCNTS_22[3]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116127, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_5, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_22[3]\);
    
    HIEFFPLA_INST_0_38235 : AND2A
      port map(A => HIEFFPLA_NET_0_119452, B => 
        \U50_PATTERNS/RD_USB_ADBUS[6]\, Y => 
        HIEFFPLA_NET_0_120129);
    
    \U200B_ELINKS/LOC_STRT_ADDR[5]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120174, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_11, Q => 
        \U200B_ELINKS/LOC_STRT_ADDR[5]\);
    
    \U50_PATTERNS/ELINK_BLKA[6]/U1\ : DFN1P0
      port map(D => HIEFFPLA_NET_0_119919, CLK => CLK60MHZ, PRE
         => P_USB_MASTER_EN_c_19, Q => 
        \U50_PATTERNS/ELINK_BLKA[6]\);
    
    \U_ELK9_CH/U_SLAVE_1ELK/RECD_SER_WORD[3]\ : DFN1C0
      port map(D => \U_ELK9_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[3]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_9[3]\);
    
    \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[0]\ : DFN1C0
      port map(D => 
        \U_ELK17_CH/U_SLAVE_1ELK/ADJ_SER_IN_R_1DEL_net_1\, CLK
         => CCC_160M_ADJ, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/ADJ_Q[0]_net_1\);
    
    HIEFFPLA_INST_0_58497 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_31[2]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_15[2]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_3[4]_net_1\, Y
         => HIEFFPLA_NET_0_116514);
    
    HIEFFPLA_INST_0_45517 : AND3A
      port map(A => HIEFFPLA_NET_0_119437, B => 
        \U50_PATTERNS/WR_XFER_TYPE[7]_net_1\, C => 
        HIEFFPLA_NET_0_119367, Y => HIEFFPLA_NET_0_118898);
    
    HIEFFPLA_INST_0_42841 : NAND2B
      port map(A => \U50_PATTERNS/REG_STATE[1]_net_1\, B => 
        \U50_PATTERNS/REG_STATE[3]_net_1\, Y => 
        HIEFFPLA_NET_0_119451);
    
    HIEFFPLA_INST_0_54426 : MX2
      port map(A => HIEFFPLA_NET_0_117294, B => 
        HIEFFPLA_NET_0_117276, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[2]_net_1\, Y => 
        HIEFFPLA_NET_0_117267);
    
    HIEFFPLA_INST_0_53038 : MX2
      port map(A => HIEFFPLA_NET_0_117453, B => 
        HIEFFPLA_NET_0_117565, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[2]\, Y => 
        HIEFFPLA_NET_0_117473);
    
    HIEFFPLA_INST_0_59456 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_27[2]\, B => 
        HIEFFPLA_NET_0_116687, S => HIEFFPLA_NET_0_117162, Y => 
        HIEFFPLA_NET_0_116392);
    
    HIEFFPLA_INST_0_58682 : NOR3A
      port map(A => HIEFFPLA_NET_0_116482, B => 
        HIEFFPLA_NET_0_116485, C => HIEFFPLA_NET_0_116487, Y => 
        HIEFFPLA_NET_0_116488);
    
    \U_MASTER_DES/U13C_MASTER_DESER/CONFIG_ONCE_TRIG\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_117193, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_24, Q => 
        \U_MASTER_DES/CCC2_CONFIG_TRIG\);
    
    \U_ELK11_CH/U_SLAVE_1ELK/Q[8]\ : DFN1C0
      port map(D => \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/Q[8]_net_1\);
    
    HIEFFPLA_INST_0_54660 : MX2
      port map(A => HIEFFPLA_NET_0_117320, B => 
        HIEFFPLA_NET_0_117224, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE[0]_net_1\, Y => 
        HIEFFPLA_NET_0_117226);
    
    HIEFFPLA_INST_0_51180 : MX2
      port map(A => \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\, B
         => \U_ELK9_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\, S => 
        \BIT_OS_SEL_2[2]\, Y => HIEFFPLA_NET_0_117816);
    
    \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[1]\ : DFN1C0
      port map(D => 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[1]_net_1\);
    
    \U_MASTER_DES/U13C_MASTER_DESER/REG40M.BIT_OS_VAL_2[2]/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_116365, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_18, Q => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_2[2]\);
    
    \U_ELK16_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]\ : DFN1C0
      port map(D => \U_ELK16_CH/U_SLAVE_1ELK/Q[1]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK16_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[1]_net_1\);
    
    \U_ELK9_CH/U_SLAVE_1ELK/RECD_SER_WORD[4]\ : DFN1C0
      port map(D => \U_ELK9_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[4]\, 
        CLK => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \ELK_RX_SER_WORD_9[4]\);
    
    \U_ELK14_CH/U_SLAVE_1ELK/Q[8]\ : DFN1C0
      port map(D => \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[8]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/Q[8]_net_1\);
    
    HIEFFPLA_INST_0_58193 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_11[2]\, B => 
        HIEFFPLA_NET_0_116550, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM_0[6]_net_1\, Y => 
        HIEFFPLA_NET_0_116552);
    
    HIEFFPLA_INST_0_55636 : MX2
      port map(A => HIEFFPLA_NET_0_115987, B => 
        HIEFFPLA_NET_0_116238, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_1[3]\, Y => 
        HIEFFPLA_NET_0_117011);
    
    \U50_PATTERNS/ELINK_ADDRA_7[7]/U1\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_119952, CLK => CLK60MHZ, CLR
         => P_USB_MASTER_EN_c_6, Q => 
        \U50_PATTERNS/ELINK_ADDRA_7[7]\);
    
    HIEFFPLA_INST_0_55360 : AOI1
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[8]_net_1\, B => 
        \OP_MODE_c[5]\, C => 
        \U_MASTER_DES/U13C_MASTER_DESER/DES_SM[2]_net_1\, Y => 
        HIEFFPLA_NET_0_117051);
    
    HIEFFPLA_INST_0_111316 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_26[0]\, B => 
        HIEFFPLA_NET_0_116735, S => HIEFFPLA_NET_0_117337, Y => 
        HIEFFPLA_NET_0_116396);
    
    \U_ELK9_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]\ : DFN1C0
      port map(D => \U_ELK9_CH/U_SLAVE_1ELK/Q[11]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK9_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]_net_1\);
    
    \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[11]\ : DFN1C0
      port map(D => 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[11]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK3_CH/U_SLAVE_1ELK/ARB_BYTE[11]_net_1\);
    
    \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_2S_17\ : DFN1C0
      port map(D => 
        \U_EXEC_MASTER/USB_MASTER_EN/USB_EN_60M_1S_0_net_1\, CLK
         => CLK60MHZ, CLR => \U_EXEC_MASTER/P_MASTER_POR_B_c_0\, 
        Q => P_USB_MASTER_EN_c_17);
    
    \U_ELK5_CH/U_ELK1_SERDAT_SOURCE/SERDAT[1]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_118012, CLK => CLK_40M_GL, CLR
         => MASTER_SALT_POR_B_i_0_i_17, Q => 
        \U_ELK5_CH/ELK_TX_DAT[1]\);
    
    \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[8]\ : DFN1C0
      port map(D => 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK2_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\);
    
    \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[8]\ : DFN1C0
      port map(D => 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK17_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\);
    
    \U_ELK14_CH/U_SLAVE_1ELK/Q[2]\ : DFN1C0
      port map(D => \U_ELK14_CH/U_SLAVE_1ELK/ADJ_Q[2]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK14_CH/U_SLAVE_1ELK/Q[2]_net_1\);
    
    \U50_PATTERNS/U4C_REGCROSS/SAMP_ONE[1]\ : DFN1C0
      port map(D => \U50_PATTERNS/ELINKS_STRT_ADDR[1]\, CLK => 
        CLK_40M_GL, CLR => P_MASTER_POR_B_c_33, Q => 
        \U50_PATTERNS/U4C_REGCROSS/SAMP_ONE[1]_net_1\);
    
    HIEFFPLA_INST_0_40810 : MX2
      port map(A => HIEFFPLA_NET_0_119578, B => 
        \U50_PATTERNS/ELINK_DINA_17[0]\, S => 
        HIEFFPLA_NET_0_119260, Y => HIEFFPLA_NET_0_119807);
    
    HIEFFPLA_INST_0_57645 : XA1B
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_5[1]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_CNT_5[0]\, C => 
        HIEFFPLA_NET_0_117179, Y => HIEFFPLA_NET_0_116644);
    
    \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[5]\ : DFN1C0
      port map(D => 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[5]_net_1\, CLK
         => CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK18_CH/U_SLAVE_1ELK/ARB_BYTE[5]_net_1\);
    
    HIEFFPLA_INST_0_48867 : NAND2B
      port map(A => \OP_MODE_c_5[1]\, B => \PATT_ELK_DAT_19[3]\, 
        Y => HIEFFPLA_NET_0_118235);
    
    HIEFFPLA_INST_0_42927 : NAND3A
      port map(A => \U50_PATTERNS/REG_STATE[2]_net_1\, B => 
        \U50_PATTERNS/REG_STATE[5]_net_1\, C => 
        HIEFFPLA_NET_0_119393, Y => HIEFFPLA_NET_0_119423);
    
    HIEFFPLA_INST_0_37219 : AO1
      port map(A => \OP_MODE_c[2]\, B => 
        \U200A_TFC/GP_PG_SM[0]_net_1\, C => 
        \U200A_TFC/GP_PG_SM[1]_net_1\, Y => HIEFFPLA_NET_0_120322);
    
    HIEFFPLA_INST_0_62568 : MX2
      port map(A => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_7[2]\, 
        B => \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_8[2]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[0]\, Y => 
        HIEFFPLA_NET_0_115973);
    
    HIEFFPLA_INST_0_52423 : MX2
      port map(A => HIEFFPLA_NET_0_117517, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_29[3]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[3]\, Y => 
        HIEFFPLA_NET_0_117565);
    
    HIEFFPLA_INST_0_45109 : MX2
      port map(A => HIEFFPLA_NET_0_118973, B => 
        \U50_PATTERNS/WR_USB_ADBUS[3]\, S => 
        HIEFFPLA_NET_0_119486, Y => HIEFFPLA_NET_0_118982);
    
    HIEFFPLA_INST_0_41962 : NAND2B
      port map(A => \U50_PATTERNS/ELINK_RWA[4]\, B => 
        HIEFFPLA_NET_0_119643, Y => HIEFFPLA_NET_0_119644);
    
    \U_ELK10_CH/U_SLAVE_1ELK/Q[6]\ : DFN1C0
      port map(D => \U_ELK10_CH/U_SLAVE_1ELK/ADJ_Q[6]_net_1\, CLK
         => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/Q[6]_net_1\);
    
    HIEFFPLA_INST_0_52648 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_13[3]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/BIT_OS_VAL_14[3]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_2[0]\, Y => 
        HIEFFPLA_NET_0_117533);
    
    HIEFFPLA_INST_0_61532 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_23[4]\, B => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_24[4]\, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[0]\, Y => 
        HIEFFPLA_NET_0_116114);
    
    HIEFFPLA_INST_0_38418 : MX2
      port map(A => \U50_PATTERNS/ELINKS_STRT_ADDR[6]\, B => 
        \U50_PATTERNS/ELINKS_STRT_ADDR_T[6]\, S => 
        HIEFFPLA_NET_0_119472, Y => HIEFFPLA_NET_0_120105);
    
    \U_ELK10_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]\ : DFN1C0
      port map(D => \U_ELK10_CH/U_SLAVE_1ELK/Q[8]_net_1\, CLK => 
        CLK_40M_GL, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK10_CH/U_SLAVE_1ELK/ARB_WRD_40M_FIXED[8]_net_1\);
    
    HIEFFPLA_INST_0_45628 : NAND3C
      port map(A => HIEFFPLA_NET_0_118721, B => 
        HIEFFPLA_NET_0_118894, C => HIEFFPLA_NET_0_118711, Y => 
        HIEFFPLA_NET_0_118878);
    
    AFLSDF_INV_33 : INV
      port map(A => DCB_SALT_SEL_c, Y => \AFLSDF_INV_33\);
    
    \U_ELK8_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U0\ : IOPADP_BI
      port map(N2PIN => 
        \U_ELK8_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/U2_N2P\, D => 
        \U_ELK8_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET1\, E => 
        \U_ELK8_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET2\, PAD => 
        ELK8_DAT_P, Y => 
        \U_ELK8_CH/U_DDR_ELK1/BIBUF_LVDS_0/U0/NET4\);
    
    HIEFFPLA_INST_0_53102 : MX2
      port map(A => HIEFFPLA_NET_0_117553, B => 
        HIEFFPLA_NET_0_117549, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[2]\, Y => 
        HIEFFPLA_NET_0_117465);
    
    HIEFFPLA_INST_0_53054 : MX2
      port map(A => HIEFFPLA_NET_0_117563, B => 
        HIEFFPLA_NET_0_117559, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT_0[2]\, Y => 
        HIEFFPLA_NET_0_117471);
    
    HIEFFPLA_INST_0_52950 : MX2
      port map(A => HIEFFPLA_NET_0_117472, B => 
        HIEFFPLA_NET_0_117468, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/INDEX_CNT[4]\, Y => 
        HIEFFPLA_NET_0_117484);
    
    HIEFFPLA_INST_0_52326 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/BEST_BIT_OS_VAL[0]\, B
         => HIEFFPLA_NET_0_117576, S => HIEFFPLA_NET_0_117111, Y
         => HIEFFPLA_NET_0_117580);
    
    HIEFFPLA_INST_0_41260 : MX2
      port map(A => \U50_PATTERNS/ELINK_DINA_4[2]\, B => 
        HIEFFPLA_NET_0_119575, S => HIEFFPLA_NET_0_119284, Y => 
        HIEFFPLA_NET_0_119757);
    
    HIEFFPLA_INST_0_47656 : MX2
      port map(A => \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[4]_net_1\, 
        B => \U_ELK14_CH/U_SLAVE_1ELK/ARB_BYTE[8]_net_1\, S => 
        \BIT_OS_SEL_2[2]\, Y => HIEFFPLA_NET_0_118451);
    
    \U_ELK11_CH/U_SLAVE_1ELK/Q[14]\ : DFN1C0
      port map(D => \U_ELK11_CH/U_SLAVE_1ELK/ADJ_Q[14]_net_1\, 
        CLK => CCC_160M_FXD, CLR => MASTER_DCB_POR_B_i_0_i, Q => 
        \U_ELK11_CH/U_SLAVE_1ELK/Q[14]_net_1\);
    
    HIEFFPLA_INST_0_60666 : MX2
      port map(A => 
        \U_MASTER_DES/U13C_MASTER_DESER/SEQCNTS_14[0]\, B => 
        HIEFFPLA_NET_0_117190, S => HIEFFPLA_NET_0_117228, Y => 
        HIEFFPLA_NET_0_116235);
    
    HIEFFPLA_INST_0_47350 : AND2
      port map(A => \U_ELK13_CH/ELK_TX_DAT[1]\, B => 
        \U_ELK13_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118513);
    
    \U200B_ELINKS/ADDR_POINTER_0[6]\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_120171, CLK => CLK_40M_GL, CLR
         => P_MASTER_POR_B_c_32_0, Q => \ELKS_ADDRB_0[6]\);
    
    HIEFFPLA_INST_0_48611 : MX2
      port map(A => 
        \U_ELK18_CH/U_ELK1_CMD_TX/SER_CMD_WORD_R[2]_net_1\, B => 
        \U_ELK18_CH/ELK_TX_DAT[7]\, S => 
        \U_ELK18_CH/U_ELK1_CMD_TX/START_RISE_net_1\, Y => 
        HIEFFPLA_NET_0_118285);
    
    HIEFFPLA_INST_0_53755 : MX2
      port map(A => HIEFFPLA_NET_0_116125, B => 
        HIEFFPLA_NET_0_116023, S => 
        \U_MASTER_DES/U13C_MASTER_DESER/CLKPHASE_0[3]_net_1\, Y
         => HIEFFPLA_NET_0_117358);
    
    HIEFFPLA_INST_0_59705 : OA1A
      port map(A => HIEFFPLA_NET_0_116687, B => 
        HIEFFPLA_NET_0_117206, C => HIEFFPLA_NET_0_116357, Y => 
        HIEFFPLA_NET_0_116358);
    
    HIEFFPLA_INST_0_49523 : MX2
      port map(A => HIEFFPLA_NET_0_118127, B => 
        HIEFFPLA_NET_0_118140, S => \BIT_OS_SEL_1[0]\, Y => 
        \U_ELK2_CH/U_SLAVE_1ELK/N_RECD_SER_WORD[5]\);
    
    \U_ELK4_CH/ELK_IN_R\ : DFN1C0
      port map(D => \AFLSDF_INV_68\, CLK => CCC_160M_ADJ, CLR => 
        DEV_RST_B_c, Q => \U_ELK4_CH/ELK_IN_R_net_1\);
    
    HIEFFPLA_INST_0_45338 : AND3A
      port map(A => HIEFFPLA_NET_0_119444, B => 
        \U50_PATTERNS/ELINK_DOUTA_18[1]\, C => 
        \U50_PATTERNS/SM_BANK_SEL[1]\, Y => HIEFFPLA_NET_0_118936);
    
    GND_power_inst1 : GND
      port map( Y => GND_power_net1);

    VCC_power_inst1 : VCC
      port map( Y => VCC_power_net1);


end DEF_ARCH; 
